/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module selector4(
    input CLK,
    input [31:0] DATA_A,
    input [31:0] DATA_B,
    output [15:0] NIBBLE_OUT,
    input RESET_L,
    input [3:0] SEL,
    input [11:0] sel_A,
    input [11:0] sel_B
);

wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _512_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire _488_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire sel_A_5_bF$buf0 ;
wire sel_A_5_bF$buf1 ;
wire sel_A_5_bF$buf2 ;
wire sel_A_5_bF$buf3 ;
wire sel_A_5_bF$buf4 ;
wire _600_ ;
wire _197_ ;
wire [15:0] NIBBLE_OUT ;
wire _7_ ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire _285_ ;
wire [3:0] _1_ ;
wire _42_ ;
wire _379_ ;
wire sel_B_5_bF$buf0 ;
wire sel_B_5_bF$buf1 ;
wire sel_B_5_bF$buf2 ;
wire sel_B_5_bF$buf3 ;
wire sel_B_5_bF$buf4 ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire sel_A_11_bF$buf0 ;
wire sel_A_11_bF$buf1 ;
wire sel_A_11_bF$buf2 ;
wire sel_A_11_bF$buf3 ;
wire sel_A_11_bF$buf4 ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _517_ ;
wire _270_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire sel_A_2_bF$buf0 ;
wire sel_A_2_bF$buf1 ;
wire sel_A_2_bF$buf2 ;
wire sel_A_2_bF$buf3 ;
wire sel_A_2_bF$buf4 ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire [3:0] SEL ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire sel_B_2_bF$buf0 ;
wire sel_B_2_bF$buf1 ;
wire sel_B_2_bF$buf2 ;
wire sel_B_2_bF$buf3 ;
wire sel_B_2_bF$buf4 ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire [3:0] _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire [15:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _240_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _272_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _269_ ;
wire _498_ ;
wire _26_ ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _228_ ;
wire RESET_L ;
wire _457_ ;
wire _266_ ;
wire CLK ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _513_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire _454_ ;
wire _263_ ;
wire [3:0] _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _260_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire [3:0] _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire [31:0] DATA_A ;
wire [31:0] DATA_B ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire [11:0] sel_A ;
wire [11:0] sel_B ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire sel_B_11_bF$buf0 ;
wire sel_B_11_bF$buf1 ;
wire sel_B_11_bF$buf2 ;
wire sel_B_11_bF$buf3 ;
wire sel_B_11_bF$buf4 ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire sel_A_8_bF$buf0 ;
wire sel_A_8_bF$buf1 ;
wire sel_A_8_bF$buf2 ;
wire sel_A_8_bF$buf3 ;
wire sel_A_8_bF$buf4 ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _524_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire sel_B_8_bF$buf0 ;
wire sel_B_8_bF$buf1 ;
wire sel_B_8_bF$buf2 ;
wire sel_B_8_bF$buf3 ;
wire sel_B_8_bF$buf4 ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _518_ ;
wire _271_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _230_ ;
wire _515_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert39 (
    .A(sel_B[11]),
    .Y(sel_B_11_bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .A(sel_B[11]),
    .Y(sel_B_11_bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .A(sel_B[11]),
    .Y(sel_B_11_bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .A(sel_B[11]),
    .Y(sel_B_11_bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .A(sel_B[11]),
    .Y(sel_B_11_bF$buf4)
);

BUFX2 BUFX2_insert34 (
    .A(sel_A[2]),
    .Y(sel_A_2_bF$buf0)
);

BUFX2 BUFX2_insert33 (
    .A(sel_A[2]),
    .Y(sel_A_2_bF$buf1)
);

BUFX2 BUFX2_insert32 (
    .A(sel_A[2]),
    .Y(sel_A_2_bF$buf2)
);

BUFX2 BUFX2_insert31 (
    .A(sel_A[2]),
    .Y(sel_A_2_bF$buf3)
);

BUFX2 BUFX2_insert30 (
    .A(sel_A[2]),
    .Y(sel_A_2_bF$buf4)
);

BUFX2 BUFX2_insert29 (
    .A(sel_A[5]),
    .Y(sel_A_5_bF$buf0)
);

BUFX2 BUFX2_insert28 (
    .A(sel_A[5]),
    .Y(sel_A_5_bF$buf1)
);

BUFX2 BUFX2_insert27 (
    .A(sel_A[5]),
    .Y(sel_A_5_bF$buf2)
);

BUFX2 BUFX2_insert26 (
    .A(sel_A[5]),
    .Y(sel_A_5_bF$buf3)
);

BUFX2 BUFX2_insert25 (
    .A(sel_A[5]),
    .Y(sel_A_5_bF$buf4)
);

BUFX2 BUFX2_insert24 (
    .A(sel_B[2]),
    .Y(sel_B_2_bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(sel_B[2]),
    .Y(sel_B_2_bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(sel_B[2]),
    .Y(sel_B_2_bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(sel_B[2]),
    .Y(sel_B_2_bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(sel_B[2]),
    .Y(sel_B_2_bF$buf4)
);

BUFX2 BUFX2_insert19 (
    .A(sel_A[8]),
    .Y(sel_A_8_bF$buf0)
);

BUFX2 BUFX2_insert18 (
    .A(sel_A[8]),
    .Y(sel_A_8_bF$buf1)
);

BUFX2 BUFX2_insert17 (
    .A(sel_A[8]),
    .Y(sel_A_8_bF$buf2)
);

BUFX2 BUFX2_insert16 (
    .A(sel_A[8]),
    .Y(sel_A_8_bF$buf3)
);

BUFX2 BUFX2_insert15 (
    .A(sel_A[8]),
    .Y(sel_A_8_bF$buf4)
);

BUFX2 BUFX2_insert14 (
    .A(sel_B[5]),
    .Y(sel_B_5_bF$buf0)
);

BUFX2 BUFX2_insert13 (
    .A(sel_B[5]),
    .Y(sel_B_5_bF$buf1)
);

BUFX2 BUFX2_insert12 (
    .A(sel_B[5]),
    .Y(sel_B_5_bF$buf2)
);

BUFX2 BUFX2_insert11 (
    .A(sel_B[5]),
    .Y(sel_B_5_bF$buf3)
);

BUFX2 BUFX2_insert10 (
    .A(sel_B[5]),
    .Y(sel_B_5_bF$buf4)
);

BUFX2 BUFX2_insert9 (
    .A(sel_B[8]),
    .Y(sel_B_8_bF$buf0)
);

BUFX2 BUFX2_insert8 (
    .A(sel_B[8]),
    .Y(sel_B_8_bF$buf1)
);

BUFX2 BUFX2_insert7 (
    .A(sel_B[8]),
    .Y(sel_B_8_bF$buf2)
);

BUFX2 BUFX2_insert6 (
    .A(sel_B[8]),
    .Y(sel_B_8_bF$buf3)
);

BUFX2 BUFX2_insert5 (
    .A(sel_B[8]),
    .Y(sel_B_8_bF$buf4)
);

BUFX2 BUFX2_insert4 (
    .A(sel_A[11]),
    .Y(sel_A_11_bF$buf0)
);

BUFX2 BUFX2_insert3 (
    .A(sel_A[11]),
    .Y(sel_A_11_bF$buf1)
);

BUFX2 BUFX2_insert2 (
    .A(sel_A[11]),
    .Y(sel_A_11_bF$buf2)
);

BUFX2 BUFX2_insert1 (
    .A(sel_A[11]),
    .Y(sel_A_11_bF$buf3)
);

BUFX2 BUFX2_insert0 (
    .A(sel_A[11]),
    .Y(sel_A_11_bF$buf4)
);

NAND2X1 _1000_ (
    .A(sel_A_8_bF$buf4),
    .B(_469_),
    .Y(_470_)
);

NAND3X1 _1001_ (
    .A(_458_),
    .B(_468_),
    .C(_470_),
    .Y(_471_)
);

INVX1 _1002_ (
    .A(DATA_A[12]),
    .Y(_472_)
);

NAND2X1 _1003_ (
    .A(sel_A_8_bF$buf3),
    .B(DATA_A[28]),
    .Y(_473_)
);

OAI21X1 _1004_ (
    .A(_472_),
    .B(sel_A_8_bF$buf2),
    .C(_473_),
    .Y(_474_)
);

NAND2X1 _1005_ (
    .A(sel_A[7]),
    .B(_474_),
    .Y(_475_)
);

NAND3X1 _1006_ (
    .A(sel_A[6]),
    .B(_471_),
    .C(_475_),
    .Y(_476_)
);

NAND3X1 _1007_ (
    .A(_456_),
    .B(_467_),
    .C(_476_),
    .Y(_477_)
);

INVX2 _1008_ (
    .A(sel_B[6]),
    .Y(_320_)
);

INVX4 _1009_ (
    .A(sel_B[7]),
    .Y(_321_)
);

OR2X2 _1010_ (
    .A(DATA_B[0]),
    .B(sel_B_8_bF$buf4),
    .Y(_322_)
);

INVX1 _1011_ (
    .A(DATA_B[16]),
    .Y(_323_)
);

NAND2X1 _1012_ (
    .A(sel_B_8_bF$buf3),
    .B(_323_),
    .Y(_324_)
);

NAND3X1 _1013_ (
    .A(_321_),
    .B(_322_),
    .C(_324_),
    .Y(_325_)
);

INVX1 _1014_ (
    .A(DATA_B[24]),
    .Y(_326_)
);

NAND2X1 _1015_ (
    .A(sel_B_8_bF$buf2),
    .B(_326_),
    .Y(_327_)
);

OR2X2 _1016_ (
    .A(sel_B_8_bF$buf1),
    .B(DATA_B[8]),
    .Y(_328_)
);

NAND3X1 _1017_ (
    .A(sel_B[7]),
    .B(_328_),
    .C(_327_),
    .Y(_329_)
);

NAND3X1 _1018_ (
    .A(_320_),
    .B(_325_),
    .C(_329_),
    .Y(_330_)
);

OR2X2 _1019_ (
    .A(sel_B_8_bF$buf0),
    .B(DATA_B[4]),
    .Y(_331_)
);

INVX1 _1020_ (
    .A(DATA_B[20]),
    .Y(_332_)
);

NAND2X1 _1021_ (
    .A(sel_B_8_bF$buf4),
    .B(_332_),
    .Y(_333_)
);

NAND3X1 _1022_ (
    .A(_321_),
    .B(_331_),
    .C(_333_),
    .Y(_334_)
);

INVX1 _1023_ (
    .A(DATA_B[12]),
    .Y(_335_)
);

NAND2X1 _1024_ (
    .A(sel_B_8_bF$buf3),
    .B(DATA_B[28]),
    .Y(_336_)
);

OAI21X1 _1025_ (
    .A(_335_),
    .B(sel_B_8_bF$buf2),
    .C(_336_),
    .Y(_337_)
);

NAND2X1 _1026_ (
    .A(sel_B[7]),
    .B(_337_),
    .Y(_338_)
);

NAND3X1 _1027_ (
    .A(sel_B[6]),
    .B(_334_),
    .C(_338_),
    .Y(_339_)
);

NAND3X1 _1028_ (
    .A(SEL[2]),
    .B(_330_),
    .C(_339_),
    .Y(_340_)
);

AOI21X1 _1029_ (
    .A(_477_),
    .B(_340_),
    .C(_455_),
    .Y(_319_[0])
);

OR2X2 _1030_ (
    .A(sel_A_8_bF$buf1),
    .B(DATA_A[1]),
    .Y(_341_)
);

INVX1 _1031_ (
    .A(DATA_A[17]),
    .Y(_342_)
);

NAND2X1 _1032_ (
    .A(sel_A_8_bF$buf0),
    .B(_342_),
    .Y(_343_)
);

NAND3X1 _1033_ (
    .A(_458_),
    .B(_341_),
    .C(_343_),
    .Y(_344_)
);

INVX1 _1034_ (
    .A(DATA_A[25]),
    .Y(_345_)
);

NAND2X1 _1035_ (
    .A(sel_A_8_bF$buf4),
    .B(_345_),
    .Y(_346_)
);

OR2X2 _1036_ (
    .A(sel_A_8_bF$buf3),
    .B(DATA_A[9]),
    .Y(_347_)
);

NAND3X1 _1037_ (
    .A(sel_A[7]),
    .B(_347_),
    .C(_346_),
    .Y(_348_)
);

NAND3X1 _1038_ (
    .A(_457_),
    .B(_344_),
    .C(_348_),
    .Y(_349_)
);

OR2X2 _1039_ (
    .A(sel_A_8_bF$buf2),
    .B(DATA_A[5]),
    .Y(_350_)
);

INVX1 _1040_ (
    .A(DATA_A[21]),
    .Y(_351_)
);

NAND2X1 _1041_ (
    .A(sel_A_8_bF$buf1),
    .B(_351_),
    .Y(_352_)
);

NAND3X1 _1042_ (
    .A(_458_),
    .B(_350_),
    .C(_352_),
    .Y(_353_)
);

INVX1 _1043_ (
    .A(DATA_A[13]),
    .Y(_354_)
);

NAND2X1 _1044_ (
    .A(sel_A_8_bF$buf0),
    .B(DATA_A[29]),
    .Y(_355_)
);

OAI21X1 _1045_ (
    .A(_354_),
    .B(sel_A_8_bF$buf4),
    .C(_355_),
    .Y(_356_)
);

NAND2X1 _1046_ (
    .A(sel_A[7]),
    .B(_356_),
    .Y(_357_)
);

NAND3X1 _1047_ (
    .A(sel_A[6]),
    .B(_353_),
    .C(_357_),
    .Y(_358_)
);

NAND3X1 _1048_ (
    .A(_456_),
    .B(_349_),
    .C(_358_),
    .Y(_359_)
);

OR2X2 _1049_ (
    .A(sel_B_8_bF$buf1),
    .B(DATA_B[1]),
    .Y(_360_)
);

INVX1 _1050_ (
    .A(DATA_B[17]),
    .Y(_361_)
);

NAND2X1 _1051_ (
    .A(sel_B_8_bF$buf0),
    .B(_361_),
    .Y(_362_)
);

NAND3X1 _1052_ (
    .A(_321_),
    .B(_360_),
    .C(_362_),
    .Y(_363_)
);

INVX1 _1053_ (
    .A(DATA_B[25]),
    .Y(_364_)
);

NAND2X1 _1054_ (
    .A(sel_B_8_bF$buf4),
    .B(_364_),
    .Y(_365_)
);

OR2X2 _1055_ (
    .A(sel_B_8_bF$buf3),
    .B(DATA_B[9]),
    .Y(_366_)
);

NAND3X1 _1056_ (
    .A(sel_B[7]),
    .B(_366_),
    .C(_365_),
    .Y(_367_)
);

NAND3X1 _1057_ (
    .A(_320_),
    .B(_363_),
    .C(_367_),
    .Y(_368_)
);

OR2X2 _1058_ (
    .A(sel_B_8_bF$buf2),
    .B(DATA_B[5]),
    .Y(_369_)
);

INVX1 _1059_ (
    .A(DATA_B[21]),
    .Y(_370_)
);

NAND2X1 _1060_ (
    .A(sel_B_8_bF$buf1),
    .B(_370_),
    .Y(_371_)
);

NAND3X1 _1061_ (
    .A(_321_),
    .B(_369_),
    .C(_371_),
    .Y(_372_)
);

INVX1 _1062_ (
    .A(DATA_B[13]),
    .Y(_373_)
);

NAND2X1 _1063_ (
    .A(sel_B_8_bF$buf0),
    .B(DATA_B[29]),
    .Y(_374_)
);

OAI21X1 _1064_ (
    .A(_373_),
    .B(sel_B_8_bF$buf4),
    .C(_374_),
    .Y(_375_)
);

NAND2X1 _1065_ (
    .A(sel_B[7]),
    .B(_375_),
    .Y(_376_)
);

NAND3X1 _1066_ (
    .A(sel_B[6]),
    .B(_372_),
    .C(_376_),
    .Y(_377_)
);

NAND3X1 _1067_ (
    .A(SEL[2]),
    .B(_368_),
    .C(_377_),
    .Y(_378_)
);

AOI21X1 _1068_ (
    .A(_359_),
    .B(_378_),
    .C(_455_),
    .Y(_319_[1])
);

OR2X2 _1069_ (
    .A(sel_A_8_bF$buf3),
    .B(DATA_A[2]),
    .Y(_379_)
);

INVX1 _1070_ (
    .A(DATA_A[18]),
    .Y(_380_)
);

NAND2X1 _1071_ (
    .A(sel_A_8_bF$buf2),
    .B(_380_),
    .Y(_381_)
);

NAND3X1 _1072_ (
    .A(_458_),
    .B(_379_),
    .C(_381_),
    .Y(_382_)
);

INVX1 _1073_ (
    .A(DATA_A[26]),
    .Y(_383_)
);

NAND2X1 _1074_ (
    .A(sel_A_8_bF$buf1),
    .B(_383_),
    .Y(_384_)
);

OR2X2 _1075_ (
    .A(sel_A_8_bF$buf0),
    .B(DATA_A[10]),
    .Y(_385_)
);

NAND3X1 _1076_ (
    .A(sel_A[7]),
    .B(_385_),
    .C(_384_),
    .Y(_386_)
);

NAND3X1 _1077_ (
    .A(_457_),
    .B(_382_),
    .C(_386_),
    .Y(_387_)
);

OR2X2 _1078_ (
    .A(sel_A_8_bF$buf4),
    .B(DATA_A[6]),
    .Y(_388_)
);

INVX1 _1079_ (
    .A(DATA_A[22]),
    .Y(_389_)
);

NAND2X1 _1080_ (
    .A(sel_A_8_bF$buf3),
    .B(_389_),
    .Y(_390_)
);

NAND3X1 _1081_ (
    .A(_458_),
    .B(_388_),
    .C(_390_),
    .Y(_391_)
);

INVX1 _1082_ (
    .A(DATA_A[14]),
    .Y(_392_)
);

NAND2X1 _1083_ (
    .A(sel_A_8_bF$buf2),
    .B(DATA_A[30]),
    .Y(_393_)
);

OAI21X1 _1084_ (
    .A(_392_),
    .B(sel_A_8_bF$buf1),
    .C(_393_),
    .Y(_394_)
);

NAND2X1 _1085_ (
    .A(sel_A[7]),
    .B(_394_),
    .Y(_395_)
);

NAND3X1 _1086_ (
    .A(sel_A[6]),
    .B(_391_),
    .C(_395_),
    .Y(_396_)
);

NAND3X1 _1087_ (
    .A(_456_),
    .B(_387_),
    .C(_396_),
    .Y(_397_)
);

OR2X2 _1088_ (
    .A(sel_B_8_bF$buf3),
    .B(DATA_B[6]),
    .Y(_398_)
);

INVX1 _1089_ (
    .A(DATA_B[22]),
    .Y(_399_)
);

NAND2X1 _1090_ (
    .A(sel_B_8_bF$buf2),
    .B(_399_),
    .Y(_400_)
);

NAND3X1 _1091_ (
    .A(_321_),
    .B(_398_),
    .C(_400_),
    .Y(_401_)
);

INVX1 _1092_ (
    .A(DATA_B[30]),
    .Y(_402_)
);

NAND2X1 _1093_ (
    .A(sel_B_8_bF$buf1),
    .B(_402_),
    .Y(_403_)
);

OR2X2 _1094_ (
    .A(sel_B_8_bF$buf0),
    .B(DATA_B[14]),
    .Y(_404_)
);

NAND3X1 _1095_ (
    .A(sel_B[7]),
    .B(_404_),
    .C(_403_),
    .Y(_405_)
);

NAND3X1 _1096_ (
    .A(sel_B[6]),
    .B(_401_),
    .C(_405_),
    .Y(_406_)
);

OR2X2 _1097_ (
    .A(sel_B_8_bF$buf4),
    .B(DATA_B[2]),
    .Y(_407_)
);

INVX1 _1098_ (
    .A(DATA_B[18]),
    .Y(_408_)
);

NAND2X1 _1099_ (
    .A(sel_B_8_bF$buf3),
    .B(_408_),
    .Y(_409_)
);

NAND3X1 _1100_ (
    .A(_321_),
    .B(_407_),
    .C(_409_),
    .Y(_410_)
);

INVX1 _1101_ (
    .A(DATA_B[10]),
    .Y(_411_)
);

NAND2X1 _1102_ (
    .A(sel_B_8_bF$buf2),
    .B(DATA_B[26]),
    .Y(_412_)
);

OAI21X1 _1103_ (
    .A(_411_),
    .B(sel_B_8_bF$buf1),
    .C(_412_),
    .Y(_413_)
);

NAND2X1 _1104_ (
    .A(sel_B[7]),
    .B(_413_),
    .Y(_414_)
);

NAND3X1 _1105_ (
    .A(_320_),
    .B(_410_),
    .C(_414_),
    .Y(_415_)
);

NAND3X1 _1106_ (
    .A(SEL[2]),
    .B(_406_),
    .C(_415_),
    .Y(_416_)
);

AOI21X1 _1107_ (
    .A(_397_),
    .B(_416_),
    .C(_455_),
    .Y(_319_[2])
);

OR2X2 _1108_ (
    .A(sel_A_8_bF$buf0),
    .B(DATA_A[3]),
    .Y(_417_)
);

INVX1 _1109_ (
    .A(DATA_A[19]),
    .Y(_418_)
);

NAND2X1 _1110_ (
    .A(sel_A_8_bF$buf4),
    .B(_418_),
    .Y(_419_)
);

NAND3X1 _1111_ (
    .A(_458_),
    .B(_417_),
    .C(_419_),
    .Y(_420_)
);

INVX1 _1112_ (
    .A(DATA_A[27]),
    .Y(_421_)
);

NAND2X1 _1113_ (
    .A(sel_A_8_bF$buf3),
    .B(_421_),
    .Y(_422_)
);

OR2X2 _1114_ (
    .A(sel_A_8_bF$buf2),
    .B(DATA_A[11]),
    .Y(_423_)
);

NAND3X1 _1115_ (
    .A(sel_A[7]),
    .B(_423_),
    .C(_422_),
    .Y(_424_)
);

NAND3X1 _1116_ (
    .A(_457_),
    .B(_420_),
    .C(_424_),
    .Y(_425_)
);

OR2X2 _1117_ (
    .A(sel_A_8_bF$buf1),
    .B(DATA_A[7]),
    .Y(_426_)
);

INVX1 _1118_ (
    .A(DATA_A[23]),
    .Y(_427_)
);

NAND2X1 _1119_ (
    .A(sel_A_8_bF$buf0),
    .B(_427_),
    .Y(_428_)
);

NAND3X1 _1120_ (
    .A(_458_),
    .B(_426_),
    .C(_428_),
    .Y(_429_)
);

INVX1 _1121_ (
    .A(DATA_A[15]),
    .Y(_430_)
);

NAND2X1 _1122_ (
    .A(sel_A_8_bF$buf4),
    .B(DATA_A[31]),
    .Y(_431_)
);

OAI21X1 _1123_ (
    .A(_430_),
    .B(sel_A_8_bF$buf3),
    .C(_431_),
    .Y(_432_)
);

NAND2X1 _1124_ (
    .A(sel_A[7]),
    .B(_432_),
    .Y(_433_)
);

NAND3X1 _1125_ (
    .A(sel_A[6]),
    .B(_429_),
    .C(_433_),
    .Y(_434_)
);

NAND3X1 _1126_ (
    .A(_456_),
    .B(_425_),
    .C(_434_),
    .Y(_435_)
);

OR2X2 _1127_ (
    .A(sel_B_8_bF$buf0),
    .B(DATA_B[3]),
    .Y(_436_)
);

INVX1 _1128_ (
    .A(DATA_B[19]),
    .Y(_437_)
);

NAND2X1 _1129_ (
    .A(sel_B_8_bF$buf4),
    .B(_437_),
    .Y(_438_)
);

NAND3X1 _1130_ (
    .A(_321_),
    .B(_436_),
    .C(_438_),
    .Y(_439_)
);

INVX1 _1131_ (
    .A(DATA_B[27]),
    .Y(_440_)
);

NAND2X1 _1132_ (
    .A(sel_B_8_bF$buf3),
    .B(_440_),
    .Y(_441_)
);

OR2X2 _1133_ (
    .A(sel_B_8_bF$buf2),
    .B(DATA_B[11]),
    .Y(_442_)
);

NAND3X1 _1134_ (
    .A(sel_B[7]),
    .B(_442_),
    .C(_441_),
    .Y(_443_)
);

NAND3X1 _1135_ (
    .A(_320_),
    .B(_439_),
    .C(_443_),
    .Y(_444_)
);

OR2X2 _1136_ (
    .A(sel_B_8_bF$buf1),
    .B(DATA_B[7]),
    .Y(_445_)
);

INVX1 _1137_ (
    .A(DATA_B[23]),
    .Y(_446_)
);

NAND2X1 _1138_ (
    .A(sel_B_8_bF$buf0),
    .B(_446_),
    .Y(_447_)
);

NAND3X1 _1139_ (
    .A(_321_),
    .B(_445_),
    .C(_447_),
    .Y(_448_)
);

INVX1 _1140_ (
    .A(DATA_B[15]),
    .Y(_449_)
);

NAND2X1 _1141_ (
    .A(sel_B_8_bF$buf4),
    .B(DATA_B[31]),
    .Y(_450_)
);

OAI21X1 _1142_ (
    .A(_449_),
    .B(sel_B_8_bF$buf3),
    .C(_450_),
    .Y(_451_)
);

NAND2X1 _1143_ (
    .A(sel_B[7]),
    .B(_451_),
    .Y(_452_)
);

NAND3X1 _1144_ (
    .A(sel_B[6]),
    .B(_448_),
    .C(_452_),
    .Y(_453_)
);

NAND3X1 _1145_ (
    .A(SEL[2]),
    .B(_444_),
    .C(_453_),
    .Y(_454_)
);

AOI21X1 _1146_ (
    .A(_435_),
    .B(_454_),
    .C(_455_),
    .Y(_319_[3])
);

DFFPOSX1 _1147_ (
    .CLK(CLK),
    .D(_319_[0]),
    .Q(_0_[8])
);

DFFPOSX1 _1148_ (
    .CLK(CLK),
    .D(_319_[1]),
    .Q(_0_[9])
);

DFFPOSX1 _1149_ (
    .CLK(CLK),
    .D(_319_[2]),
    .Q(_0_[10])
);

DFFPOSX1 _1150_ (
    .CLK(CLK),
    .D(_319_[3]),
    .Q(_0_[11])
);

INVX2 _1151_ (
    .A(RESET_L),
    .Y(_614_)
);

INVX2 _1152_ (
    .A(SEL[3]),
    .Y(_615_)
);

INVX2 _1153_ (
    .A(sel_A[9]),
    .Y(_616_)
);

INVX4 _1154_ (
    .A(sel_A[10]),
    .Y(_617_)
);

OR2X2 _1155_ (
    .A(DATA_A[0]),
    .B(sel_A_11_bF$buf4),
    .Y(_618_)
);

INVX1 _1156_ (
    .A(DATA_A[16]),
    .Y(_619_)
);

NAND2X1 _1157_ (
    .A(sel_A_11_bF$buf3),
    .B(_619_),
    .Y(_620_)
);

NAND3X1 _1158_ (
    .A(_617_),
    .B(_618_),
    .C(_620_),
    .Y(_621_)
);

INVX1 _1159_ (
    .A(DATA_A[24]),
    .Y(_622_)
);

NAND2X1 _1160_ (
    .A(sel_A_11_bF$buf2),
    .B(_622_),
    .Y(_623_)
);

OR2X2 _1161_ (
    .A(sel_A_11_bF$buf1),
    .B(DATA_A[8]),
    .Y(_624_)
);

NAND3X1 _1162_ (
    .A(sel_A[10]),
    .B(_624_),
    .C(_623_),
    .Y(_625_)
);

NAND3X1 _1163_ (
    .A(_616_),
    .B(_621_),
    .C(_625_),
    .Y(_626_)
);

OR2X2 _1164_ (
    .A(sel_A_11_bF$buf0),
    .B(DATA_A[4]),
    .Y(_627_)
);

INVX1 _1165_ (
    .A(DATA_A[20]),
    .Y(_628_)
);

NAND2X1 _1166_ (
    .A(sel_A_11_bF$buf4),
    .B(_628_),
    .Y(_629_)
);

NAND3X1 _1167_ (
    .A(_617_),
    .B(_627_),
    .C(_629_),
    .Y(_630_)
);

INVX1 _1168_ (
    .A(DATA_A[12]),
    .Y(_631_)
);

NAND2X1 _1169_ (
    .A(sel_A_11_bF$buf3),
    .B(DATA_A[28]),
    .Y(_632_)
);

OAI21X1 _1170_ (
    .A(_631_),
    .B(sel_A_11_bF$buf2),
    .C(_632_),
    .Y(_633_)
);

NAND2X1 _1171_ (
    .A(sel_A[10]),
    .B(_633_),
    .Y(_634_)
);

NAND3X1 _1172_ (
    .A(sel_A[9]),
    .B(_630_),
    .C(_634_),
    .Y(_635_)
);

NAND3X1 _1173_ (
    .A(_615_),
    .B(_626_),
    .C(_635_),
    .Y(_636_)
);

INVX2 _1174_ (
    .A(sel_B[9]),
    .Y(_479_)
);

INVX4 _1175_ (
    .A(sel_B[10]),
    .Y(_480_)
);

OR2X2 _1176_ (
    .A(DATA_B[0]),
    .B(sel_B_11_bF$buf4),
    .Y(_481_)
);

INVX1 _1177_ (
    .A(DATA_B[16]),
    .Y(_482_)
);

NAND2X1 _1178_ (
    .A(sel_B_11_bF$buf3),
    .B(_482_),
    .Y(_483_)
);

NAND3X1 _1179_ (
    .A(_480_),
    .B(_481_),
    .C(_483_),
    .Y(_484_)
);

INVX1 _1180_ (
    .A(DATA_B[24]),
    .Y(_485_)
);

NAND2X1 _1181_ (
    .A(sel_B_11_bF$buf2),
    .B(_485_),
    .Y(_486_)
);

OR2X2 _1182_ (
    .A(sel_B_11_bF$buf1),
    .B(DATA_B[8]),
    .Y(_487_)
);

NAND3X1 _1183_ (
    .A(sel_B[10]),
    .B(_487_),
    .C(_486_),
    .Y(_488_)
);

NAND3X1 _1184_ (
    .A(_479_),
    .B(_484_),
    .C(_488_),
    .Y(_489_)
);

OR2X2 _1185_ (
    .A(sel_B_11_bF$buf0),
    .B(DATA_B[4]),
    .Y(_490_)
);

INVX1 _1186_ (
    .A(DATA_B[20]),
    .Y(_491_)
);

NAND2X1 _1187_ (
    .A(sel_B_11_bF$buf4),
    .B(_491_),
    .Y(_492_)
);

NAND3X1 _1188_ (
    .A(_480_),
    .B(_490_),
    .C(_492_),
    .Y(_493_)
);

INVX1 _1189_ (
    .A(DATA_B[12]),
    .Y(_494_)
);

NAND2X1 _1190_ (
    .A(sel_B_11_bF$buf3),
    .B(DATA_B[28]),
    .Y(_495_)
);

OAI21X1 _1191_ (
    .A(_494_),
    .B(sel_B_11_bF$buf2),
    .C(_495_),
    .Y(_496_)
);

NAND2X1 _1192_ (
    .A(sel_B[10]),
    .B(_496_),
    .Y(_497_)
);

NAND3X1 _1193_ (
    .A(sel_B[9]),
    .B(_493_),
    .C(_497_),
    .Y(_498_)
);

NAND3X1 _1194_ (
    .A(SEL[3]),
    .B(_489_),
    .C(_498_),
    .Y(_499_)
);

AOI21X1 _1195_ (
    .A(_636_),
    .B(_499_),
    .C(_614_),
    .Y(_478_[0])
);

OR2X2 _1196_ (
    .A(sel_A_11_bF$buf1),
    .B(DATA_A[1]),
    .Y(_500_)
);

INVX1 _1197_ (
    .A(DATA_A[17]),
    .Y(_501_)
);

NAND2X1 _1198_ (
    .A(sel_A_11_bF$buf0),
    .B(_501_),
    .Y(_502_)
);

NAND3X1 _1199_ (
    .A(_617_),
    .B(_500_),
    .C(_502_),
    .Y(_503_)
);

INVX1 _1200_ (
    .A(DATA_A[25]),
    .Y(_504_)
);

NAND2X1 _1201_ (
    .A(sel_A_11_bF$buf4),
    .B(_504_),
    .Y(_505_)
);

OR2X2 _1202_ (
    .A(sel_A_11_bF$buf3),
    .B(DATA_A[9]),
    .Y(_506_)
);

NAND3X1 _1203_ (
    .A(sel_A[10]),
    .B(_506_),
    .C(_505_),
    .Y(_507_)
);

NAND3X1 _1204_ (
    .A(_616_),
    .B(_503_),
    .C(_507_),
    .Y(_508_)
);

OR2X2 _1205_ (
    .A(sel_A_11_bF$buf2),
    .B(DATA_A[5]),
    .Y(_509_)
);

INVX1 _1206_ (
    .A(DATA_A[21]),
    .Y(_510_)
);

NAND2X1 _1207_ (
    .A(sel_A_11_bF$buf1),
    .B(_510_),
    .Y(_511_)
);

NAND3X1 _1208_ (
    .A(_617_),
    .B(_509_),
    .C(_511_),
    .Y(_512_)
);

INVX1 _1209_ (
    .A(DATA_A[13]),
    .Y(_513_)
);

NAND2X1 _1210_ (
    .A(sel_A_11_bF$buf0),
    .B(DATA_A[29]),
    .Y(_514_)
);

OAI21X1 _1211_ (
    .A(_513_),
    .B(sel_A_11_bF$buf4),
    .C(_514_),
    .Y(_515_)
);

NAND2X1 _1212_ (
    .A(sel_A[10]),
    .B(_515_),
    .Y(_516_)
);

NAND3X1 _1213_ (
    .A(sel_A[9]),
    .B(_512_),
    .C(_516_),
    .Y(_517_)
);

NAND3X1 _1214_ (
    .A(_615_),
    .B(_508_),
    .C(_517_),
    .Y(_518_)
);

OR2X2 _1215_ (
    .A(sel_B_11_bF$buf1),
    .B(DATA_B[1]),
    .Y(_519_)
);

INVX1 _1216_ (
    .A(DATA_B[17]),
    .Y(_520_)
);

NAND2X1 _1217_ (
    .A(sel_B_11_bF$buf0),
    .B(_520_),
    .Y(_521_)
);

NAND3X1 _1218_ (
    .A(_480_),
    .B(_519_),
    .C(_521_),
    .Y(_522_)
);

INVX1 _1219_ (
    .A(DATA_B[25]),
    .Y(_523_)
);

NAND2X1 _1220_ (
    .A(sel_B_11_bF$buf4),
    .B(_523_),
    .Y(_524_)
);

OR2X2 _1221_ (
    .A(sel_B_11_bF$buf3),
    .B(DATA_B[9]),
    .Y(_525_)
);

NAND3X1 _1222_ (
    .A(sel_B[10]),
    .B(_525_),
    .C(_524_),
    .Y(_526_)
);

NAND3X1 _1223_ (
    .A(_479_),
    .B(_522_),
    .C(_526_),
    .Y(_527_)
);

OR2X2 _1224_ (
    .A(sel_B_11_bF$buf2),
    .B(DATA_B[5]),
    .Y(_528_)
);

INVX1 _1225_ (
    .A(DATA_B[21]),
    .Y(_529_)
);

NAND2X1 _1226_ (
    .A(sel_B_11_bF$buf1),
    .B(_529_),
    .Y(_530_)
);

NAND3X1 _1227_ (
    .A(_480_),
    .B(_528_),
    .C(_530_),
    .Y(_531_)
);

INVX1 _1228_ (
    .A(DATA_B[13]),
    .Y(_532_)
);

NAND2X1 _1229_ (
    .A(sel_B_11_bF$buf0),
    .B(DATA_B[29]),
    .Y(_533_)
);

OAI21X1 _1230_ (
    .A(_532_),
    .B(sel_B_11_bF$buf4),
    .C(_533_),
    .Y(_534_)
);

NAND2X1 _1231_ (
    .A(sel_B[10]),
    .B(_534_),
    .Y(_535_)
);

NAND3X1 _1232_ (
    .A(sel_B[9]),
    .B(_531_),
    .C(_535_),
    .Y(_536_)
);

NAND3X1 _1233_ (
    .A(SEL[3]),
    .B(_527_),
    .C(_536_),
    .Y(_537_)
);

AOI21X1 _1234_ (
    .A(_518_),
    .B(_537_),
    .C(_614_),
    .Y(_478_[1])
);

OR2X2 _1235_ (
    .A(sel_A_11_bF$buf3),
    .B(DATA_A[2]),
    .Y(_538_)
);

INVX1 _1236_ (
    .A(DATA_A[18]),
    .Y(_539_)
);

NAND2X1 _1237_ (
    .A(sel_A_11_bF$buf2),
    .B(_539_),
    .Y(_540_)
);

NAND3X1 _1238_ (
    .A(_617_),
    .B(_538_),
    .C(_540_),
    .Y(_541_)
);

INVX1 _1239_ (
    .A(DATA_A[26]),
    .Y(_542_)
);

NAND2X1 _1240_ (
    .A(sel_A_11_bF$buf1),
    .B(_542_),
    .Y(_543_)
);

OR2X2 _1241_ (
    .A(sel_A_11_bF$buf0),
    .B(DATA_A[10]),
    .Y(_544_)
);

NAND3X1 _1242_ (
    .A(sel_A[10]),
    .B(_544_),
    .C(_543_),
    .Y(_545_)
);

NAND3X1 _1243_ (
    .A(_616_),
    .B(_541_),
    .C(_545_),
    .Y(_546_)
);

OR2X2 _1244_ (
    .A(sel_A_11_bF$buf4),
    .B(DATA_A[6]),
    .Y(_547_)
);

INVX1 _1245_ (
    .A(DATA_A[22]),
    .Y(_548_)
);

NAND2X1 _1246_ (
    .A(sel_A_11_bF$buf3),
    .B(_548_),
    .Y(_549_)
);

NAND3X1 _1247_ (
    .A(_617_),
    .B(_547_),
    .C(_549_),
    .Y(_550_)
);

INVX1 _1248_ (
    .A(DATA_A[14]),
    .Y(_551_)
);

NAND2X1 _1249_ (
    .A(sel_A_11_bF$buf2),
    .B(DATA_A[30]),
    .Y(_552_)
);

OAI21X1 _1250_ (
    .A(_551_),
    .B(sel_A_11_bF$buf1),
    .C(_552_),
    .Y(_553_)
);

NAND2X1 _1251_ (
    .A(sel_A[10]),
    .B(_553_),
    .Y(_554_)
);

NAND3X1 _1252_ (
    .A(sel_A[9]),
    .B(_550_),
    .C(_554_),
    .Y(_555_)
);

NAND3X1 _1253_ (
    .A(_615_),
    .B(_546_),
    .C(_555_),
    .Y(_556_)
);

OR2X2 _1254_ (
    .A(sel_B_11_bF$buf3),
    .B(DATA_B[6]),
    .Y(_557_)
);

INVX1 _1255_ (
    .A(DATA_B[22]),
    .Y(_558_)
);

NAND2X1 _1256_ (
    .A(sel_B_11_bF$buf2),
    .B(_558_),
    .Y(_559_)
);

NAND3X1 _1257_ (
    .A(_480_),
    .B(_557_),
    .C(_559_),
    .Y(_560_)
);

INVX1 _1258_ (
    .A(DATA_B[30]),
    .Y(_561_)
);

NAND2X1 _1259_ (
    .A(sel_B_11_bF$buf1),
    .B(_561_),
    .Y(_562_)
);

OR2X2 _1260_ (
    .A(sel_B_11_bF$buf0),
    .B(DATA_B[14]),
    .Y(_563_)
);

NAND3X1 _1261_ (
    .A(sel_B[10]),
    .B(_563_),
    .C(_562_),
    .Y(_564_)
);

NAND3X1 _1262_ (
    .A(sel_B[9]),
    .B(_560_),
    .C(_564_),
    .Y(_565_)
);

OR2X2 _1263_ (
    .A(sel_B_11_bF$buf4),
    .B(DATA_B[2]),
    .Y(_566_)
);

INVX1 _1264_ (
    .A(DATA_B[18]),
    .Y(_567_)
);

NAND2X1 _1265_ (
    .A(sel_B_11_bF$buf3),
    .B(_567_),
    .Y(_568_)
);

NAND3X1 _1266_ (
    .A(_480_),
    .B(_566_),
    .C(_568_),
    .Y(_569_)
);

INVX1 _1267_ (
    .A(DATA_B[10]),
    .Y(_570_)
);

NAND2X1 _1268_ (
    .A(sel_B_11_bF$buf2),
    .B(DATA_B[26]),
    .Y(_571_)
);

OAI21X1 _1269_ (
    .A(_570_),
    .B(sel_B_11_bF$buf1),
    .C(_571_),
    .Y(_572_)
);

NAND2X1 _1270_ (
    .A(sel_B[10]),
    .B(_572_),
    .Y(_573_)
);

NAND3X1 _1271_ (
    .A(_479_),
    .B(_569_),
    .C(_573_),
    .Y(_574_)
);

NAND3X1 _1272_ (
    .A(SEL[3]),
    .B(_565_),
    .C(_574_),
    .Y(_575_)
);

AOI21X1 _1273_ (
    .A(_556_),
    .B(_575_),
    .C(_614_),
    .Y(_478_[2])
);

OR2X2 _1274_ (
    .A(sel_A_11_bF$buf0),
    .B(DATA_A[3]),
    .Y(_576_)
);

INVX1 _1275_ (
    .A(DATA_A[19]),
    .Y(_577_)
);

NAND2X1 _1276_ (
    .A(sel_A_11_bF$buf4),
    .B(_577_),
    .Y(_578_)
);

NAND3X1 _1277_ (
    .A(_617_),
    .B(_576_),
    .C(_578_),
    .Y(_579_)
);

INVX1 _1278_ (
    .A(DATA_A[27]),
    .Y(_580_)
);

NAND2X1 _1279_ (
    .A(sel_A_11_bF$buf3),
    .B(_580_),
    .Y(_581_)
);

OR2X2 _1280_ (
    .A(sel_A_11_bF$buf2),
    .B(DATA_A[11]),
    .Y(_582_)
);

NAND3X1 _1281_ (
    .A(sel_A[10]),
    .B(_582_),
    .C(_581_),
    .Y(_583_)
);

NAND3X1 _1282_ (
    .A(_616_),
    .B(_579_),
    .C(_583_),
    .Y(_584_)
);

OR2X2 _1283_ (
    .A(sel_A_11_bF$buf1),
    .B(DATA_A[7]),
    .Y(_585_)
);

INVX1 _1284_ (
    .A(DATA_A[23]),
    .Y(_586_)
);

NAND2X1 _1285_ (
    .A(sel_A_11_bF$buf0),
    .B(_586_),
    .Y(_587_)
);

NAND3X1 _1286_ (
    .A(_617_),
    .B(_585_),
    .C(_587_),
    .Y(_588_)
);

INVX1 _1287_ (
    .A(DATA_A[15]),
    .Y(_589_)
);

NAND2X1 _1288_ (
    .A(sel_A_11_bF$buf4),
    .B(DATA_A[31]),
    .Y(_590_)
);

OAI21X1 _1289_ (
    .A(_589_),
    .B(sel_A_11_bF$buf3),
    .C(_590_),
    .Y(_591_)
);

NAND2X1 _1290_ (
    .A(sel_A[10]),
    .B(_591_),
    .Y(_592_)
);

NAND3X1 _1291_ (
    .A(sel_A[9]),
    .B(_588_),
    .C(_592_),
    .Y(_593_)
);

NAND3X1 _1292_ (
    .A(_615_),
    .B(_584_),
    .C(_593_),
    .Y(_594_)
);

OR2X2 _1293_ (
    .A(sel_B_11_bF$buf0),
    .B(DATA_B[3]),
    .Y(_595_)
);

INVX1 _1294_ (
    .A(DATA_B[19]),
    .Y(_596_)
);

NAND2X1 _1295_ (
    .A(sel_B_11_bF$buf4),
    .B(_596_),
    .Y(_597_)
);

NAND3X1 _1296_ (
    .A(_480_),
    .B(_595_),
    .C(_597_),
    .Y(_598_)
);

INVX1 _1297_ (
    .A(DATA_B[27]),
    .Y(_599_)
);

NAND2X1 _1298_ (
    .A(sel_B_11_bF$buf3),
    .B(_599_),
    .Y(_600_)
);

OR2X2 _1299_ (
    .A(sel_B_11_bF$buf2),
    .B(DATA_B[11]),
    .Y(_601_)
);

NAND3X1 _1300_ (
    .A(sel_B[10]),
    .B(_601_),
    .C(_600_),
    .Y(_602_)
);

NAND3X1 _1301_ (
    .A(_479_),
    .B(_598_),
    .C(_602_),
    .Y(_603_)
);

OR2X2 _1302_ (
    .A(sel_B_11_bF$buf1),
    .B(DATA_B[7]),
    .Y(_604_)
);

INVX1 _1303_ (
    .A(DATA_B[23]),
    .Y(_605_)
);

NAND2X1 _1304_ (
    .A(sel_B_11_bF$buf0),
    .B(_605_),
    .Y(_606_)
);

NAND3X1 _1305_ (
    .A(_480_),
    .B(_604_),
    .C(_606_),
    .Y(_607_)
);

INVX1 _1306_ (
    .A(DATA_B[15]),
    .Y(_608_)
);

NAND2X1 _1307_ (
    .A(sel_B_11_bF$buf4),
    .B(DATA_B[31]),
    .Y(_609_)
);

OAI21X1 _1308_ (
    .A(_608_),
    .B(sel_B_11_bF$buf3),
    .C(_609_),
    .Y(_610_)
);

NAND2X1 _1309_ (
    .A(sel_B[10]),
    .B(_610_),
    .Y(_611_)
);

NAND3X1 _1310_ (
    .A(sel_B[9]),
    .B(_607_),
    .C(_611_),
    .Y(_612_)
);

NAND3X1 _1311_ (
    .A(SEL[3]),
    .B(_603_),
    .C(_612_),
    .Y(_613_)
);

AOI21X1 _1312_ (
    .A(_594_),
    .B(_613_),
    .C(_614_),
    .Y(_478_[3])
);

DFFPOSX1 _1313_ (
    .CLK(CLK),
    .D(_478_[0]),
    .Q(_0_[12])
);

DFFPOSX1 _1314_ (
    .CLK(CLK),
    .D(_478_[1]),
    .Q(_0_[13])
);

DFFPOSX1 _1315_ (
    .CLK(CLK),
    .D(_478_[2]),
    .Q(_0_[14])
);

DFFPOSX1 _1316_ (
    .CLK(CLK),
    .D(_478_[3]),
    .Q(_0_[15])
);

BUFX2 _637_ (
    .A(_0_[0]),
    .Y(NIBBLE_OUT[0])
);

BUFX2 _638_ (
    .A(_0_[1]),
    .Y(NIBBLE_OUT[1])
);

BUFX2 _639_ (
    .A(_0_[2]),
    .Y(NIBBLE_OUT[2])
);

BUFX2 _640_ (
    .A(_0_[3]),
    .Y(NIBBLE_OUT[3])
);

BUFX2 _641_ (
    .A(_0_[4]),
    .Y(NIBBLE_OUT[4])
);

BUFX2 _642_ (
    .A(_0_[5]),
    .Y(NIBBLE_OUT[5])
);

BUFX2 _643_ (
    .A(_0_[6]),
    .Y(NIBBLE_OUT[6])
);

BUFX2 _644_ (
    .A(_0_[7]),
    .Y(NIBBLE_OUT[7])
);

BUFX2 _645_ (
    .A(_0_[8]),
    .Y(NIBBLE_OUT[8])
);

BUFX2 _646_ (
    .A(_0_[9]),
    .Y(NIBBLE_OUT[9])
);

BUFX2 _647_ (
    .A(_0_[10]),
    .Y(NIBBLE_OUT[10])
);

BUFX2 _648_ (
    .A(_0_[11]),
    .Y(NIBBLE_OUT[11])
);

BUFX2 _649_ (
    .A(_0_[12]),
    .Y(NIBBLE_OUT[12])
);

BUFX2 _650_ (
    .A(_0_[13]),
    .Y(NIBBLE_OUT[13])
);

BUFX2 _651_ (
    .A(_0_[14]),
    .Y(NIBBLE_OUT[14])
);

BUFX2 _652_ (
    .A(_0_[15]),
    .Y(NIBBLE_OUT[15])
);

INVX2 _653_ (
    .A(RESET_L),
    .Y(_137_)
);

INVX2 _654_ (
    .A(SEL[0]),
    .Y(_138_)
);

INVX2 _655_ (
    .A(sel_A[0]),
    .Y(_139_)
);

INVX4 _656_ (
    .A(sel_A[1]),
    .Y(_140_)
);

OR2X2 _657_ (
    .A(DATA_A[0]),
    .B(sel_A_2_bF$buf4),
    .Y(_141_)
);

INVX1 _658_ (
    .A(DATA_A[16]),
    .Y(_142_)
);

NAND2X1 _659_ (
    .A(sel_A_2_bF$buf3),
    .B(_142_),
    .Y(_143_)
);

NAND3X1 _660_ (
    .A(_140_),
    .B(_141_),
    .C(_143_),
    .Y(_144_)
);

INVX1 _661_ (
    .A(DATA_A[24]),
    .Y(_145_)
);

NAND2X1 _662_ (
    .A(sel_A_2_bF$buf2),
    .B(_145_),
    .Y(_146_)
);

OR2X2 _663_ (
    .A(sel_A_2_bF$buf1),
    .B(DATA_A[8]),
    .Y(_147_)
);

NAND3X1 _664_ (
    .A(sel_A[1]),
    .B(_147_),
    .C(_146_),
    .Y(_148_)
);

NAND3X1 _665_ (
    .A(_139_),
    .B(_144_),
    .C(_148_),
    .Y(_149_)
);

OR2X2 _666_ (
    .A(sel_A_2_bF$buf0),
    .B(DATA_A[4]),
    .Y(_150_)
);

INVX1 _667_ (
    .A(DATA_A[20]),
    .Y(_151_)
);

NAND2X1 _668_ (
    .A(sel_A_2_bF$buf4),
    .B(_151_),
    .Y(_152_)
);

NAND3X1 _669_ (
    .A(_140_),
    .B(_150_),
    .C(_152_),
    .Y(_153_)
);

INVX1 _670_ (
    .A(DATA_A[12]),
    .Y(_154_)
);

NAND2X1 _671_ (
    .A(sel_A_2_bF$buf3),
    .B(DATA_A[28]),
    .Y(_155_)
);

OAI21X1 _672_ (
    .A(_154_),
    .B(sel_A_2_bF$buf2),
    .C(_155_),
    .Y(_156_)
);

NAND2X1 _673_ (
    .A(sel_A[1]),
    .B(_156_),
    .Y(_157_)
);

NAND3X1 _674_ (
    .A(sel_A[0]),
    .B(_153_),
    .C(_157_),
    .Y(_158_)
);

NAND3X1 _675_ (
    .A(_138_),
    .B(_149_),
    .C(_158_),
    .Y(_159_)
);

INVX2 _676_ (
    .A(sel_B[0]),
    .Y(_2_)
);

INVX4 _677_ (
    .A(sel_B[1]),
    .Y(_3_)
);

OR2X2 _678_ (
    .A(DATA_B[0]),
    .B(sel_B_2_bF$buf4),
    .Y(_4_)
);

INVX1 _679_ (
    .A(DATA_B[16]),
    .Y(_5_)
);

NAND2X1 _680_ (
    .A(sel_B_2_bF$buf3),
    .B(_5_),
    .Y(_6_)
);

NAND3X1 _681_ (
    .A(_3_),
    .B(_4_),
    .C(_6_),
    .Y(_7_)
);

INVX1 _682_ (
    .A(DATA_B[24]),
    .Y(_8_)
);

NAND2X1 _683_ (
    .A(sel_B_2_bF$buf2),
    .B(_8_),
    .Y(_9_)
);

OR2X2 _684_ (
    .A(sel_B_2_bF$buf1),
    .B(DATA_B[8]),
    .Y(_10_)
);

NAND3X1 _685_ (
    .A(sel_B[1]),
    .B(_10_),
    .C(_9_),
    .Y(_11_)
);

NAND3X1 _686_ (
    .A(_2_),
    .B(_7_),
    .C(_11_),
    .Y(_12_)
);

OR2X2 _687_ (
    .A(sel_B_2_bF$buf0),
    .B(DATA_B[4]),
    .Y(_13_)
);

INVX1 _688_ (
    .A(DATA_B[20]),
    .Y(_14_)
);

NAND2X1 _689_ (
    .A(sel_B_2_bF$buf4),
    .B(_14_),
    .Y(_15_)
);

NAND3X1 _690_ (
    .A(_3_),
    .B(_13_),
    .C(_15_),
    .Y(_16_)
);

INVX1 _691_ (
    .A(DATA_B[12]),
    .Y(_17_)
);

NAND2X1 _692_ (
    .A(sel_B_2_bF$buf3),
    .B(DATA_B[28]),
    .Y(_18_)
);

OAI21X1 _693_ (
    .A(_17_),
    .B(sel_B_2_bF$buf2),
    .C(_18_),
    .Y(_19_)
);

NAND2X1 _694_ (
    .A(sel_B[1]),
    .B(_19_),
    .Y(_20_)
);

NAND3X1 _695_ (
    .A(sel_B[0]),
    .B(_16_),
    .C(_20_),
    .Y(_21_)
);

NAND3X1 _696_ (
    .A(SEL[0]),
    .B(_12_),
    .C(_21_),
    .Y(_22_)
);

AOI21X1 _697_ (
    .A(_159_),
    .B(_22_),
    .C(_137_),
    .Y(_1_[0])
);

OR2X2 _698_ (
    .A(sel_A_2_bF$buf1),
    .B(DATA_A[1]),
    .Y(_23_)
);

INVX1 _699_ (
    .A(DATA_A[17]),
    .Y(_24_)
);

NAND2X1 _700_ (
    .A(sel_A_2_bF$buf0),
    .B(_24_),
    .Y(_25_)
);

NAND3X1 _701_ (
    .A(_140_),
    .B(_23_),
    .C(_25_),
    .Y(_26_)
);

INVX1 _702_ (
    .A(DATA_A[25]),
    .Y(_27_)
);

NAND2X1 _703_ (
    .A(sel_A_2_bF$buf4),
    .B(_27_),
    .Y(_28_)
);

OR2X2 _704_ (
    .A(sel_A_2_bF$buf3),
    .B(DATA_A[9]),
    .Y(_29_)
);

NAND3X1 _705_ (
    .A(sel_A[1]),
    .B(_29_),
    .C(_28_),
    .Y(_30_)
);

NAND3X1 _706_ (
    .A(_139_),
    .B(_26_),
    .C(_30_),
    .Y(_31_)
);

OR2X2 _707_ (
    .A(sel_A_2_bF$buf2),
    .B(DATA_A[5]),
    .Y(_32_)
);

INVX1 _708_ (
    .A(DATA_A[21]),
    .Y(_33_)
);

NAND2X1 _709_ (
    .A(sel_A_2_bF$buf1),
    .B(_33_),
    .Y(_34_)
);

NAND3X1 _710_ (
    .A(_140_),
    .B(_32_),
    .C(_34_),
    .Y(_35_)
);

INVX1 _711_ (
    .A(DATA_A[13]),
    .Y(_36_)
);

NAND2X1 _712_ (
    .A(sel_A_2_bF$buf0),
    .B(DATA_A[29]),
    .Y(_37_)
);

OAI21X1 _713_ (
    .A(_36_),
    .B(sel_A_2_bF$buf4),
    .C(_37_),
    .Y(_38_)
);

NAND2X1 _714_ (
    .A(sel_A[1]),
    .B(_38_),
    .Y(_39_)
);

NAND3X1 _715_ (
    .A(sel_A[0]),
    .B(_35_),
    .C(_39_),
    .Y(_40_)
);

NAND3X1 _716_ (
    .A(_138_),
    .B(_31_),
    .C(_40_),
    .Y(_41_)
);

OR2X2 _717_ (
    .A(sel_B_2_bF$buf1),
    .B(DATA_B[1]),
    .Y(_42_)
);

INVX1 _718_ (
    .A(DATA_B[17]),
    .Y(_43_)
);

NAND2X1 _719_ (
    .A(sel_B_2_bF$buf0),
    .B(_43_),
    .Y(_44_)
);

NAND3X1 _720_ (
    .A(_3_),
    .B(_42_),
    .C(_44_),
    .Y(_45_)
);

INVX1 _721_ (
    .A(DATA_B[25]),
    .Y(_46_)
);

NAND2X1 _722_ (
    .A(sel_B_2_bF$buf4),
    .B(_46_),
    .Y(_47_)
);

OR2X2 _723_ (
    .A(sel_B_2_bF$buf3),
    .B(DATA_B[9]),
    .Y(_48_)
);

NAND3X1 _724_ (
    .A(sel_B[1]),
    .B(_48_),
    .C(_47_),
    .Y(_49_)
);

NAND3X1 _725_ (
    .A(_2_),
    .B(_45_),
    .C(_49_),
    .Y(_50_)
);

OR2X2 _726_ (
    .A(sel_B_2_bF$buf2),
    .B(DATA_B[5]),
    .Y(_51_)
);

INVX1 _727_ (
    .A(DATA_B[21]),
    .Y(_52_)
);

NAND2X1 _728_ (
    .A(sel_B_2_bF$buf1),
    .B(_52_),
    .Y(_53_)
);

NAND3X1 _729_ (
    .A(_3_),
    .B(_51_),
    .C(_53_),
    .Y(_54_)
);

INVX1 _730_ (
    .A(DATA_B[13]),
    .Y(_55_)
);

NAND2X1 _731_ (
    .A(sel_B_2_bF$buf0),
    .B(DATA_B[29]),
    .Y(_56_)
);

OAI21X1 _732_ (
    .A(_55_),
    .B(sel_B_2_bF$buf4),
    .C(_56_),
    .Y(_57_)
);

NAND2X1 _733_ (
    .A(sel_B[1]),
    .B(_57_),
    .Y(_58_)
);

NAND3X1 _734_ (
    .A(sel_B[0]),
    .B(_54_),
    .C(_58_),
    .Y(_59_)
);

NAND3X1 _735_ (
    .A(SEL[0]),
    .B(_50_),
    .C(_59_),
    .Y(_60_)
);

AOI21X1 _736_ (
    .A(_41_),
    .B(_60_),
    .C(_137_),
    .Y(_1_[1])
);

OR2X2 _737_ (
    .A(sel_A_2_bF$buf3),
    .B(DATA_A[2]),
    .Y(_61_)
);

INVX1 _738_ (
    .A(DATA_A[18]),
    .Y(_62_)
);

NAND2X1 _739_ (
    .A(sel_A_2_bF$buf2),
    .B(_62_),
    .Y(_63_)
);

NAND3X1 _740_ (
    .A(_140_),
    .B(_61_),
    .C(_63_),
    .Y(_64_)
);

INVX1 _741_ (
    .A(DATA_A[26]),
    .Y(_65_)
);

NAND2X1 _742_ (
    .A(sel_A_2_bF$buf1),
    .B(_65_),
    .Y(_66_)
);

OR2X2 _743_ (
    .A(sel_A_2_bF$buf0),
    .B(DATA_A[10]),
    .Y(_67_)
);

NAND3X1 _744_ (
    .A(sel_A[1]),
    .B(_67_),
    .C(_66_),
    .Y(_68_)
);

NAND3X1 _745_ (
    .A(_139_),
    .B(_64_),
    .C(_68_),
    .Y(_69_)
);

OR2X2 _746_ (
    .A(sel_A_2_bF$buf4),
    .B(DATA_A[6]),
    .Y(_70_)
);

INVX1 _747_ (
    .A(DATA_A[22]),
    .Y(_71_)
);

NAND2X1 _748_ (
    .A(sel_A_2_bF$buf3),
    .B(_71_),
    .Y(_72_)
);

NAND3X1 _749_ (
    .A(_140_),
    .B(_70_),
    .C(_72_),
    .Y(_73_)
);

INVX1 _750_ (
    .A(DATA_A[14]),
    .Y(_74_)
);

NAND2X1 _751_ (
    .A(sel_A_2_bF$buf2),
    .B(DATA_A[30]),
    .Y(_75_)
);

OAI21X1 _752_ (
    .A(_74_),
    .B(sel_A_2_bF$buf1),
    .C(_75_),
    .Y(_76_)
);

NAND2X1 _753_ (
    .A(sel_A[1]),
    .B(_76_),
    .Y(_77_)
);

NAND3X1 _754_ (
    .A(sel_A[0]),
    .B(_73_),
    .C(_77_),
    .Y(_78_)
);

NAND3X1 _755_ (
    .A(_138_),
    .B(_69_),
    .C(_78_),
    .Y(_79_)
);

OR2X2 _756_ (
    .A(sel_B_2_bF$buf3),
    .B(DATA_B[6]),
    .Y(_80_)
);

INVX1 _757_ (
    .A(DATA_B[22]),
    .Y(_81_)
);

NAND2X1 _758_ (
    .A(sel_B_2_bF$buf2),
    .B(_81_),
    .Y(_82_)
);

NAND3X1 _759_ (
    .A(_3_),
    .B(_80_),
    .C(_82_),
    .Y(_83_)
);

INVX1 _760_ (
    .A(DATA_B[30]),
    .Y(_84_)
);

NAND2X1 _761_ (
    .A(sel_B_2_bF$buf1),
    .B(_84_),
    .Y(_85_)
);

OR2X2 _762_ (
    .A(sel_B_2_bF$buf0),
    .B(DATA_B[14]),
    .Y(_86_)
);

NAND3X1 _763_ (
    .A(sel_B[1]),
    .B(_86_),
    .C(_85_),
    .Y(_87_)
);

NAND3X1 _764_ (
    .A(sel_B[0]),
    .B(_83_),
    .C(_87_),
    .Y(_88_)
);

OR2X2 _765_ (
    .A(sel_B_2_bF$buf4),
    .B(DATA_B[2]),
    .Y(_89_)
);

INVX1 _766_ (
    .A(DATA_B[18]),
    .Y(_90_)
);

NAND2X1 _767_ (
    .A(sel_B_2_bF$buf3),
    .B(_90_),
    .Y(_91_)
);

NAND3X1 _768_ (
    .A(_3_),
    .B(_89_),
    .C(_91_),
    .Y(_92_)
);

INVX1 _769_ (
    .A(DATA_B[10]),
    .Y(_93_)
);

NAND2X1 _770_ (
    .A(sel_B_2_bF$buf2),
    .B(DATA_B[26]),
    .Y(_94_)
);

OAI21X1 _771_ (
    .A(_93_),
    .B(sel_B_2_bF$buf1),
    .C(_94_),
    .Y(_95_)
);

NAND2X1 _772_ (
    .A(sel_B[1]),
    .B(_95_),
    .Y(_96_)
);

NAND3X1 _773_ (
    .A(_2_),
    .B(_92_),
    .C(_96_),
    .Y(_97_)
);

NAND3X1 _774_ (
    .A(SEL[0]),
    .B(_88_),
    .C(_97_),
    .Y(_98_)
);

AOI21X1 _775_ (
    .A(_79_),
    .B(_98_),
    .C(_137_),
    .Y(_1_[2])
);

OR2X2 _776_ (
    .A(sel_A_2_bF$buf0),
    .B(DATA_A[3]),
    .Y(_99_)
);

INVX1 _777_ (
    .A(DATA_A[19]),
    .Y(_100_)
);

NAND2X1 _778_ (
    .A(sel_A_2_bF$buf4),
    .B(_100_),
    .Y(_101_)
);

NAND3X1 _779_ (
    .A(_140_),
    .B(_99_),
    .C(_101_),
    .Y(_102_)
);

INVX1 _780_ (
    .A(DATA_A[27]),
    .Y(_103_)
);

NAND2X1 _781_ (
    .A(sel_A_2_bF$buf3),
    .B(_103_),
    .Y(_104_)
);

OR2X2 _782_ (
    .A(sel_A_2_bF$buf2),
    .B(DATA_A[11]),
    .Y(_105_)
);

NAND3X1 _783_ (
    .A(sel_A[1]),
    .B(_105_),
    .C(_104_),
    .Y(_106_)
);

NAND3X1 _784_ (
    .A(_139_),
    .B(_102_),
    .C(_106_),
    .Y(_107_)
);

OR2X2 _785_ (
    .A(sel_A_2_bF$buf1),
    .B(DATA_A[7]),
    .Y(_108_)
);

INVX1 _786_ (
    .A(DATA_A[23]),
    .Y(_109_)
);

NAND2X1 _787_ (
    .A(sel_A_2_bF$buf0),
    .B(_109_),
    .Y(_110_)
);

NAND3X1 _788_ (
    .A(_140_),
    .B(_108_),
    .C(_110_),
    .Y(_111_)
);

INVX1 _789_ (
    .A(DATA_A[15]),
    .Y(_112_)
);

NAND2X1 _790_ (
    .A(sel_A_2_bF$buf4),
    .B(DATA_A[31]),
    .Y(_113_)
);

OAI21X1 _791_ (
    .A(_112_),
    .B(sel_A_2_bF$buf3),
    .C(_113_),
    .Y(_114_)
);

NAND2X1 _792_ (
    .A(sel_A[1]),
    .B(_114_),
    .Y(_115_)
);

NAND3X1 _793_ (
    .A(sel_A[0]),
    .B(_111_),
    .C(_115_),
    .Y(_116_)
);

NAND3X1 _794_ (
    .A(_138_),
    .B(_107_),
    .C(_116_),
    .Y(_117_)
);

OR2X2 _795_ (
    .A(sel_B_2_bF$buf0),
    .B(DATA_B[3]),
    .Y(_118_)
);

INVX1 _796_ (
    .A(DATA_B[19]),
    .Y(_119_)
);

NAND2X1 _797_ (
    .A(sel_B_2_bF$buf4),
    .B(_119_),
    .Y(_120_)
);

NAND3X1 _798_ (
    .A(_3_),
    .B(_118_),
    .C(_120_),
    .Y(_121_)
);

INVX1 _799_ (
    .A(DATA_B[27]),
    .Y(_122_)
);

NAND2X1 _800_ (
    .A(sel_B_2_bF$buf3),
    .B(_122_),
    .Y(_123_)
);

OR2X2 _801_ (
    .A(sel_B_2_bF$buf2),
    .B(DATA_B[11]),
    .Y(_124_)
);

NAND3X1 _802_ (
    .A(sel_B[1]),
    .B(_124_),
    .C(_123_),
    .Y(_125_)
);

NAND3X1 _803_ (
    .A(_2_),
    .B(_121_),
    .C(_125_),
    .Y(_126_)
);

OR2X2 _804_ (
    .A(sel_B_2_bF$buf1),
    .B(DATA_B[7]),
    .Y(_127_)
);

INVX1 _805_ (
    .A(DATA_B[23]),
    .Y(_128_)
);

NAND2X1 _806_ (
    .A(sel_B_2_bF$buf0),
    .B(_128_),
    .Y(_129_)
);

NAND3X1 _807_ (
    .A(_3_),
    .B(_127_),
    .C(_129_),
    .Y(_130_)
);

INVX1 _808_ (
    .A(DATA_B[15]),
    .Y(_131_)
);

NAND2X1 _809_ (
    .A(sel_B_2_bF$buf4),
    .B(DATA_B[31]),
    .Y(_132_)
);

OAI21X1 _810_ (
    .A(_131_),
    .B(sel_B_2_bF$buf3),
    .C(_132_),
    .Y(_133_)
);

NAND2X1 _811_ (
    .A(sel_B[1]),
    .B(_133_),
    .Y(_134_)
);

NAND3X1 _812_ (
    .A(sel_B[0]),
    .B(_130_),
    .C(_134_),
    .Y(_135_)
);

NAND3X1 _813_ (
    .A(SEL[0]),
    .B(_126_),
    .C(_135_),
    .Y(_136_)
);

AOI21X1 _814_ (
    .A(_117_),
    .B(_136_),
    .C(_137_),
    .Y(_1_[3])
);

DFFPOSX1 _815_ (
    .CLK(CLK),
    .D(_1_[0]),
    .Q(_0_[0])
);

DFFPOSX1 _816_ (
    .CLK(CLK),
    .D(_1_[1]),
    .Q(_0_[1])
);

DFFPOSX1 _817_ (
    .CLK(CLK),
    .D(_1_[2]),
    .Q(_0_[2])
);

DFFPOSX1 _818_ (
    .CLK(CLK),
    .D(_1_[3]),
    .Q(_0_[3])
);

INVX2 _819_ (
    .A(RESET_L),
    .Y(_296_)
);

INVX2 _820_ (
    .A(SEL[1]),
    .Y(_297_)
);

INVX2 _821_ (
    .A(sel_A[3]),
    .Y(_298_)
);

INVX4 _822_ (
    .A(sel_A[4]),
    .Y(_299_)
);

OR2X2 _823_ (
    .A(DATA_A[0]),
    .B(sel_A_5_bF$buf4),
    .Y(_300_)
);

INVX1 _824_ (
    .A(DATA_A[16]),
    .Y(_301_)
);

NAND2X1 _825_ (
    .A(sel_A_5_bF$buf3),
    .B(_301_),
    .Y(_302_)
);

NAND3X1 _826_ (
    .A(_299_),
    .B(_300_),
    .C(_302_),
    .Y(_303_)
);

INVX1 _827_ (
    .A(DATA_A[24]),
    .Y(_304_)
);

NAND2X1 _828_ (
    .A(sel_A_5_bF$buf2),
    .B(_304_),
    .Y(_305_)
);

OR2X2 _829_ (
    .A(sel_A_5_bF$buf1),
    .B(DATA_A[8]),
    .Y(_306_)
);

NAND3X1 _830_ (
    .A(sel_A[4]),
    .B(_306_),
    .C(_305_),
    .Y(_307_)
);

NAND3X1 _831_ (
    .A(_298_),
    .B(_303_),
    .C(_307_),
    .Y(_308_)
);

OR2X2 _832_ (
    .A(sel_A_5_bF$buf0),
    .B(DATA_A[4]),
    .Y(_309_)
);

INVX1 _833_ (
    .A(DATA_A[20]),
    .Y(_310_)
);

NAND2X1 _834_ (
    .A(sel_A_5_bF$buf4),
    .B(_310_),
    .Y(_311_)
);

NAND3X1 _835_ (
    .A(_299_),
    .B(_309_),
    .C(_311_),
    .Y(_312_)
);

INVX1 _836_ (
    .A(DATA_A[12]),
    .Y(_313_)
);

NAND2X1 _837_ (
    .A(sel_A_5_bF$buf3),
    .B(DATA_A[28]),
    .Y(_314_)
);

OAI21X1 _838_ (
    .A(_313_),
    .B(sel_A_5_bF$buf2),
    .C(_314_),
    .Y(_315_)
);

NAND2X1 _839_ (
    .A(sel_A[4]),
    .B(_315_),
    .Y(_316_)
);

NAND3X1 _840_ (
    .A(sel_A[3]),
    .B(_312_),
    .C(_316_),
    .Y(_317_)
);

NAND3X1 _841_ (
    .A(_297_),
    .B(_308_),
    .C(_317_),
    .Y(_318_)
);

INVX2 _842_ (
    .A(sel_B[3]),
    .Y(_161_)
);

INVX4 _843_ (
    .A(sel_B[4]),
    .Y(_162_)
);

OR2X2 _844_ (
    .A(DATA_B[0]),
    .B(sel_B_5_bF$buf4),
    .Y(_163_)
);

INVX1 _845_ (
    .A(DATA_B[16]),
    .Y(_164_)
);

NAND2X1 _846_ (
    .A(sel_B_5_bF$buf3),
    .B(_164_),
    .Y(_165_)
);

NAND3X1 _847_ (
    .A(_162_),
    .B(_163_),
    .C(_165_),
    .Y(_166_)
);

INVX1 _848_ (
    .A(DATA_B[24]),
    .Y(_167_)
);

NAND2X1 _849_ (
    .A(sel_B_5_bF$buf2),
    .B(_167_),
    .Y(_168_)
);

OR2X2 _850_ (
    .A(sel_B_5_bF$buf1),
    .B(DATA_B[8]),
    .Y(_169_)
);

NAND3X1 _851_ (
    .A(sel_B[4]),
    .B(_169_),
    .C(_168_),
    .Y(_170_)
);

NAND3X1 _852_ (
    .A(_161_),
    .B(_166_),
    .C(_170_),
    .Y(_171_)
);

OR2X2 _853_ (
    .A(sel_B_5_bF$buf0),
    .B(DATA_B[4]),
    .Y(_172_)
);

INVX1 _854_ (
    .A(DATA_B[20]),
    .Y(_173_)
);

NAND2X1 _855_ (
    .A(sel_B_5_bF$buf4),
    .B(_173_),
    .Y(_174_)
);

NAND3X1 _856_ (
    .A(_162_),
    .B(_172_),
    .C(_174_),
    .Y(_175_)
);

INVX1 _857_ (
    .A(DATA_B[12]),
    .Y(_176_)
);

NAND2X1 _858_ (
    .A(sel_B_5_bF$buf3),
    .B(DATA_B[28]),
    .Y(_177_)
);

OAI21X1 _859_ (
    .A(_176_),
    .B(sel_B_5_bF$buf2),
    .C(_177_),
    .Y(_178_)
);

NAND2X1 _860_ (
    .A(sel_B[4]),
    .B(_178_),
    .Y(_179_)
);

NAND3X1 _861_ (
    .A(sel_B[3]),
    .B(_175_),
    .C(_179_),
    .Y(_180_)
);

NAND3X1 _862_ (
    .A(SEL[1]),
    .B(_171_),
    .C(_180_),
    .Y(_181_)
);

AOI21X1 _863_ (
    .A(_318_),
    .B(_181_),
    .C(_296_),
    .Y(_160_[0])
);

OR2X2 _864_ (
    .A(sel_A_5_bF$buf1),
    .B(DATA_A[1]),
    .Y(_182_)
);

INVX1 _865_ (
    .A(DATA_A[17]),
    .Y(_183_)
);

NAND2X1 _866_ (
    .A(sel_A_5_bF$buf0),
    .B(_183_),
    .Y(_184_)
);

NAND3X1 _867_ (
    .A(_299_),
    .B(_182_),
    .C(_184_),
    .Y(_185_)
);

INVX1 _868_ (
    .A(DATA_A[25]),
    .Y(_186_)
);

NAND2X1 _869_ (
    .A(sel_A_5_bF$buf4),
    .B(_186_),
    .Y(_187_)
);

OR2X2 _870_ (
    .A(sel_A_5_bF$buf3),
    .B(DATA_A[9]),
    .Y(_188_)
);

NAND3X1 _871_ (
    .A(sel_A[4]),
    .B(_188_),
    .C(_187_),
    .Y(_189_)
);

NAND3X1 _872_ (
    .A(_298_),
    .B(_185_),
    .C(_189_),
    .Y(_190_)
);

OR2X2 _873_ (
    .A(sel_A_5_bF$buf2),
    .B(DATA_A[5]),
    .Y(_191_)
);

INVX1 _874_ (
    .A(DATA_A[21]),
    .Y(_192_)
);

NAND2X1 _875_ (
    .A(sel_A_5_bF$buf1),
    .B(_192_),
    .Y(_193_)
);

NAND3X1 _876_ (
    .A(_299_),
    .B(_191_),
    .C(_193_),
    .Y(_194_)
);

INVX1 _877_ (
    .A(DATA_A[13]),
    .Y(_195_)
);

NAND2X1 _878_ (
    .A(sel_A_5_bF$buf0),
    .B(DATA_A[29]),
    .Y(_196_)
);

OAI21X1 _879_ (
    .A(_195_),
    .B(sel_A_5_bF$buf4),
    .C(_196_),
    .Y(_197_)
);

NAND2X1 _880_ (
    .A(sel_A[4]),
    .B(_197_),
    .Y(_198_)
);

NAND3X1 _881_ (
    .A(sel_A[3]),
    .B(_194_),
    .C(_198_),
    .Y(_199_)
);

NAND3X1 _882_ (
    .A(_297_),
    .B(_190_),
    .C(_199_),
    .Y(_200_)
);

OR2X2 _883_ (
    .A(sel_B_5_bF$buf1),
    .B(DATA_B[1]),
    .Y(_201_)
);

INVX1 _884_ (
    .A(DATA_B[17]),
    .Y(_202_)
);

NAND2X1 _885_ (
    .A(sel_B_5_bF$buf0),
    .B(_202_),
    .Y(_203_)
);

NAND3X1 _886_ (
    .A(_162_),
    .B(_201_),
    .C(_203_),
    .Y(_204_)
);

INVX1 _887_ (
    .A(DATA_B[25]),
    .Y(_205_)
);

NAND2X1 _888_ (
    .A(sel_B_5_bF$buf4),
    .B(_205_),
    .Y(_206_)
);

OR2X2 _889_ (
    .A(sel_B_5_bF$buf3),
    .B(DATA_B[9]),
    .Y(_207_)
);

NAND3X1 _890_ (
    .A(sel_B[4]),
    .B(_207_),
    .C(_206_),
    .Y(_208_)
);

NAND3X1 _891_ (
    .A(_161_),
    .B(_204_),
    .C(_208_),
    .Y(_209_)
);

OR2X2 _892_ (
    .A(sel_B_5_bF$buf2),
    .B(DATA_B[5]),
    .Y(_210_)
);

INVX1 _893_ (
    .A(DATA_B[21]),
    .Y(_211_)
);

NAND2X1 _894_ (
    .A(sel_B_5_bF$buf1),
    .B(_211_),
    .Y(_212_)
);

NAND3X1 _895_ (
    .A(_162_),
    .B(_210_),
    .C(_212_),
    .Y(_213_)
);

INVX1 _896_ (
    .A(DATA_B[13]),
    .Y(_214_)
);

NAND2X1 _897_ (
    .A(sel_B_5_bF$buf0),
    .B(DATA_B[29]),
    .Y(_215_)
);

OAI21X1 _898_ (
    .A(_214_),
    .B(sel_B_5_bF$buf4),
    .C(_215_),
    .Y(_216_)
);

NAND2X1 _899_ (
    .A(sel_B[4]),
    .B(_216_),
    .Y(_217_)
);

NAND3X1 _900_ (
    .A(sel_B[3]),
    .B(_213_),
    .C(_217_),
    .Y(_218_)
);

NAND3X1 _901_ (
    .A(SEL[1]),
    .B(_209_),
    .C(_218_),
    .Y(_219_)
);

AOI21X1 _902_ (
    .A(_200_),
    .B(_219_),
    .C(_296_),
    .Y(_160_[1])
);

OR2X2 _903_ (
    .A(sel_A_5_bF$buf3),
    .B(DATA_A[2]),
    .Y(_220_)
);

INVX1 _904_ (
    .A(DATA_A[18]),
    .Y(_221_)
);

NAND2X1 _905_ (
    .A(sel_A_5_bF$buf2),
    .B(_221_),
    .Y(_222_)
);

NAND3X1 _906_ (
    .A(_299_),
    .B(_220_),
    .C(_222_),
    .Y(_223_)
);

INVX1 _907_ (
    .A(DATA_A[26]),
    .Y(_224_)
);

NAND2X1 _908_ (
    .A(sel_A_5_bF$buf1),
    .B(_224_),
    .Y(_225_)
);

OR2X2 _909_ (
    .A(sel_A_5_bF$buf0),
    .B(DATA_A[10]),
    .Y(_226_)
);

NAND3X1 _910_ (
    .A(sel_A[4]),
    .B(_226_),
    .C(_225_),
    .Y(_227_)
);

NAND3X1 _911_ (
    .A(_298_),
    .B(_223_),
    .C(_227_),
    .Y(_228_)
);

OR2X2 _912_ (
    .A(sel_A_5_bF$buf4),
    .B(DATA_A[6]),
    .Y(_229_)
);

INVX1 _913_ (
    .A(DATA_A[22]),
    .Y(_230_)
);

NAND2X1 _914_ (
    .A(sel_A_5_bF$buf3),
    .B(_230_),
    .Y(_231_)
);

NAND3X1 _915_ (
    .A(_299_),
    .B(_229_),
    .C(_231_),
    .Y(_232_)
);

INVX1 _916_ (
    .A(DATA_A[14]),
    .Y(_233_)
);

NAND2X1 _917_ (
    .A(sel_A_5_bF$buf2),
    .B(DATA_A[30]),
    .Y(_234_)
);

OAI21X1 _918_ (
    .A(_233_),
    .B(sel_A_5_bF$buf1),
    .C(_234_),
    .Y(_235_)
);

NAND2X1 _919_ (
    .A(sel_A[4]),
    .B(_235_),
    .Y(_236_)
);

NAND3X1 _920_ (
    .A(sel_A[3]),
    .B(_232_),
    .C(_236_),
    .Y(_237_)
);

NAND3X1 _921_ (
    .A(_297_),
    .B(_228_),
    .C(_237_),
    .Y(_238_)
);

OR2X2 _922_ (
    .A(sel_B_5_bF$buf3),
    .B(DATA_B[6]),
    .Y(_239_)
);

INVX1 _923_ (
    .A(DATA_B[22]),
    .Y(_240_)
);

NAND2X1 _924_ (
    .A(sel_B_5_bF$buf2),
    .B(_240_),
    .Y(_241_)
);

NAND3X1 _925_ (
    .A(_162_),
    .B(_239_),
    .C(_241_),
    .Y(_242_)
);

INVX1 _926_ (
    .A(DATA_B[30]),
    .Y(_243_)
);

NAND2X1 _927_ (
    .A(sel_B_5_bF$buf1),
    .B(_243_),
    .Y(_244_)
);

OR2X2 _928_ (
    .A(sel_B_5_bF$buf0),
    .B(DATA_B[14]),
    .Y(_245_)
);

NAND3X1 _929_ (
    .A(sel_B[4]),
    .B(_245_),
    .C(_244_),
    .Y(_246_)
);

NAND3X1 _930_ (
    .A(sel_B[3]),
    .B(_242_),
    .C(_246_),
    .Y(_247_)
);

OR2X2 _931_ (
    .A(sel_B_5_bF$buf4),
    .B(DATA_B[2]),
    .Y(_248_)
);

INVX1 _932_ (
    .A(DATA_B[18]),
    .Y(_249_)
);

NAND2X1 _933_ (
    .A(sel_B_5_bF$buf3),
    .B(_249_),
    .Y(_250_)
);

NAND3X1 _934_ (
    .A(_162_),
    .B(_248_),
    .C(_250_),
    .Y(_251_)
);

INVX1 _935_ (
    .A(DATA_B[10]),
    .Y(_252_)
);

NAND2X1 _936_ (
    .A(sel_B_5_bF$buf2),
    .B(DATA_B[26]),
    .Y(_253_)
);

OAI21X1 _937_ (
    .A(_252_),
    .B(sel_B_5_bF$buf1),
    .C(_253_),
    .Y(_254_)
);

NAND2X1 _938_ (
    .A(sel_B[4]),
    .B(_254_),
    .Y(_255_)
);

NAND3X1 _939_ (
    .A(_161_),
    .B(_251_),
    .C(_255_),
    .Y(_256_)
);

NAND3X1 _940_ (
    .A(SEL[1]),
    .B(_247_),
    .C(_256_),
    .Y(_257_)
);

AOI21X1 _941_ (
    .A(_238_),
    .B(_257_),
    .C(_296_),
    .Y(_160_[2])
);

OR2X2 _942_ (
    .A(sel_A_5_bF$buf0),
    .B(DATA_A[3]),
    .Y(_258_)
);

INVX1 _943_ (
    .A(DATA_A[19]),
    .Y(_259_)
);

NAND2X1 _944_ (
    .A(sel_A_5_bF$buf4),
    .B(_259_),
    .Y(_260_)
);

NAND3X1 _945_ (
    .A(_299_),
    .B(_258_),
    .C(_260_),
    .Y(_261_)
);

INVX1 _946_ (
    .A(DATA_A[27]),
    .Y(_262_)
);

NAND2X1 _947_ (
    .A(sel_A_5_bF$buf3),
    .B(_262_),
    .Y(_263_)
);

OR2X2 _948_ (
    .A(sel_A_5_bF$buf2),
    .B(DATA_A[11]),
    .Y(_264_)
);

NAND3X1 _949_ (
    .A(sel_A[4]),
    .B(_264_),
    .C(_263_),
    .Y(_265_)
);

NAND3X1 _950_ (
    .A(_298_),
    .B(_261_),
    .C(_265_),
    .Y(_266_)
);

OR2X2 _951_ (
    .A(sel_A_5_bF$buf1),
    .B(DATA_A[7]),
    .Y(_267_)
);

INVX1 _952_ (
    .A(DATA_A[23]),
    .Y(_268_)
);

NAND2X1 _953_ (
    .A(sel_A_5_bF$buf0),
    .B(_268_),
    .Y(_269_)
);

NAND3X1 _954_ (
    .A(_299_),
    .B(_267_),
    .C(_269_),
    .Y(_270_)
);

INVX1 _955_ (
    .A(DATA_A[15]),
    .Y(_271_)
);

NAND2X1 _956_ (
    .A(sel_A_5_bF$buf4),
    .B(DATA_A[31]),
    .Y(_272_)
);

OAI21X1 _957_ (
    .A(_271_),
    .B(sel_A_5_bF$buf3),
    .C(_272_),
    .Y(_273_)
);

NAND2X1 _958_ (
    .A(sel_A[4]),
    .B(_273_),
    .Y(_274_)
);

NAND3X1 _959_ (
    .A(sel_A[3]),
    .B(_270_),
    .C(_274_),
    .Y(_275_)
);

NAND3X1 _960_ (
    .A(_297_),
    .B(_266_),
    .C(_275_),
    .Y(_276_)
);

OR2X2 _961_ (
    .A(sel_B_5_bF$buf0),
    .B(DATA_B[3]),
    .Y(_277_)
);

INVX1 _962_ (
    .A(DATA_B[19]),
    .Y(_278_)
);

NAND2X1 _963_ (
    .A(sel_B_5_bF$buf4),
    .B(_278_),
    .Y(_279_)
);

NAND3X1 _964_ (
    .A(_162_),
    .B(_277_),
    .C(_279_),
    .Y(_280_)
);

INVX1 _965_ (
    .A(DATA_B[27]),
    .Y(_281_)
);

NAND2X1 _966_ (
    .A(sel_B_5_bF$buf3),
    .B(_281_),
    .Y(_282_)
);

OR2X2 _967_ (
    .A(sel_B_5_bF$buf2),
    .B(DATA_B[11]),
    .Y(_283_)
);

NAND3X1 _968_ (
    .A(sel_B[4]),
    .B(_283_),
    .C(_282_),
    .Y(_284_)
);

NAND3X1 _969_ (
    .A(_161_),
    .B(_280_),
    .C(_284_),
    .Y(_285_)
);

OR2X2 _970_ (
    .A(sel_B_5_bF$buf1),
    .B(DATA_B[7]),
    .Y(_286_)
);

INVX1 _971_ (
    .A(DATA_B[23]),
    .Y(_287_)
);

NAND2X1 _972_ (
    .A(sel_B_5_bF$buf0),
    .B(_287_),
    .Y(_288_)
);

NAND3X1 _973_ (
    .A(_162_),
    .B(_286_),
    .C(_288_),
    .Y(_289_)
);

INVX1 _974_ (
    .A(DATA_B[15]),
    .Y(_290_)
);

NAND2X1 _975_ (
    .A(sel_B_5_bF$buf4),
    .B(DATA_B[31]),
    .Y(_291_)
);

OAI21X1 _976_ (
    .A(_290_),
    .B(sel_B_5_bF$buf3),
    .C(_291_),
    .Y(_292_)
);

NAND2X1 _977_ (
    .A(sel_B[4]),
    .B(_292_),
    .Y(_293_)
);

NAND3X1 _978_ (
    .A(sel_B[3]),
    .B(_289_),
    .C(_293_),
    .Y(_294_)
);

NAND3X1 _979_ (
    .A(SEL[1]),
    .B(_285_),
    .C(_294_),
    .Y(_295_)
);

AOI21X1 _980_ (
    .A(_276_),
    .B(_295_),
    .C(_296_),
    .Y(_160_[3])
);

DFFPOSX1 _981_ (
    .CLK(CLK),
    .D(_160_[0]),
    .Q(_0_[4])
);

DFFPOSX1 _982_ (
    .CLK(CLK),
    .D(_160_[1]),
    .Q(_0_[5])
);

DFFPOSX1 _983_ (
    .CLK(CLK),
    .D(_160_[2]),
    .Q(_0_[6])
);

DFFPOSX1 _984_ (
    .CLK(CLK),
    .D(_160_[3]),
    .Q(_0_[7])
);

INVX2 _985_ (
    .A(RESET_L),
    .Y(_455_)
);

INVX2 _986_ (
    .A(SEL[2]),
    .Y(_456_)
);

INVX2 _987_ (
    .A(sel_A[6]),
    .Y(_457_)
);

INVX4 _988_ (
    .A(sel_A[7]),
    .Y(_458_)
);

OR2X2 _989_ (
    .A(DATA_A[0]),
    .B(sel_A_8_bF$buf2),
    .Y(_459_)
);

INVX1 _990_ (
    .A(DATA_A[16]),
    .Y(_460_)
);

NAND2X1 _991_ (
    .A(sel_A_8_bF$buf1),
    .B(_460_),
    .Y(_461_)
);

NAND3X1 _992_ (
    .A(_458_),
    .B(_459_),
    .C(_461_),
    .Y(_462_)
);

INVX1 _993_ (
    .A(DATA_A[24]),
    .Y(_463_)
);

NAND2X1 _994_ (
    .A(sel_A_8_bF$buf0),
    .B(_463_),
    .Y(_464_)
);

OR2X2 _995_ (
    .A(sel_A_8_bF$buf4),
    .B(DATA_A[8]),
    .Y(_465_)
);

NAND3X1 _996_ (
    .A(sel_A[7]),
    .B(_465_),
    .C(_464_),
    .Y(_466_)
);

NAND3X1 _997_ (
    .A(_457_),
    .B(_462_),
    .C(_466_),
    .Y(_467_)
);

OR2X2 _998_ (
    .A(sel_A_8_bF$buf3),
    .B(DATA_A[4]),
    .Y(_468_)
);

INVX1 _999_ (
    .A(DATA_A[20]),
    .Y(_469_)
);

endmodule
