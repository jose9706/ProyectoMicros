magic
tech scmos
timestamp 1560018123
<< metal1 >>
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 485 1403 488 1407
rect 286 1368 297 1371
rect 1386 1368 1393 1371
rect 286 1366 290 1368
rect 294 1362 297 1368
rect 14 1358 25 1361
rect 118 1358 129 1361
rect 142 1358 150 1361
rect 158 1358 177 1361
rect 246 1352 249 1361
rect 302 1358 313 1361
rect 214 1348 222 1351
rect 446 1351 449 1361
rect 510 1358 521 1361
rect 446 1348 465 1351
rect 550 1348 558 1351
rect 718 1351 721 1361
rect 814 1358 825 1361
rect 854 1358 865 1361
rect 910 1358 921 1361
rect 966 1358 982 1361
rect 1178 1358 1185 1361
rect 1226 1358 1230 1362
rect 1278 1358 1289 1361
rect 1318 1358 1329 1361
rect 1438 1358 1446 1361
rect 718 1348 737 1351
rect 774 1348 785 1351
rect 974 1348 1006 1351
rect 42 1338 49 1341
rect 98 1338 105 1341
rect 222 1338 233 1341
rect 242 1338 257 1341
rect 266 1338 270 1341
rect 358 1341 361 1348
rect 350 1338 361 1341
rect 378 1338 385 1341
rect 414 1338 425 1341
rect 446 1338 454 1341
rect 470 1338 494 1341
rect 526 1341 529 1348
rect 774 1342 777 1348
rect 526 1338 537 1341
rect 650 1338 657 1341
rect 750 1338 761 1341
rect 790 1338 798 1341
rect 870 1341 873 1348
rect 870 1338 881 1341
rect 942 1338 950 1341
rect 974 1338 977 1348
rect 1022 1338 1025 1348
rect 1170 1338 1177 1341
rect 1342 1338 1358 1341
rect 6 1328 9 1338
rect 46 1328 49 1338
rect 150 1328 153 1338
rect 85 1318 86 1322
rect 282 1318 283 1322
rect 850 1318 851 1322
rect 925 1318 926 1322
rect 1133 1318 1134 1322
rect 1157 1318 1158 1322
rect 1253 1318 1254 1322
rect 1293 1318 1294 1322
rect 1333 1318 1334 1322
rect 1418 1318 1425 1321
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 22 1278 30 1281
rect 34 1268 41 1271
rect 174 1268 182 1271
rect 274 1268 281 1271
rect 326 1268 334 1271
rect 382 1268 393 1271
rect 466 1268 489 1271
rect 510 1268 521 1271
rect 710 1271 713 1278
rect 702 1268 713 1271
rect 750 1271 754 1272
rect 758 1271 761 1278
rect 750 1268 761 1271
rect 1038 1271 1041 1281
rect 1034 1268 1041 1271
rect 1134 1271 1138 1272
rect 1142 1271 1145 1278
rect 1134 1268 1145 1271
rect 306 1258 313 1261
rect 1086 1261 1089 1268
rect 1078 1258 1089 1261
rect 646 1248 657 1251
rect 678 1248 689 1251
rect 906 1248 913 1251
rect 1070 1251 1073 1258
rect 1006 1248 1017 1251
rect 1062 1248 1073 1251
rect 1190 1251 1193 1258
rect 1154 1248 1161 1251
rect 1182 1248 1193 1251
rect 1198 1248 1209 1251
rect 546 1238 553 1241
rect 634 1238 641 1241
rect 1214 1238 1222 1241
rect 822 1228 825 1238
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 485 1203 488 1207
rect 94 1168 102 1171
rect 830 1171 833 1181
rect 1134 1172 1137 1181
rect 830 1168 838 1171
rect 1198 1168 1209 1171
rect 138 1158 145 1161
rect 166 1158 177 1161
rect 214 1158 233 1161
rect 294 1158 305 1161
rect 422 1158 430 1161
rect 654 1161 657 1168
rect 1206 1162 1209 1168
rect 558 1158 569 1161
rect 630 1158 641 1161
rect 646 1158 657 1161
rect 750 1158 761 1161
rect 874 1158 881 1161
rect 974 1158 1009 1161
rect 1046 1158 1057 1161
rect 1158 1158 1169 1161
rect 1374 1158 1385 1161
rect 718 1151 722 1154
rect 718 1148 737 1151
rect 22 1141 25 1148
rect 22 1138 33 1141
rect 246 1138 257 1141
rect 518 1138 529 1141
rect 778 1138 785 1141
rect 1026 1138 1033 1141
rect 1206 1141 1209 1148
rect 1206 1138 1217 1141
rect 1244 1138 1246 1142
rect 182 1128 185 1138
rect 254 1132 257 1138
rect 518 1132 521 1138
rect 470 1128 478 1131
rect 782 1128 785 1138
rect 126 1118 134 1121
rect 237 1118 238 1122
rect 309 1118 310 1122
rect 573 1118 574 1122
rect 765 1118 766 1122
rect 850 1118 852 1122
rect 900 1118 902 1122
rect 1173 1118 1174 1122
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 6 1072 9 1081
rect 38 1068 49 1071
rect 538 1068 545 1071
rect 630 1071 633 1078
rect 630 1068 641 1071
rect 854 1071 857 1078
rect 844 1068 857 1071
rect 1086 1071 1089 1078
rect 1078 1068 1089 1071
rect 1190 1071 1194 1072
rect 1198 1071 1201 1078
rect 1190 1068 1201 1071
rect 222 1058 230 1061
rect 302 1058 313 1061
rect 550 1061 553 1068
rect 550 1058 561 1061
rect 1206 1058 1225 1061
rect 302 1052 305 1058
rect 14 1048 25 1051
rect 130 1048 137 1051
rect 286 1048 297 1051
rect 462 1048 494 1051
rect 654 1048 665 1051
rect 710 1048 718 1051
rect 758 1048 769 1051
rect 974 1048 982 1051
rect 1078 1051 1081 1058
rect 1206 1056 1210 1058
rect 1070 1048 1081 1051
rect 1406 1048 1417 1051
rect 518 1041 521 1048
rect 518 1038 529 1041
rect 742 1041 745 1048
rect 742 1038 753 1041
rect 1246 1038 1262 1041
rect 1422 1038 1430 1041
rect 86 1028 89 1038
rect 246 1028 249 1038
rect 878 1028 881 1038
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 485 1003 488 1007
rect 1190 972 1193 981
rect 98 968 105 971
rect 158 968 174 971
rect 326 968 334 971
rect 1366 971 1369 981
rect 1362 968 1369 971
rect 1394 968 1401 971
rect 94 958 105 961
rect 334 958 345 961
rect 718 958 729 961
rect 914 958 921 961
rect 926 958 937 961
rect 334 952 337 958
rect 1134 952 1137 961
rect 1322 958 1326 961
rect 1406 958 1417 961
rect 794 948 801 951
rect 994 948 1001 951
rect 122 938 129 941
rect 362 938 377 941
rect 902 938 910 941
rect 1034 938 1041 941
rect 1158 938 1169 941
rect 1270 938 1281 941
rect 166 931 169 938
rect 158 928 169 931
rect 766 931 769 938
rect 766 928 777 931
rect 194 918 201 921
rect 306 918 307 922
rect 386 918 387 922
rect 422 918 430 921
rect 454 918 462 921
rect 498 918 500 922
rect 650 918 657 921
rect 674 918 676 922
rect 714 918 715 922
rect 826 918 828 922
rect 1302 918 1310 921
rect 1338 918 1345 921
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 258 888 259 892
rect 738 888 739 892
rect 1181 888 1182 892
rect 1210 888 1211 892
rect 1250 888 1251 892
rect 1274 888 1275 892
rect 1386 888 1387 892
rect 622 878 630 881
rect 1010 878 1017 881
rect 382 868 390 871
rect 838 871 841 878
rect 838 868 849 871
rect 742 861 745 868
rect 742 858 753 861
rect 886 858 894 861
rect 938 858 953 861
rect 974 861 977 871
rect 962 858 977 861
rect 1046 861 1049 871
rect 1034 858 1049 861
rect 1062 868 1073 871
rect 1106 868 1113 871
rect 1134 868 1145 871
rect 1194 868 1201 871
rect 1310 868 1321 871
rect 1422 868 1433 871
rect 1062 862 1065 868
rect 1094 858 1113 861
rect 1390 858 1409 861
rect 1438 858 1457 861
rect 94 848 105 851
rect 542 848 553 851
rect 862 848 873 851
rect 918 848 929 851
rect 974 848 985 851
rect 990 848 998 851
rect 1110 848 1113 858
rect 1214 848 1225 851
rect 1342 848 1361 851
rect 1390 848 1393 858
rect 1438 852 1441 858
rect 102 842 105 848
rect 902 841 905 848
rect 974 842 977 848
rect 1062 842 1066 844
rect 902 838 913 841
rect 278 828 281 838
rect 1330 828 1331 832
rect 472 803 474 807
rect 478 803 481 807
rect 485 803 488 807
rect 750 768 761 771
rect 750 762 753 768
rect 30 751 34 753
rect 22 748 34 751
rect 150 742 153 751
rect 434 738 441 741
rect 470 738 494 741
rect 598 738 601 748
rect 1026 748 1041 751
rect 1094 751 1097 758
rect 1094 748 1105 751
rect 1230 751 1234 753
rect 1230 748 1241 751
rect 1262 742 1265 751
rect 1414 751 1418 753
rect 1414 748 1425 751
rect 770 738 777 741
rect 1086 738 1094 741
rect 154 728 161 731
rect 790 731 793 738
rect 450 728 457 731
rect 782 728 793 731
rect 1066 728 1070 732
rect 634 718 641 721
rect 666 718 673 721
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 474 688 481 691
rect 874 688 876 692
rect 914 688 921 691
rect 946 688 953 691
rect 602 678 609 681
rect 1290 678 1297 681
rect 718 671 721 678
rect 710 668 721 671
rect 1238 671 1242 672
rect 1246 671 1249 678
rect 1238 668 1249 671
rect 1298 668 1305 671
rect 1462 668 1470 671
rect 22 658 34 661
rect 214 658 217 668
rect 266 658 281 661
rect 334 658 346 661
rect 394 658 401 661
rect 454 658 470 661
rect 598 658 601 668
rect 30 657 34 658
rect 342 657 346 658
rect 654 651 657 658
rect 1198 657 1202 658
rect 1102 652 1106 654
rect 646 648 657 651
rect 662 648 673 651
rect 834 648 841 651
rect 894 648 902 651
rect 678 638 686 641
rect 890 638 921 641
rect 1238 638 1246 641
rect 1395 638 1398 642
rect 974 628 977 638
rect 472 603 474 607
rect 478 603 481 607
rect 485 603 488 607
rect 806 572 809 581
rect 942 572 945 581
rect 1222 572 1225 581
rect 470 568 502 571
rect 550 568 558 571
rect 606 568 617 571
rect 630 568 646 571
rect 6 566 10 568
rect 614 562 617 568
rect 70 558 81 561
rect 142 558 153 561
rect 190 558 201 561
rect 222 558 233 561
rect 262 558 273 561
rect 278 558 286 561
rect 410 558 417 561
rect 534 558 545 561
rect 574 558 585 561
rect 590 558 601 561
rect 666 558 673 561
rect 846 558 854 561
rect 894 558 905 561
rect 1230 558 1238 561
rect 1318 558 1329 561
rect 414 551 418 554
rect 582 552 585 558
rect 902 552 906 554
rect 414 548 422 551
rect 22 538 33 541
rect 166 538 174 541
rect 286 538 297 541
rect 438 538 449 541
rect 690 538 697 541
rect 1454 538 1478 541
rect 30 532 33 538
rect 62 528 65 538
rect 206 531 209 538
rect 294 532 297 538
rect 446 532 449 538
rect 206 528 217 531
rect 694 528 697 538
rect 990 528 1006 531
rect 13 518 14 522
rect 186 518 187 522
rect 237 518 238 522
rect 429 518 430 522
rect 677 518 678 522
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 914 488 921 491
rect 946 488 947 492
rect 1162 488 1163 492
rect 1274 488 1275 492
rect 202 478 209 481
rect 994 478 1001 481
rect 14 468 25 471
rect 190 468 198 471
rect 354 468 361 471
rect 534 468 545 471
rect 554 468 561 471
rect 610 468 617 471
rect 746 468 753 471
rect 798 468 809 471
rect 830 468 838 471
rect 878 471 882 472
rect 886 471 889 478
rect 878 468 889 471
rect 1090 468 1092 472
rect 1254 468 1262 471
rect 86 461 89 468
rect 534 462 537 468
rect 78 458 89 461
rect 574 458 593 461
rect 774 458 790 461
rect 810 458 817 461
rect 1018 458 1025 461
rect 1398 458 1418 461
rect 590 448 593 458
rect 894 456 898 458
rect 1414 456 1418 458
rect 718 448 729 451
rect 770 448 774 452
rect 94 438 129 441
rect 358 441 361 448
rect 358 438 369 441
rect 534 441 537 448
rect 526 438 537 441
rect 702 441 705 448
rect 702 438 713 441
rect 894 441 897 451
rect 1054 448 1065 451
rect 1182 448 1193 451
rect 1222 448 1230 451
rect 1290 448 1297 451
rect 894 438 910 441
rect 1078 441 1081 448
rect 1070 438 1081 441
rect 1106 438 1121 441
rect 472 403 474 407
rect 478 403 481 407
rect 485 403 488 407
rect 786 388 787 392
rect 638 372 641 381
rect 158 368 166 371
rect 230 368 265 371
rect 350 368 361 371
rect 922 368 929 371
rect 358 362 361 368
rect 98 358 105 361
rect 270 358 281 361
rect 334 358 345 361
rect 470 358 478 361
rect 30 352 34 354
rect 286 351 289 358
rect 286 348 297 351
rect 494 351 497 361
rect 726 358 737 361
rect 1226 358 1233 361
rect 450 348 457 351
rect 462 348 497 351
rect 982 348 1014 351
rect 1454 348 1465 351
rect 310 338 326 341
rect 438 338 449 341
rect 766 338 777 341
rect 814 338 822 341
rect 894 338 905 341
rect 982 338 985 348
rect 1030 338 1033 348
rect 1454 342 1457 348
rect 1190 338 1201 341
rect 902 332 905 338
rect 1198 332 1201 338
rect 973 318 974 322
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 14 288 22 291
rect 74 288 81 291
rect 122 288 123 292
rect 170 288 177 291
rect 454 288 462 291
rect 482 288 497 291
rect 526 288 534 291
rect 634 288 641 291
rect 666 288 667 292
rect 746 288 747 292
rect 893 288 894 292
rect 1021 288 1022 292
rect 1082 288 1089 291
rect 1362 288 1369 291
rect 1442 288 1443 292
rect 414 272 417 281
rect 702 278 713 281
rect 1222 278 1233 281
rect 294 268 302 271
rect 334 262 337 271
rect 358 268 369 271
rect 378 268 385 271
rect 596 268 598 272
rect 926 268 934 271
rect 974 271 978 272
rect 982 271 985 278
rect 1230 272 1233 278
rect 974 268 985 271
rect 154 258 162 261
rect 726 258 734 261
rect 766 258 777 261
rect 1334 258 1354 261
rect 1402 258 1409 261
rect 62 256 66 258
rect 158 256 162 258
rect 386 248 393 251
rect 398 248 401 258
rect 774 252 777 258
rect 1350 256 1354 258
rect 846 248 857 251
rect 878 248 889 251
rect 990 248 1006 251
rect 1102 248 1113 251
rect 1118 248 1129 251
rect 1322 248 1329 251
rect 1102 242 1105 248
rect 238 238 246 241
rect 318 238 326 241
rect 526 238 550 241
rect 1282 238 1289 241
rect 472 203 474 207
rect 478 203 481 207
rect 485 203 488 207
rect 381 188 382 192
rect 893 188 894 192
rect 1218 188 1219 192
rect 210 168 217 171
rect 294 168 305 171
rect 774 168 782 171
rect 802 168 809 171
rect 978 168 990 171
rect 1058 168 1073 171
rect 1418 168 1441 171
rect 294 162 297 168
rect 326 161 329 168
rect 310 158 321 161
rect 326 158 337 161
rect 398 161 401 168
rect 398 158 409 161
rect 654 158 665 161
rect 758 158 769 161
rect 1146 158 1153 161
rect 1230 158 1249 161
rect 1410 158 1417 161
rect 1422 158 1430 161
rect 386 148 401 151
rect 982 151 986 154
rect 982 148 998 151
rect 350 138 358 141
rect 398 138 401 148
rect 498 138 513 141
rect 598 138 606 141
rect 682 138 689 141
rect 902 138 913 141
rect 994 138 1009 141
rect 1198 138 1209 141
rect 686 128 689 138
rect 1322 128 1329 131
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 93 88 94 92
rect 122 88 123 92
rect 146 88 147 92
rect 210 88 211 92
rect 234 88 241 91
rect 421 88 422 92
rect 733 88 734 92
rect 757 88 758 92
rect 797 88 798 92
rect 1093 88 1094 92
rect 1117 88 1118 92
rect 1157 88 1158 92
rect 1202 88 1203 92
rect 1349 88 1350 92
rect 474 78 489 81
rect 998 81 1001 88
rect 986 78 1001 81
rect 1446 78 1462 81
rect 38 68 49 71
rect 190 68 198 71
rect 278 71 281 78
rect 278 68 289 71
rect 366 68 374 71
rect 430 68 446 71
rect 542 68 553 71
rect 686 68 697 71
rect 742 68 750 71
rect 830 68 838 71
rect 846 68 857 71
rect 878 68 886 71
rect 1078 68 1086 71
rect 1254 68 1265 71
rect 1278 68 1289 71
rect 1390 68 1401 71
rect 358 61 361 68
rect 1262 62 1265 68
rect 346 58 361 61
rect 522 58 529 61
rect 878 58 897 61
rect 1050 58 1057 61
rect 1182 58 1193 61
rect 1310 58 1329 61
rect 14 48 25 51
rect 78 48 89 51
rect 150 48 161 51
rect 302 48 313 51
rect 502 51 505 58
rect 406 48 417 51
rect 494 48 505 51
rect 566 48 585 51
rect 646 48 665 51
rect 718 48 729 51
rect 746 48 753 51
rect 782 48 793 51
rect 878 48 881 58
rect 1190 52 1193 58
rect 950 48 961 51
rect 990 48 1017 51
rect 1134 48 1153 51
rect 1310 48 1313 58
rect 1338 48 1345 51
rect 286 41 289 48
rect 374 42 378 44
rect 286 38 297 41
rect 506 38 513 41
rect 472 3 474 7
rect 478 3 481 7
rect 485 3 488 7
<< m2contact >>
rect 474 1403 478 1407
rect 481 1403 485 1407
rect 574 1378 578 1382
rect 630 1378 634 1382
rect 622 1368 626 1372
rect 678 1368 682 1372
rect 1382 1368 1386 1372
rect 1422 1368 1426 1372
rect 78 1358 82 1362
rect 150 1358 154 1362
rect 198 1358 202 1362
rect 294 1358 298 1362
rect 358 1358 362 1362
rect 398 1358 402 1362
rect 222 1348 226 1352
rect 246 1348 250 1352
rect 334 1348 338 1352
rect 358 1348 362 1352
rect 430 1348 434 1352
rect 454 1358 458 1362
rect 638 1358 642 1362
rect 646 1358 650 1362
rect 694 1358 698 1362
rect 526 1348 530 1352
rect 558 1348 562 1352
rect 606 1348 610 1352
rect 622 1348 626 1352
rect 686 1348 690 1352
rect 726 1358 730 1362
rect 774 1358 778 1362
rect 958 1358 962 1362
rect 982 1358 986 1362
rect 1022 1358 1026 1362
rect 1094 1358 1098 1362
rect 1126 1358 1130 1362
rect 1150 1358 1154 1362
rect 1174 1358 1178 1362
rect 1190 1358 1194 1362
rect 1214 1358 1218 1362
rect 1230 1358 1234 1362
rect 1246 1358 1250 1362
rect 1398 1358 1402 1362
rect 1406 1358 1410 1362
rect 1446 1358 1450 1362
rect 742 1348 746 1352
rect 870 1348 874 1352
rect 894 1348 898 1352
rect 1006 1348 1010 1352
rect 1022 1348 1026 1352
rect 1046 1348 1050 1352
rect 1102 1348 1106 1352
rect 1230 1348 1234 1352
rect 1414 1348 1418 1352
rect 6 1338 10 1342
rect 38 1338 42 1342
rect 54 1338 58 1342
rect 94 1338 98 1342
rect 150 1338 154 1342
rect 190 1338 194 1342
rect 238 1338 242 1342
rect 262 1338 266 1342
rect 270 1338 274 1342
rect 326 1338 330 1342
rect 374 1338 378 1342
rect 454 1338 458 1342
rect 494 1338 498 1342
rect 590 1338 594 1342
rect 646 1338 650 1342
rect 662 1338 666 1342
rect 702 1338 706 1342
rect 774 1338 778 1342
rect 798 1338 802 1342
rect 838 1338 842 1342
rect 934 1338 938 1342
rect 950 1338 954 1342
rect 998 1338 1002 1342
rect 1062 1338 1066 1342
rect 1142 1338 1146 1342
rect 1166 1338 1170 1342
rect 1238 1338 1242 1342
rect 1262 1338 1266 1342
rect 1302 1338 1306 1342
rect 1358 1338 1362 1342
rect 1382 1338 1386 1342
rect 134 1328 138 1332
rect 166 1328 170 1332
rect 238 1328 242 1332
rect 294 1328 298 1332
rect 318 1328 322 1332
rect 406 1328 410 1332
rect 526 1328 530 1332
rect 582 1328 586 1332
rect 766 1328 770 1332
rect 830 1328 834 1332
rect 870 1328 874 1332
rect 902 1328 906 1332
rect 950 1328 954 1332
rect 1054 1328 1058 1332
rect 1086 1328 1090 1332
rect 1118 1328 1122 1332
rect 1198 1328 1202 1332
rect 1206 1328 1210 1332
rect 1270 1328 1274 1332
rect 1310 1328 1314 1332
rect 1350 1328 1354 1332
rect 1446 1328 1450 1332
rect 22 1318 26 1322
rect 70 1318 74 1322
rect 86 1318 90 1322
rect 118 1318 122 1322
rect 174 1318 178 1322
rect 198 1318 202 1322
rect 278 1318 282 1322
rect 358 1318 362 1322
rect 398 1318 402 1322
rect 510 1318 514 1322
rect 678 1318 682 1322
rect 718 1318 722 1322
rect 814 1318 818 1322
rect 846 1318 850 1322
rect 926 1318 930 1322
rect 1030 1318 1034 1322
rect 1078 1318 1082 1322
rect 1134 1318 1138 1322
rect 1158 1318 1162 1322
rect 1254 1318 1258 1322
rect 1294 1318 1298 1322
rect 1334 1318 1338 1322
rect 1374 1318 1378 1322
rect 1414 1318 1418 1322
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 222 1288 226 1292
rect 686 1288 690 1292
rect 30 1278 34 1282
rect 182 1278 186 1282
rect 270 1278 274 1282
rect 334 1278 338 1282
rect 342 1278 346 1282
rect 350 1278 354 1282
rect 398 1278 402 1282
rect 462 1278 466 1282
rect 526 1278 530 1282
rect 542 1278 546 1282
rect 558 1278 562 1282
rect 566 1278 570 1282
rect 662 1278 666 1282
rect 670 1278 674 1282
rect 710 1278 714 1282
rect 758 1278 762 1282
rect 894 1278 898 1282
rect 902 1278 906 1282
rect 974 1278 978 1282
rect 998 1278 1002 1282
rect 30 1268 34 1272
rect 182 1268 186 1272
rect 262 1268 266 1272
rect 270 1268 274 1272
rect 302 1268 306 1272
rect 334 1268 338 1272
rect 454 1268 458 1272
rect 462 1268 466 1272
rect 574 1268 578 1272
rect 630 1268 634 1272
rect 718 1268 722 1272
rect 886 1268 890 1272
rect 966 1268 970 1272
rect 1030 1268 1034 1272
rect 1094 1278 1098 1282
rect 1118 1278 1122 1282
rect 1142 1278 1146 1282
rect 1190 1278 1194 1282
rect 1318 1278 1322 1282
rect 1358 1278 1362 1282
rect 1046 1268 1050 1272
rect 1070 1268 1074 1272
rect 1086 1268 1090 1272
rect 1102 1268 1106 1272
rect 1222 1268 1226 1272
rect 1310 1268 1314 1272
rect 1366 1268 1370 1272
rect 6 1258 10 1262
rect 54 1258 58 1262
rect 78 1258 82 1262
rect 102 1258 106 1262
rect 142 1258 146 1262
rect 158 1258 162 1262
rect 206 1258 210 1262
rect 238 1258 242 1262
rect 294 1258 298 1262
rect 302 1258 306 1262
rect 366 1258 370 1262
rect 374 1258 378 1262
rect 422 1258 426 1262
rect 438 1258 442 1262
rect 502 1258 506 1262
rect 590 1258 594 1262
rect 614 1258 618 1262
rect 734 1258 738 1262
rect 758 1258 762 1262
rect 790 1258 794 1262
rect 822 1258 826 1262
rect 854 1258 858 1262
rect 870 1258 874 1262
rect 934 1258 938 1262
rect 950 1258 954 1262
rect 1070 1258 1074 1262
rect 1142 1258 1146 1262
rect 1166 1258 1170 1262
rect 1190 1258 1194 1262
rect 1246 1258 1250 1262
rect 1278 1258 1282 1262
rect 1294 1258 1298 1262
rect 1342 1258 1346 1262
rect 1382 1258 1386 1262
rect 1398 1258 1402 1262
rect 1430 1258 1434 1262
rect 86 1248 90 1252
rect 94 1248 98 1252
rect 150 1248 154 1252
rect 214 1248 218 1252
rect 278 1248 282 1252
rect 358 1248 362 1252
rect 430 1248 434 1252
rect 486 1248 490 1252
rect 622 1248 626 1252
rect 766 1248 770 1252
rect 798 1248 802 1252
rect 830 1248 834 1252
rect 862 1248 866 1252
rect 902 1248 906 1252
rect 942 1248 946 1252
rect 1086 1248 1090 1252
rect 1150 1248 1154 1252
rect 1254 1248 1258 1252
rect 1286 1248 1290 1252
rect 1350 1248 1354 1252
rect 1390 1248 1394 1252
rect 1422 1248 1426 1252
rect 70 1238 74 1242
rect 110 1238 114 1242
rect 134 1238 138 1242
rect 198 1238 202 1242
rect 414 1238 418 1242
rect 542 1238 546 1242
rect 606 1238 610 1242
rect 630 1238 634 1242
rect 750 1238 754 1242
rect 782 1238 786 1242
rect 814 1238 818 1242
rect 822 1238 826 1242
rect 846 1238 850 1242
rect 926 1238 930 1242
rect 1134 1238 1138 1242
rect 1174 1238 1178 1242
rect 1222 1238 1226 1242
rect 1238 1238 1242 1242
rect 1270 1238 1274 1242
rect 1334 1238 1338 1242
rect 1406 1238 1410 1242
rect 1438 1238 1442 1242
rect 918 1228 922 1232
rect 78 1218 82 1222
rect 102 1218 106 1222
rect 126 1218 130 1222
rect 190 1218 194 1222
rect 246 1218 250 1222
rect 422 1218 426 1222
rect 534 1218 538 1222
rect 614 1218 618 1222
rect 790 1218 794 1222
rect 854 1218 858 1222
rect 1022 1218 1026 1222
rect 1246 1218 1250 1222
rect 1278 1218 1282 1222
rect 1342 1218 1346 1222
rect 1398 1218 1402 1222
rect 1430 1218 1434 1222
rect 474 1203 478 1207
rect 481 1203 485 1207
rect 14 1188 18 1192
rect 710 1188 714 1192
rect 1390 1188 1394 1192
rect 70 1178 74 1182
rect 678 1178 682 1182
rect 62 1168 66 1172
rect 102 1168 106 1172
rect 126 1168 130 1172
rect 654 1168 658 1172
rect 670 1168 674 1172
rect 702 1168 706 1172
rect 822 1168 826 1172
rect 1286 1178 1290 1182
rect 838 1168 842 1172
rect 854 1168 858 1172
rect 894 1168 898 1172
rect 942 1168 946 1172
rect 950 1168 954 1172
rect 1014 1168 1018 1172
rect 1126 1168 1130 1172
rect 1134 1168 1138 1172
rect 1246 1168 1250 1172
rect 1278 1168 1282 1172
rect 1310 1168 1314 1172
rect 1342 1168 1346 1172
rect 1398 1168 1402 1172
rect 46 1158 50 1162
rect 78 1158 82 1162
rect 110 1158 114 1162
rect 134 1158 138 1162
rect 206 1158 210 1162
rect 366 1158 370 1162
rect 430 1158 434 1162
rect 446 1158 450 1162
rect 542 1158 546 1162
rect 686 1158 690 1162
rect 838 1158 842 1162
rect 870 1158 874 1162
rect 966 1158 970 1162
rect 1078 1158 1082 1162
rect 1142 1158 1146 1162
rect 1190 1158 1194 1162
rect 1206 1158 1210 1162
rect 1262 1158 1266 1162
rect 1294 1158 1298 1162
rect 1326 1158 1330 1162
rect 1358 1158 1362 1162
rect 22 1148 26 1152
rect 70 1148 74 1152
rect 102 1148 106 1152
rect 134 1148 138 1152
rect 342 1148 346 1152
rect 454 1148 458 1152
rect 678 1148 682 1152
rect 710 1148 714 1152
rect 806 1148 810 1152
rect 822 1148 826 1152
rect 862 1148 866 1152
rect 886 1148 890 1152
rect 934 1148 938 1152
rect 958 1148 962 1152
rect 1110 1148 1114 1152
rect 1134 1148 1138 1152
rect 1206 1148 1210 1152
rect 1230 1148 1234 1152
rect 1254 1148 1258 1152
rect 1286 1148 1290 1152
rect 1318 1148 1322 1152
rect 1350 1148 1354 1152
rect 1390 1148 1394 1152
rect 1430 1148 1434 1152
rect 1454 1148 1458 1152
rect 150 1138 154 1142
rect 182 1138 186 1142
rect 190 1138 194 1142
rect 262 1138 266 1142
rect 318 1138 322 1142
rect 350 1138 354 1142
rect 382 1138 386 1142
rect 406 1138 410 1142
rect 430 1138 434 1142
rect 510 1138 514 1142
rect 582 1138 586 1142
rect 598 1138 602 1142
rect 654 1138 658 1142
rect 726 1138 730 1142
rect 774 1138 778 1142
rect 790 1138 794 1142
rect 918 1138 922 1142
rect 1022 1138 1026 1142
rect 1094 1138 1098 1142
rect 1182 1138 1186 1142
rect 1246 1138 1250 1142
rect 1366 1138 1370 1142
rect 158 1128 162 1132
rect 222 1128 226 1132
rect 254 1128 258 1132
rect 286 1128 290 1132
rect 374 1128 378 1132
rect 478 1128 482 1132
rect 518 1128 522 1132
rect 550 1128 554 1132
rect 590 1128 594 1132
rect 622 1128 626 1132
rect 742 1128 746 1132
rect 910 1128 914 1132
rect 982 1128 986 1132
rect 1062 1128 1066 1132
rect 1070 1128 1074 1132
rect 1086 1128 1090 1132
rect 1150 1128 1154 1132
rect 1374 1128 1378 1132
rect 46 1118 50 1122
rect 94 1118 98 1122
rect 134 1118 138 1122
rect 206 1118 210 1122
rect 238 1118 242 1122
rect 278 1118 282 1122
rect 310 1118 314 1122
rect 326 1118 330 1122
rect 366 1118 370 1122
rect 398 1118 402 1122
rect 422 1118 426 1122
rect 446 1118 450 1122
rect 494 1118 498 1122
rect 542 1118 546 1122
rect 574 1118 578 1122
rect 614 1118 618 1122
rect 734 1118 738 1122
rect 766 1118 770 1122
rect 846 1118 850 1122
rect 902 1118 906 1122
rect 1046 1118 1050 1122
rect 1174 1118 1178 1122
rect 1310 1118 1314 1122
rect 1342 1118 1346 1122
rect 1414 1118 1418 1122
rect 1438 1118 1442 1122
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 790 1088 794 1092
rect 1222 1088 1226 1092
rect 1462 1088 1466 1092
rect 230 1078 234 1082
rect 302 1078 306 1082
rect 334 1078 338 1082
rect 374 1078 378 1082
rect 550 1078 554 1082
rect 566 1078 570 1082
rect 630 1078 634 1082
rect 670 1078 674 1082
rect 678 1078 682 1082
rect 774 1078 778 1082
rect 854 1078 858 1082
rect 958 1078 962 1082
rect 966 1078 970 1082
rect 998 1078 1002 1082
rect 1086 1078 1090 1082
rect 1150 1078 1154 1082
rect 1198 1078 1202 1082
rect 1390 1078 1394 1082
rect 1398 1078 1402 1082
rect 1438 1078 1442 1082
rect 6 1068 10 1072
rect 166 1068 170 1072
rect 270 1068 274 1072
rect 326 1068 330 1072
rect 382 1068 386 1072
rect 518 1068 522 1072
rect 534 1068 538 1072
rect 550 1068 554 1072
rect 622 1068 626 1072
rect 686 1068 690 1072
rect 742 1068 746 1072
rect 782 1068 786 1072
rect 950 1068 954 1072
rect 1006 1068 1010 1072
rect 1094 1068 1098 1072
rect 1158 1068 1162 1072
rect 1214 1068 1218 1072
rect 1382 1068 1386 1072
rect 1430 1068 1434 1072
rect 1446 1068 1450 1072
rect 62 1058 66 1062
rect 86 1058 90 1062
rect 118 1058 122 1062
rect 142 1058 146 1062
rect 198 1058 202 1062
rect 230 1058 234 1062
rect 254 1058 258 1062
rect 358 1058 362 1062
rect 398 1058 402 1062
rect 422 1058 426 1062
rect 454 1058 458 1062
rect 494 1058 498 1062
rect 590 1058 594 1062
rect 606 1058 610 1062
rect 702 1058 706 1062
rect 718 1058 722 1062
rect 822 1058 826 1062
rect 854 1058 858 1062
rect 878 1058 882 1062
rect 918 1058 922 1062
rect 1022 1058 1026 1062
rect 1038 1058 1042 1062
rect 1078 1058 1082 1062
rect 1110 1058 1114 1062
rect 1134 1058 1138 1062
rect 1174 1058 1178 1062
rect 1198 1058 1202 1062
rect 1254 1058 1258 1062
rect 1286 1058 1290 1062
rect 1310 1058 1314 1062
rect 1342 1058 1346 1062
rect 1366 1058 1370 1062
rect 94 1048 98 1052
rect 126 1048 130 1052
rect 182 1048 186 1052
rect 190 1048 194 1052
rect 238 1048 242 1052
rect 302 1048 306 1052
rect 366 1048 370 1052
rect 430 1048 434 1052
rect 494 1048 498 1052
rect 518 1048 522 1052
rect 534 1048 538 1052
rect 598 1048 602 1052
rect 718 1048 722 1052
rect 742 1048 746 1052
rect 830 1048 834 1052
rect 862 1048 866 1052
rect 870 1048 874 1052
rect 926 1048 930 1052
rect 934 1048 938 1052
rect 982 1048 986 1052
rect 1030 1048 1034 1052
rect 1062 1048 1066 1052
rect 1142 1048 1146 1052
rect 1262 1048 1266 1052
rect 1294 1048 1298 1052
rect 1302 1048 1306 1052
rect 1334 1048 1338 1052
rect 78 1038 82 1042
rect 86 1038 90 1042
rect 110 1038 114 1042
rect 150 1038 154 1042
rect 206 1038 210 1042
rect 246 1038 250 1042
rect 254 1038 258 1042
rect 350 1038 354 1042
rect 414 1038 418 1042
rect 446 1038 450 1042
rect 502 1038 506 1042
rect 582 1038 586 1042
rect 726 1038 730 1042
rect 814 1038 818 1042
rect 846 1038 850 1042
rect 878 1038 882 1042
rect 886 1038 890 1042
rect 910 1038 914 1042
rect 1046 1038 1050 1042
rect 1126 1038 1130 1042
rect 1190 1038 1194 1042
rect 1262 1038 1266 1042
rect 1278 1038 1282 1042
rect 1318 1038 1322 1042
rect 1350 1038 1354 1042
rect 1430 1038 1434 1042
rect 278 1028 282 1032
rect 1134 1028 1138 1032
rect 1342 1028 1346 1032
rect 30 1018 34 1022
rect 46 1018 50 1022
rect 118 1018 122 1022
rect 158 1018 162 1022
rect 174 1018 178 1022
rect 198 1018 202 1022
rect 358 1018 362 1022
rect 422 1018 426 1022
rect 454 1018 458 1022
rect 510 1018 514 1022
rect 574 1018 578 1022
rect 646 1018 650 1022
rect 718 1018 722 1022
rect 806 1018 810 1022
rect 902 1018 906 1022
rect 1038 1018 1042 1022
rect 1254 1018 1258 1022
rect 1286 1018 1290 1022
rect 1310 1018 1314 1022
rect 474 1003 478 1007
rect 481 1003 485 1007
rect 222 988 226 992
rect 398 988 402 992
rect 950 988 954 992
rect 1062 988 1066 992
rect 22 978 26 982
rect 558 978 562 982
rect 14 968 18 972
rect 78 968 82 972
rect 94 968 98 972
rect 174 968 178 972
rect 198 968 202 972
rect 230 968 234 972
rect 334 968 338 972
rect 422 968 426 972
rect 454 968 458 972
rect 502 968 506 972
rect 534 968 538 972
rect 622 968 626 972
rect 654 968 658 972
rect 678 968 682 972
rect 830 968 834 972
rect 870 968 874 972
rect 958 968 962 972
rect 1070 968 1074 972
rect 1094 968 1098 972
rect 1190 968 1194 972
rect 1198 968 1202 972
rect 1302 968 1306 972
rect 1342 968 1346 972
rect 1358 968 1362 972
rect 1438 978 1442 982
rect 1374 968 1378 972
rect 1390 968 1394 972
rect 1446 968 1450 972
rect 30 958 34 962
rect 174 958 178 962
rect 182 958 186 962
rect 214 958 218 962
rect 310 958 314 962
rect 318 958 322 962
rect 390 958 394 962
rect 438 958 442 962
rect 470 958 474 962
rect 518 958 522 962
rect 550 958 554 962
rect 606 958 610 962
rect 638 958 642 962
rect 694 958 698 962
rect 846 958 850 962
rect 854 958 858 962
rect 910 958 914 962
rect 974 958 978 962
rect 1030 958 1034 962
rect 1054 958 1058 962
rect 1102 958 1106 962
rect 1182 958 1186 962
rect 1246 958 1250 962
rect 1318 958 1322 962
rect 1326 958 1330 962
rect 1358 958 1362 962
rect 1430 958 1434 962
rect 22 948 26 952
rect 38 948 42 952
rect 86 948 90 952
rect 142 948 146 952
rect 166 948 170 952
rect 190 948 194 952
rect 222 948 226 952
rect 246 948 250 952
rect 270 948 274 952
rect 334 948 338 952
rect 430 948 434 952
rect 462 948 466 952
rect 510 948 514 952
rect 542 948 546 952
rect 598 948 602 952
rect 614 948 618 952
rect 630 948 634 952
rect 646 948 650 952
rect 686 948 690 952
rect 742 948 746 952
rect 790 948 794 952
rect 838 948 842 952
rect 862 948 866 952
rect 886 948 890 952
rect 966 948 970 952
rect 990 948 994 952
rect 1062 948 1066 952
rect 1110 948 1114 952
rect 1134 948 1138 952
rect 1150 948 1154 952
rect 1190 948 1194 952
rect 1214 948 1218 952
rect 1262 948 1266 952
rect 1310 948 1314 952
rect 1334 948 1338 952
rect 1366 948 1370 952
rect 1438 948 1442 952
rect 54 938 58 942
rect 110 938 114 942
rect 118 938 122 942
rect 166 938 170 942
rect 262 938 266 942
rect 294 938 298 942
rect 334 938 338 942
rect 358 938 362 942
rect 582 938 586 942
rect 702 938 706 942
rect 758 938 762 942
rect 766 938 770 942
rect 870 938 874 942
rect 910 938 914 942
rect 1014 938 1018 942
rect 1030 938 1034 942
rect 1046 938 1050 942
rect 1086 938 1090 942
rect 1126 938 1130 942
rect 1134 938 1138 942
rect 1230 938 1234 942
rect 1254 938 1258 942
rect 1390 938 1394 942
rect 62 928 66 932
rect 118 928 122 932
rect 366 928 370 932
rect 406 928 410 932
rect 566 928 570 932
rect 574 928 578 932
rect 734 928 738 932
rect 942 928 946 932
rect 1022 928 1026 932
rect 1174 928 1178 932
rect 1238 928 1242 932
rect 1286 928 1290 932
rect 1422 928 1426 932
rect 78 918 82 922
rect 190 918 194 922
rect 286 918 290 922
rect 302 918 306 922
rect 382 918 386 922
rect 430 918 434 922
rect 462 918 466 922
rect 494 918 498 922
rect 534 918 538 922
rect 646 918 650 922
rect 670 918 674 922
rect 710 918 714 922
rect 814 918 818 922
rect 822 918 826 922
rect 1310 918 1314 922
rect 1334 918 1338 922
rect 986 903 990 907
rect 993 903 997 907
rect 30 888 34 892
rect 254 888 258 892
rect 518 888 522 892
rect 654 888 658 892
rect 734 888 738 892
rect 1182 888 1186 892
rect 1206 888 1210 892
rect 1246 888 1250 892
rect 1270 888 1274 892
rect 1382 888 1386 892
rect 358 878 362 882
rect 390 878 394 882
rect 558 878 562 882
rect 630 878 634 882
rect 774 878 778 882
rect 838 878 842 882
rect 878 878 882 882
rect 934 878 938 882
rect 1006 878 1010 882
rect 1054 878 1058 882
rect 1078 878 1082 882
rect 1150 878 1154 882
rect 1158 878 1162 882
rect 1166 878 1170 882
rect 1230 878 1234 882
rect 1302 878 1306 882
rect 1438 878 1442 882
rect 6 868 10 872
rect 54 868 58 872
rect 70 868 74 872
rect 190 868 194 872
rect 246 868 250 872
rect 350 868 354 872
rect 390 868 394 872
rect 510 868 514 872
rect 526 868 530 872
rect 614 868 618 872
rect 638 868 642 872
rect 726 868 730 872
rect 742 868 746 872
rect 766 868 770 872
rect 830 868 834 872
rect 894 868 898 872
rect 902 868 906 872
rect 966 868 970 872
rect 22 858 26 862
rect 46 858 50 862
rect 86 858 90 862
rect 102 858 106 862
rect 134 858 138 862
rect 166 858 170 862
rect 222 858 226 862
rect 278 858 282 862
rect 310 858 314 862
rect 334 858 338 862
rect 366 858 370 862
rect 406 858 410 862
rect 446 858 450 862
rect 494 858 498 862
rect 582 858 586 862
rect 598 858 602 862
rect 670 858 674 862
rect 702 858 706 862
rect 798 858 802 862
rect 814 858 818 862
rect 894 858 898 862
rect 934 858 938 862
rect 958 858 962 862
rect 1038 868 1042 872
rect 1030 858 1034 862
rect 1086 868 1090 872
rect 1102 868 1106 872
rect 1190 868 1194 872
rect 1238 868 1242 872
rect 1262 868 1266 872
rect 1286 868 1290 872
rect 1350 868 1354 872
rect 1374 868 1378 872
rect 1446 868 1450 872
rect 1062 858 1066 862
rect 1126 858 1130 862
rect 1326 858 1330 862
rect 1414 858 1418 862
rect 126 848 130 852
rect 158 848 162 852
rect 206 848 210 852
rect 214 848 218 852
rect 262 848 266 852
rect 270 848 274 852
rect 302 848 306 852
rect 398 848 402 852
rect 454 848 458 852
rect 502 848 506 852
rect 590 848 594 852
rect 662 848 666 852
rect 694 848 698 852
rect 742 848 746 852
rect 782 848 786 852
rect 902 848 906 852
rect 942 848 946 852
rect 998 848 1002 852
rect 1014 848 1018 852
rect 1102 848 1106 852
rect 1174 848 1178 852
rect 1254 848 1258 852
rect 1278 848 1282 852
rect 1366 848 1370 852
rect 1398 848 1402 852
rect 1438 848 1442 852
rect 1462 848 1466 852
rect 102 838 106 842
rect 110 838 114 842
rect 142 838 146 842
rect 174 838 178 842
rect 230 838 234 842
rect 278 838 282 842
rect 286 838 290 842
rect 318 838 322 842
rect 414 838 418 842
rect 438 838 442 842
rect 486 838 490 842
rect 574 838 578 842
rect 678 838 682 842
rect 710 838 714 842
rect 798 838 802 842
rect 974 838 978 842
rect 1062 838 1066 842
rect 166 828 170 832
rect 198 828 202 832
rect 310 828 314 832
rect 534 828 538 832
rect 854 828 858 832
rect 1326 828 1330 832
rect 62 818 66 822
rect 118 818 122 822
rect 134 818 138 822
rect 222 818 226 822
rect 406 818 410 822
rect 430 818 434 822
rect 494 818 498 822
rect 582 818 586 822
rect 670 818 674 822
rect 718 818 722 822
rect 790 818 794 822
rect 1294 818 1298 822
rect 474 803 478 807
rect 481 803 485 807
rect 174 788 178 792
rect 270 788 274 792
rect 294 788 298 792
rect 606 788 610 792
rect 726 788 730 792
rect 1254 788 1258 792
rect 1470 788 1474 792
rect 6 778 10 782
rect 694 778 698 782
rect 1438 778 1442 782
rect 502 768 506 772
rect 638 768 642 772
rect 670 768 674 772
rect 702 768 706 772
rect 734 768 738 772
rect 1006 768 1010 772
rect 1118 768 1122 772
rect 622 758 626 762
rect 654 758 658 762
rect 686 758 690 762
rect 718 758 722 762
rect 750 758 754 762
rect 766 758 770 762
rect 1030 758 1034 762
rect 1062 758 1066 762
rect 1094 758 1098 762
rect 94 747 98 751
rect 126 748 130 752
rect 206 748 210 752
rect 230 748 234 752
rect 286 748 290 752
rect 326 748 330 752
rect 350 748 354 752
rect 406 748 410 752
rect 478 748 482 752
rect 566 747 570 751
rect 598 748 602 752
rect 630 748 634 752
rect 662 748 666 752
rect 694 748 698 752
rect 726 748 730 752
rect 814 748 818 752
rect 846 748 850 752
rect 878 748 882 752
rect 910 748 914 752
rect 134 738 138 742
rect 150 738 154 742
rect 166 738 170 742
rect 374 738 378 742
rect 390 738 394 742
rect 414 738 418 742
rect 430 738 434 742
rect 494 738 498 742
rect 558 738 562 742
rect 942 747 946 751
rect 1022 748 1026 752
rect 1046 748 1050 752
rect 1174 748 1178 752
rect 1286 748 1290 752
rect 1302 748 1306 752
rect 1318 748 1322 752
rect 1350 747 1354 751
rect 750 738 754 742
rect 766 738 770 742
rect 790 738 794 742
rect 806 738 810 742
rect 838 738 842 742
rect 870 738 874 742
rect 902 738 906 742
rect 926 738 930 742
rect 1054 738 1058 742
rect 1078 738 1082 742
rect 1094 738 1098 742
rect 1126 738 1130 742
rect 1262 738 1266 742
rect 1278 738 1282 742
rect 1310 738 1314 742
rect 1454 738 1458 742
rect 94 728 98 732
rect 150 728 154 732
rect 430 728 434 732
rect 446 728 450 732
rect 822 728 826 732
rect 854 728 858 732
rect 886 728 890 732
rect 1062 728 1066 732
rect 1094 728 1098 732
rect 1134 728 1138 732
rect 1166 728 1170 732
rect 1262 728 1266 732
rect 1294 728 1298 732
rect 1350 728 1354 732
rect 1446 728 1450 732
rect 398 718 402 722
rect 422 718 426 722
rect 462 718 466 722
rect 630 718 634 722
rect 662 718 666 722
rect 798 718 802 722
rect 830 718 834 722
rect 862 718 866 722
rect 894 718 898 722
rect 986 703 990 707
rect 993 703 997 707
rect 142 688 146 692
rect 174 688 178 692
rect 222 688 226 692
rect 470 688 474 692
rect 870 688 874 692
rect 910 688 914 692
rect 942 688 946 692
rect 1222 688 1226 692
rect 94 678 98 682
rect 150 678 154 682
rect 182 678 186 682
rect 214 678 218 682
rect 598 678 602 682
rect 614 678 618 682
rect 638 678 642 682
rect 654 678 658 682
rect 718 678 722 682
rect 782 678 786 682
rect 846 678 850 682
rect 1246 678 1250 682
rect 1286 678 1290 682
rect 1350 678 1354 682
rect 6 668 10 672
rect 134 668 138 672
rect 166 668 170 672
rect 198 668 202 672
rect 214 668 218 672
rect 270 668 274 672
rect 558 668 562 672
rect 582 668 586 672
rect 598 668 602 672
rect 622 668 626 672
rect 686 668 690 672
rect 726 668 730 672
rect 790 668 794 672
rect 1022 668 1026 672
rect 1118 668 1122 672
rect 1166 668 1170 672
rect 1270 668 1274 672
rect 1294 668 1298 672
rect 1310 668 1314 672
rect 1470 668 1474 672
rect 86 658 90 662
rect 126 658 130 662
rect 158 658 162 662
rect 190 658 194 662
rect 262 658 266 662
rect 374 658 378 662
rect 390 658 394 662
rect 470 658 474 662
rect 510 658 514 662
rect 542 659 546 663
rect 574 658 578 662
rect 630 658 634 662
rect 654 658 658 662
rect 766 658 770 662
rect 806 658 810 662
rect 830 658 834 662
rect 862 658 866 662
rect 886 658 890 662
rect 910 658 914 662
rect 942 658 946 662
rect 974 658 978 662
rect 1038 659 1042 663
rect 1134 659 1138 663
rect 1198 658 1202 662
rect 1206 658 1210 662
rect 1246 658 1250 662
rect 1262 658 1266 662
rect 1318 658 1322 662
rect 1350 659 1354 663
rect 1422 658 1426 662
rect 1446 658 1450 662
rect 694 648 698 652
rect 742 648 746 652
rect 774 648 778 652
rect 830 648 834 652
rect 902 648 906 652
rect 934 648 938 652
rect 966 648 970 652
rect 1102 648 1106 652
rect 1254 648 1258 652
rect 318 638 322 642
rect 686 638 690 642
rect 758 638 762 642
rect 822 638 826 642
rect 878 638 882 642
rect 886 638 890 642
rect 950 638 954 642
rect 974 638 978 642
rect 982 638 986 642
rect 1246 638 1250 642
rect 1398 638 1402 642
rect 1414 638 1418 642
rect 1438 638 1442 642
rect 438 628 442 632
rect 702 628 706 632
rect 766 618 770 622
rect 830 618 834 622
rect 846 618 850 622
rect 1286 618 1290 622
rect 474 603 478 607
rect 481 603 485 607
rect 126 588 130 592
rect 406 588 410 592
rect 838 588 842 592
rect 878 588 882 592
rect 910 588 914 592
rect 1022 588 1026 592
rect 1246 588 1250 592
rect 1286 588 1290 592
rect 342 578 346 582
rect 374 578 378 582
rect 742 578 746 582
rect 1054 578 1058 582
rect 6 568 10 572
rect 118 568 122 572
rect 334 568 338 572
rect 366 568 370 572
rect 398 568 402 572
rect 502 568 506 572
rect 510 568 514 572
rect 558 568 562 572
rect 646 568 650 572
rect 734 568 738 572
rect 798 568 802 572
rect 806 568 810 572
rect 830 568 834 572
rect 870 568 874 572
rect 918 568 922 572
rect 942 568 946 572
rect 950 568 954 572
rect 1030 568 1034 572
rect 1062 568 1066 572
rect 1198 568 1202 572
rect 1214 568 1218 572
rect 1222 568 1226 572
rect 1254 568 1258 572
rect 1278 568 1282 572
rect 102 558 106 562
rect 286 558 290 562
rect 350 558 354 562
rect 382 558 386 562
rect 406 558 410 562
rect 422 558 426 562
rect 494 558 498 562
rect 614 558 618 562
rect 622 558 626 562
rect 662 558 666 562
rect 750 558 754 562
rect 814 558 818 562
rect 854 558 858 562
rect 934 558 938 562
rect 1014 558 1018 562
rect 1046 558 1050 562
rect 1238 558 1242 562
rect 1294 558 1298 562
rect 110 548 114 552
rect 318 548 322 552
rect 334 548 338 552
rect 374 548 378 552
rect 406 548 410 552
rect 422 548 426 552
rect 502 548 506 552
rect 582 548 586 552
rect 718 548 722 552
rect 742 548 746 552
rect 806 548 810 552
rect 838 548 842 552
rect 862 548 866 552
rect 902 548 906 552
rect 910 548 914 552
rect 942 548 946 552
rect 1022 548 1026 552
rect 1054 548 1058 552
rect 1078 548 1082 552
rect 1134 547 1138 551
rect 1166 548 1170 552
rect 1222 548 1226 552
rect 1246 548 1250 552
rect 1286 548 1290 552
rect 1366 547 1370 551
rect 1398 548 1402 552
rect 1438 548 1442 552
rect 38 538 42 542
rect 62 538 66 542
rect 94 538 98 542
rect 174 538 178 542
rect 206 538 210 542
rect 246 538 250 542
rect 302 538 306 542
rect 454 538 458 542
rect 558 538 562 542
rect 614 538 618 542
rect 638 538 642 542
rect 646 538 650 542
rect 686 538 690 542
rect 702 538 706 542
rect 766 538 770 542
rect 782 538 786 542
rect 886 538 890 542
rect 966 538 970 542
rect 982 538 986 542
rect 1094 538 1098 542
rect 1302 538 1306 542
rect 1478 538 1482 542
rect 30 528 34 532
rect 134 528 138 532
rect 254 528 258 532
rect 294 528 298 532
rect 446 528 450 532
rect 526 528 530 532
rect 566 528 570 532
rect 582 528 586 532
rect 758 528 762 532
rect 1006 528 1010 532
rect 1102 528 1106 532
rect 1334 528 1338 532
rect 14 518 18 522
rect 54 518 58 522
rect 78 518 82 522
rect 150 518 154 522
rect 182 518 186 522
rect 238 518 242 522
rect 430 518 434 522
rect 510 518 514 522
rect 662 518 666 522
rect 678 518 682 522
rect 1318 518 1322 522
rect 1430 518 1434 522
rect 986 503 990 507
rect 993 503 997 507
rect 126 488 130 492
rect 454 488 458 492
rect 590 488 594 492
rect 910 488 914 492
rect 942 488 946 492
rect 958 488 962 492
rect 1158 488 1162 492
rect 1190 488 1194 492
rect 1238 488 1242 492
rect 1270 488 1274 492
rect 6 478 10 482
rect 198 478 202 482
rect 286 478 290 482
rect 350 478 354 482
rect 382 478 386 482
rect 534 478 538 482
rect 550 478 554 482
rect 638 478 642 482
rect 734 478 738 482
rect 742 478 746 482
rect 790 478 794 482
rect 838 478 842 482
rect 886 478 890 482
rect 990 478 994 482
rect 1038 478 1042 482
rect 1046 478 1050 482
rect 1142 478 1146 482
rect 1174 478 1178 482
rect 1286 478 1290 482
rect 1302 478 1306 482
rect 1326 478 1330 482
rect 1470 478 1474 482
rect 46 468 50 472
rect 86 468 90 472
rect 102 468 106 472
rect 198 468 202 472
rect 278 468 282 472
rect 326 468 330 472
rect 342 468 346 472
rect 350 468 354 472
rect 390 468 394 472
rect 550 468 554 472
rect 606 468 610 472
rect 646 468 650 472
rect 702 468 706 472
rect 742 468 746 472
rect 782 468 786 472
rect 838 468 842 472
rect 846 468 850 472
rect 934 468 938 472
rect 974 468 978 472
rect 1078 468 1082 472
rect 1086 468 1090 472
rect 1134 468 1138 472
rect 1150 468 1154 472
rect 1206 468 1210 472
rect 1230 468 1234 472
rect 1262 468 1266 472
rect 1310 468 1314 472
rect 1382 468 1386 472
rect 1390 468 1394 472
rect 1462 468 1466 472
rect 30 458 34 462
rect 62 458 66 462
rect 118 458 122 462
rect 158 458 162 462
rect 174 458 178 462
rect 222 458 226 462
rect 238 458 242 462
rect 262 458 266 462
rect 302 458 306 462
rect 406 458 410 462
rect 422 458 426 462
rect 462 458 466 462
rect 510 458 514 462
rect 534 458 538 462
rect 566 458 570 462
rect 662 458 666 462
rect 678 458 682 462
rect 790 458 794 462
rect 806 458 810 462
rect 862 458 866 462
rect 878 458 882 462
rect 894 458 898 462
rect 910 458 914 462
rect 1014 458 1018 462
rect 1102 458 1106 462
rect 1342 458 1346 462
rect 1422 458 1426 462
rect 1446 458 1450 462
rect 46 448 50 452
rect 54 448 58 452
rect 86 448 90 452
rect 110 448 114 452
rect 166 448 170 452
rect 230 448 234 452
rect 294 448 298 452
rect 358 448 362 452
rect 374 448 378 452
rect 438 448 442 452
rect 470 448 474 452
rect 518 448 522 452
rect 534 448 538 452
rect 582 448 586 452
rect 622 448 626 452
rect 670 448 674 452
rect 702 448 706 452
rect 758 448 762 452
rect 774 448 778 452
rect 830 448 834 452
rect 70 438 74 442
rect 150 438 154 442
rect 246 438 250 442
rect 310 438 314 442
rect 422 438 426 442
rect 454 438 458 442
rect 502 438 506 442
rect 686 438 690 442
rect 878 438 882 442
rect 902 448 906 452
rect 950 448 954 452
rect 958 448 962 452
rect 1078 448 1082 452
rect 1110 448 1114 452
rect 1166 448 1170 452
rect 1214 448 1218 452
rect 1230 448 1234 452
rect 1238 448 1242 452
rect 1278 448 1282 452
rect 1286 448 1290 452
rect 1334 448 1338 452
rect 1366 448 1370 452
rect 910 438 914 442
rect 918 438 922 442
rect 1094 438 1098 442
rect 1102 438 1106 442
rect 1350 438 1354 442
rect 1430 438 1434 442
rect 430 428 434 432
rect 1374 428 1378 432
rect 142 418 146 422
rect 238 418 242 422
rect 302 418 306 422
rect 510 418 514 422
rect 678 418 682 422
rect 1342 418 1346 422
rect 1398 418 1402 422
rect 1422 418 1426 422
rect 474 403 478 407
rect 481 403 485 407
rect 22 388 26 392
rect 86 388 90 392
rect 126 388 130 392
rect 174 388 178 392
rect 382 388 386 392
rect 502 388 506 392
rect 534 388 538 392
rect 558 388 562 392
rect 574 388 578 392
rect 606 388 610 392
rect 670 388 674 392
rect 694 388 698 392
rect 742 388 746 392
rect 782 388 786 392
rect 870 388 874 392
rect 934 388 938 392
rect 1038 388 1042 392
rect 1070 388 1074 392
rect 1214 388 1218 392
rect 1278 388 1282 392
rect 1302 388 1306 392
rect 1334 388 1338 392
rect 1430 388 1434 392
rect 54 378 58 382
rect 1366 378 1370 382
rect 14 368 18 372
rect 46 368 50 372
rect 78 368 82 372
rect 118 368 122 372
rect 150 368 154 372
rect 166 368 170 372
rect 182 368 186 372
rect 374 368 378 372
rect 526 368 530 372
rect 582 368 586 372
rect 614 368 618 372
rect 638 368 642 372
rect 646 368 650 372
rect 678 368 682 372
rect 862 368 866 372
rect 894 368 898 372
rect 918 368 922 372
rect 942 368 946 372
rect 1078 368 1082 372
rect 1190 368 1194 372
rect 1238 368 1242 372
rect 1270 368 1274 372
rect 1310 368 1314 372
rect 1342 368 1346 372
rect 1374 368 1378 372
rect 1438 368 1442 372
rect 62 358 66 362
rect 94 358 98 362
rect 134 358 138 362
rect 166 358 170 362
rect 246 358 250 362
rect 286 358 290 362
rect 358 358 362 362
rect 390 358 394 362
rect 478 358 482 362
rect 22 348 26 352
rect 30 348 34 352
rect 54 348 58 352
rect 86 348 90 352
rect 110 348 114 352
rect 142 348 146 352
rect 174 348 178 352
rect 198 348 202 352
rect 222 348 226 352
rect 238 348 242 352
rect 382 348 386 352
rect 398 348 402 352
rect 446 348 450 352
rect 542 358 546 362
rect 566 358 570 362
rect 598 358 602 362
rect 630 358 634 362
rect 662 358 666 362
rect 798 358 802 362
rect 878 358 882 362
rect 910 358 914 362
rect 958 358 962 362
rect 966 358 970 362
rect 1030 358 1034 362
rect 1062 358 1066 362
rect 1206 358 1210 362
rect 1222 358 1226 362
rect 1254 358 1258 362
rect 1286 358 1290 362
rect 1294 358 1298 362
rect 1326 358 1330 362
rect 1358 358 1362 362
rect 1422 358 1426 362
rect 1454 358 1458 362
rect 534 348 538 352
rect 574 348 578 352
rect 606 348 610 352
rect 638 348 642 352
rect 670 348 674 352
rect 710 348 714 352
rect 782 348 786 352
rect 846 348 850 352
rect 870 348 874 352
rect 894 348 898 352
rect 950 348 954 352
rect 1014 348 1018 352
rect 1030 348 1034 352
rect 1054 348 1058 352
rect 1078 348 1082 352
rect 1110 348 1114 352
rect 1142 348 1146 352
rect 1174 348 1178 352
rect 1198 348 1202 352
rect 1246 348 1250 352
rect 1278 348 1282 352
rect 1302 348 1306 352
rect 1334 348 1338 352
rect 1366 348 1370 352
rect 1390 348 1394 352
rect 1430 348 1434 352
rect 214 338 218 342
rect 254 338 258 342
rect 326 338 330 342
rect 358 338 362 342
rect 414 338 418 342
rect 510 338 514 342
rect 550 338 554 342
rect 750 338 754 342
rect 822 338 826 342
rect 830 338 834 342
rect 1006 338 1010 342
rect 1126 338 1130 342
rect 1158 338 1162 342
rect 1406 338 1410 342
rect 1454 338 1458 342
rect 1470 338 1474 342
rect 286 328 290 332
rect 318 328 322 332
rect 326 328 330 332
rect 422 328 426 332
rect 430 328 434 332
rect 718 328 722 332
rect 758 328 762 332
rect 806 328 810 332
rect 822 328 826 332
rect 902 328 906 332
rect 918 328 922 332
rect 1094 328 1098 332
rect 1118 328 1122 332
rect 1150 328 1154 332
rect 1198 328 1202 332
rect 1222 328 1226 332
rect 1414 328 1418 332
rect 558 318 562 322
rect 974 318 978 322
rect 986 303 990 307
rect 993 303 997 307
rect 22 288 26 292
rect 70 288 74 292
rect 118 288 122 292
rect 150 288 154 292
rect 166 288 170 292
rect 206 288 210 292
rect 406 288 410 292
rect 422 288 426 292
rect 462 288 466 292
rect 478 288 482 292
rect 534 288 538 292
rect 630 288 634 292
rect 662 288 666 292
rect 742 288 746 292
rect 790 288 794 292
rect 822 288 826 292
rect 846 288 850 292
rect 894 288 898 292
rect 1022 288 1026 292
rect 1078 288 1082 292
rect 1190 288 1194 292
rect 1246 288 1250 292
rect 1310 288 1314 292
rect 1334 288 1338 292
rect 1358 288 1362 292
rect 1382 288 1386 292
rect 1422 288 1426 292
rect 1438 288 1442 292
rect 302 278 306 282
rect 374 278 378 282
rect 550 278 554 282
rect 558 278 562 282
rect 678 278 682 282
rect 758 278 762 282
rect 798 278 802 282
rect 862 278 866 282
rect 870 278 874 282
rect 934 278 938 282
rect 982 278 986 282
rect 1038 278 1042 282
rect 1134 278 1138 282
rect 1142 278 1146 282
rect 1174 278 1178 282
rect 38 268 42 272
rect 94 268 98 272
rect 110 268 114 272
rect 134 268 138 272
rect 302 268 306 272
rect 326 268 330 272
rect 374 268 378 272
rect 414 268 418 272
rect 510 268 514 272
rect 566 268 570 272
rect 598 268 602 272
rect 654 268 658 272
rect 694 268 698 272
rect 734 268 738 272
rect 774 268 778 272
rect 806 268 810 272
rect 830 268 834 272
rect 902 268 906 272
rect 934 268 938 272
rect 942 268 946 272
rect 1030 268 1034 272
rect 1046 268 1050 272
rect 1102 268 1106 272
rect 1150 268 1154 272
rect 1206 268 1210 272
rect 1230 268 1234 272
rect 1262 268 1266 272
rect 1342 268 1346 272
rect 1430 268 1434 272
rect 22 258 26 262
rect 62 258 66 262
rect 70 258 74 262
rect 102 258 106 262
rect 150 258 154 262
rect 166 258 170 262
rect 198 258 202 262
rect 222 258 226 262
rect 254 258 258 262
rect 278 258 282 262
rect 334 258 338 262
rect 350 258 354 262
rect 398 258 402 262
rect 438 258 442 262
rect 462 258 466 262
rect 534 258 538 262
rect 606 258 610 262
rect 630 258 634 262
rect 734 258 738 262
rect 910 258 914 262
rect 958 258 962 262
rect 982 258 986 262
rect 1078 258 1082 262
rect 1230 258 1234 262
rect 1278 258 1282 262
rect 1294 258 1298 262
rect 1310 258 1314 262
rect 1358 258 1362 262
rect 1398 258 1402 262
rect 30 248 34 252
rect 126 248 130 252
rect 150 248 154 252
rect 190 248 194 252
rect 246 248 250 252
rect 310 248 314 252
rect 334 248 338 252
rect 382 248 386 252
rect 470 248 474 252
rect 494 248 498 252
rect 542 248 546 252
rect 582 248 586 252
rect 614 248 618 252
rect 622 248 626 252
rect 670 248 674 252
rect 750 248 754 252
rect 774 248 778 252
rect 790 248 794 252
rect 1006 248 1010 252
rect 1014 248 1018 252
rect 1062 248 1066 252
rect 1070 248 1074 252
rect 1166 248 1170 252
rect 1190 248 1194 252
rect 1238 248 1242 252
rect 1246 248 1250 252
rect 1270 248 1274 252
rect 1318 248 1322 252
rect 1446 248 1450 252
rect 14 238 18 242
rect 78 238 82 242
rect 174 238 178 242
rect 206 238 210 242
rect 246 238 250 242
rect 262 238 266 242
rect 326 238 330 242
rect 454 238 458 242
rect 550 238 554 242
rect 574 238 578 242
rect 598 238 602 242
rect 638 238 642 242
rect 974 238 978 242
rect 1086 238 1090 242
rect 1102 238 1106 242
rect 1222 238 1226 242
rect 1278 238 1282 242
rect 1310 238 1314 242
rect 1366 238 1370 242
rect 254 228 258 232
rect 1182 228 1186 232
rect 46 218 50 222
rect 710 218 714 222
rect 1422 218 1426 222
rect 474 203 478 207
rect 481 203 485 207
rect 14 188 18 192
rect 78 188 82 192
rect 134 188 138 192
rect 206 188 210 192
rect 270 188 274 192
rect 382 188 386 192
rect 438 188 442 192
rect 462 188 466 192
rect 534 188 538 192
rect 558 188 562 192
rect 622 188 626 192
rect 726 188 730 192
rect 798 188 802 192
rect 894 188 898 192
rect 942 188 946 192
rect 958 188 962 192
rect 1126 188 1130 192
rect 1214 188 1218 192
rect 1278 188 1282 192
rect 1366 188 1370 192
rect 1430 188 1434 192
rect 22 168 26 172
rect 86 168 90 172
rect 142 168 146 172
rect 206 168 210 172
rect 278 168 282 172
rect 326 168 330 172
rect 398 168 402 172
rect 430 168 434 172
rect 470 168 474 172
rect 566 168 570 172
rect 630 168 634 172
rect 734 168 738 172
rect 782 168 786 172
rect 798 168 802 172
rect 934 168 938 172
rect 966 168 970 172
rect 974 168 978 172
rect 990 168 994 172
rect 1038 168 1042 172
rect 1046 168 1050 172
rect 1054 168 1058 172
rect 1110 168 1114 172
rect 1134 168 1138 172
rect 1270 168 1274 172
rect 1374 168 1378 172
rect 1398 168 1402 172
rect 1414 168 1418 172
rect 6 158 10 162
rect 70 158 74 162
rect 158 158 162 162
rect 198 158 202 162
rect 262 158 266 162
rect 294 158 298 162
rect 366 158 370 162
rect 414 158 418 162
rect 446 158 450 162
rect 454 158 458 162
rect 550 158 554 162
rect 614 158 618 162
rect 718 158 722 162
rect 790 158 794 162
rect 878 158 882 162
rect 950 158 954 162
rect 982 158 986 162
rect 1062 158 1066 162
rect 1142 158 1146 162
rect 1254 158 1258 162
rect 1286 158 1290 162
rect 1294 158 1298 162
rect 1358 158 1362 162
rect 1406 158 1410 162
rect 1430 158 1434 162
rect 14 148 18 152
rect 86 148 90 152
rect 102 148 106 152
rect 150 148 154 152
rect 166 148 170 152
rect 214 148 218 152
rect 230 148 234 152
rect 270 148 274 152
rect 382 148 386 152
rect 438 148 442 152
rect 462 148 466 152
rect 558 148 562 152
rect 622 148 626 152
rect 710 148 714 152
rect 726 148 730 152
rect 806 148 810 152
rect 822 148 826 152
rect 846 148 850 152
rect 894 148 898 152
rect 942 148 946 152
rect 974 148 978 152
rect 998 148 1002 152
rect 1054 148 1058 152
rect 1142 148 1146 152
rect 1158 148 1162 152
rect 1214 148 1218 152
rect 1278 148 1282 152
rect 1350 148 1354 152
rect 1366 148 1370 152
rect 1406 148 1410 152
rect 1430 148 1434 152
rect 38 138 42 142
rect 54 138 58 142
rect 118 138 122 142
rect 182 138 186 142
rect 246 138 250 142
rect 294 138 298 142
rect 358 138 362 142
rect 390 138 394 142
rect 494 138 498 142
rect 606 138 610 142
rect 678 138 682 142
rect 694 138 698 142
rect 782 138 786 142
rect 862 138 866 142
rect 990 138 994 142
rect 1022 138 1026 142
rect 1086 138 1090 142
rect 1102 138 1106 142
rect 1174 138 1178 142
rect 1238 138 1242 142
rect 1310 138 1314 142
rect 1334 138 1338 142
rect 62 128 66 132
rect 126 128 130 132
rect 190 128 194 132
rect 254 128 258 132
rect 326 128 330 132
rect 358 128 362 132
rect 502 128 506 132
rect 542 128 546 132
rect 606 128 610 132
rect 646 128 650 132
rect 750 128 754 132
rect 838 128 842 132
rect 870 128 874 132
rect 918 128 922 132
rect 1030 128 1034 132
rect 1094 128 1098 132
rect 1182 128 1186 132
rect 1190 128 1194 132
rect 1318 128 1322 132
rect 1398 128 1402 132
rect 526 118 530 122
rect 582 118 586 122
rect 662 118 666 122
rect 986 103 990 107
rect 993 103 997 107
rect 22 88 26 92
rect 46 88 50 92
rect 94 88 98 92
rect 118 88 122 92
rect 142 88 146 92
rect 206 88 210 92
rect 230 88 234 92
rect 382 88 386 92
rect 422 88 426 92
rect 462 88 466 92
rect 566 88 570 92
rect 614 88 618 92
rect 662 88 666 92
rect 734 88 738 92
rect 758 88 762 92
rect 798 88 802 92
rect 910 88 914 92
rect 950 88 954 92
rect 998 88 1002 92
rect 1094 88 1098 92
rect 1118 88 1122 92
rect 1158 88 1162 92
rect 1198 88 1202 92
rect 1238 88 1242 92
rect 1350 88 1354 92
rect 1366 88 1370 92
rect 1438 88 1442 92
rect 6 78 10 82
rect 70 78 74 82
rect 166 78 170 82
rect 278 78 282 82
rect 318 78 322 82
rect 390 78 394 82
rect 398 78 402 82
rect 438 78 442 82
rect 470 78 474 82
rect 542 78 546 82
rect 574 78 578 82
rect 590 78 594 82
rect 630 78 634 82
rect 702 78 706 82
rect 710 78 714 82
rect 774 78 778 82
rect 838 78 842 82
rect 966 78 970 82
rect 1022 78 1026 82
rect 1030 78 1034 82
rect 1046 78 1050 82
rect 1142 78 1146 82
rect 1174 78 1178 82
rect 1214 78 1218 82
rect 1270 78 1274 82
rect 1406 78 1410 82
rect 1462 78 1466 82
rect 102 68 106 72
rect 110 68 114 72
rect 134 68 138 72
rect 198 68 202 72
rect 254 68 258 72
rect 270 68 274 72
rect 350 68 354 72
rect 358 68 362 72
rect 374 68 378 72
rect 446 68 450 72
rect 502 68 506 72
rect 598 68 602 72
rect 622 68 626 72
rect 654 68 658 72
rect 750 68 754 72
rect 766 68 770 72
rect 806 68 810 72
rect 838 68 842 72
rect 886 68 890 72
rect 902 68 906 72
rect 926 68 930 72
rect 934 68 938 72
rect 974 68 978 72
rect 1086 68 1090 72
rect 1102 68 1106 72
rect 1126 68 1130 72
rect 1166 68 1170 72
rect 1190 68 1194 72
rect 1222 68 1226 72
rect 1246 68 1250 72
rect 1310 68 1314 72
rect 1334 68 1338 72
rect 1358 68 1362 72
rect 62 58 66 62
rect 174 58 178 62
rect 230 58 234 62
rect 334 58 338 62
rect 342 58 346 62
rect 502 58 506 62
rect 518 58 522 62
rect 678 58 682 62
rect 814 58 818 62
rect 862 58 866 62
rect 1038 58 1042 62
rect 1046 58 1050 62
rect 1062 58 1066 62
rect 1262 58 1266 62
rect 1294 58 1298 62
rect 1382 58 1386 62
rect 1430 58 1434 62
rect 126 48 130 52
rect 214 48 218 52
rect 222 48 226 52
rect 286 48 290 52
rect 326 48 330 52
rect 518 48 522 52
rect 638 48 642 52
rect 742 48 746 52
rect 886 48 890 52
rect 910 48 914 52
rect 1086 48 1090 52
rect 1110 48 1114 52
rect 1190 48 1194 52
rect 1206 48 1210 52
rect 1262 48 1266 52
rect 1318 48 1322 52
rect 1334 48 1338 52
rect 1366 48 1370 52
rect 238 38 242 42
rect 374 38 378 42
rect 502 38 506 42
rect 1414 38 1418 42
rect 474 3 478 7
rect 481 3 485 7
<< metal2 >>
rect 142 1441 146 1442
rect 134 1438 146 1441
rect 342 1438 346 1442
rect 438 1438 442 1442
rect 518 1438 522 1442
rect 542 1438 546 1442
rect 566 1441 570 1442
rect 590 1441 594 1442
rect 558 1438 570 1441
rect 582 1438 594 1441
rect 614 1438 618 1442
rect 654 1441 658 1442
rect 654 1438 665 1441
rect 82 1358 86 1361
rect 54 1342 57 1348
rect 30 1338 38 1341
rect 90 1338 94 1341
rect 6 1332 9 1338
rect 6 1312 9 1328
rect 6 1252 9 1258
rect 6 1232 9 1248
rect 6 1092 9 1228
rect 14 1192 17 1248
rect 22 1242 25 1318
rect 30 1282 33 1338
rect 134 1332 137 1438
rect 146 1358 150 1361
rect 150 1332 153 1338
rect 166 1332 169 1388
rect 294 1362 297 1368
rect 202 1358 206 1361
rect 222 1342 225 1348
rect 238 1342 241 1358
rect 246 1352 249 1358
rect 342 1352 345 1438
rect 438 1412 441 1438
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 485 1403 488 1407
rect 518 1392 521 1438
rect 358 1362 361 1368
rect 398 1362 401 1368
rect 454 1362 457 1368
rect 394 1358 398 1361
rect 338 1348 342 1351
rect 358 1342 361 1348
rect 194 1338 198 1341
rect 258 1338 262 1341
rect 330 1338 334 1341
rect 370 1338 374 1341
rect 70 1272 73 1318
rect 34 1268 38 1271
rect 38 1192 41 1268
rect 54 1262 57 1268
rect 86 1262 89 1318
rect 102 1262 105 1268
rect 74 1258 78 1261
rect 82 1248 86 1251
rect 66 1238 70 1241
rect 46 1162 49 1198
rect 70 1172 73 1178
rect 78 1171 81 1218
rect 78 1168 89 1171
rect 22 1142 25 1148
rect 62 1132 65 1168
rect 70 1152 73 1158
rect 78 1142 81 1158
rect 78 1122 81 1138
rect 6 1072 9 1078
rect 46 1052 49 1118
rect 62 1062 65 1088
rect 86 1062 89 1168
rect 94 1142 97 1248
rect 110 1242 113 1258
rect 118 1242 121 1318
rect 134 1302 137 1328
rect 158 1262 161 1268
rect 146 1258 150 1261
rect 146 1248 150 1251
rect 174 1242 177 1318
rect 182 1282 185 1338
rect 130 1238 134 1241
rect 102 1172 105 1218
rect 126 1191 129 1218
rect 118 1188 129 1191
rect 102 1152 105 1158
rect 110 1121 113 1158
rect 118 1152 121 1188
rect 126 1172 129 1178
rect 182 1172 185 1268
rect 198 1262 201 1318
rect 222 1292 225 1338
rect 238 1322 241 1328
rect 270 1282 273 1338
rect 290 1328 294 1331
rect 322 1328 326 1331
rect 210 1258 214 1261
rect 210 1248 214 1251
rect 194 1238 198 1241
rect 130 1158 134 1161
rect 190 1152 193 1218
rect 202 1158 206 1161
rect 138 1148 142 1151
rect 102 1118 113 1121
rect 94 1062 97 1118
rect 6 1012 9 1048
rect 46 1022 49 1038
rect 6 922 9 998
rect 30 992 33 1018
rect 14 972 17 988
rect 26 978 41 981
rect 38 972 41 978
rect 30 962 33 968
rect 38 952 41 958
rect 26 948 30 951
rect 46 932 49 1018
rect 54 1002 57 1018
rect 62 1002 65 1058
rect 78 1042 81 1048
rect 86 1032 89 1038
rect 94 1012 97 1048
rect 54 942 57 998
rect 74 968 78 971
rect 86 952 89 988
rect 102 972 105 1118
rect 114 1058 118 1061
rect 134 1061 137 1118
rect 150 1112 153 1138
rect 182 1132 185 1138
rect 162 1128 166 1131
rect 190 1122 193 1138
rect 166 1072 169 1108
rect 134 1058 142 1061
rect 110 1032 113 1038
rect 98 968 102 971
rect 110 942 113 1008
rect 118 962 121 1018
rect 126 982 129 1048
rect 166 1042 169 1068
rect 182 1052 185 1058
rect 150 1032 153 1038
rect 142 952 145 958
rect 122 938 126 941
rect 58 928 62 931
rect 114 928 118 931
rect 30 882 33 888
rect 10 868 14 871
rect 22 802 25 858
rect 46 812 49 858
rect 54 852 57 868
rect 70 862 73 868
rect 78 862 81 918
rect 98 858 102 861
rect 138 858 142 861
rect 6 782 9 788
rect 6 732 9 748
rect 6 672 9 678
rect 6 582 9 608
rect 6 572 9 578
rect 6 482 9 488
rect 14 452 17 518
rect 22 392 25 658
rect 62 612 65 818
rect 86 792 89 858
rect 122 848 126 851
rect 150 851 153 1008
rect 158 962 161 1018
rect 174 972 177 1018
rect 190 1012 193 1048
rect 198 1032 201 1058
rect 206 1042 209 1118
rect 214 1052 217 1248
rect 238 1232 241 1258
rect 262 1222 265 1268
rect 246 1212 249 1218
rect 262 1142 265 1218
rect 270 1202 273 1268
rect 278 1252 281 1318
rect 334 1282 337 1288
rect 342 1282 345 1288
rect 350 1282 353 1288
rect 294 1262 297 1278
rect 302 1272 305 1278
rect 334 1262 337 1268
rect 306 1258 310 1261
rect 358 1252 361 1318
rect 374 1282 377 1338
rect 406 1332 409 1358
rect 430 1342 433 1348
rect 454 1342 457 1348
rect 498 1338 502 1341
rect 518 1331 521 1388
rect 542 1362 545 1438
rect 558 1362 561 1438
rect 574 1382 577 1388
rect 582 1371 585 1438
rect 614 1412 617 1438
rect 574 1368 585 1371
rect 526 1342 529 1348
rect 518 1328 526 1331
rect 406 1322 409 1328
rect 398 1301 401 1318
rect 398 1298 409 1301
rect 398 1282 401 1288
rect 374 1262 377 1278
rect 302 1132 305 1238
rect 366 1162 369 1258
rect 322 1138 326 1141
rect 342 1132 345 1148
rect 374 1142 377 1258
rect 382 1142 385 1188
rect 226 1128 230 1131
rect 290 1128 294 1131
rect 254 1122 257 1128
rect 230 1082 233 1088
rect 238 1062 241 1118
rect 278 1112 281 1118
rect 302 1082 305 1128
rect 326 1122 329 1128
rect 226 1058 230 1061
rect 258 1058 262 1061
rect 234 1048 238 1051
rect 198 1011 201 1018
rect 198 1008 206 1011
rect 182 962 185 968
rect 174 952 177 958
rect 162 948 166 951
rect 166 932 169 938
rect 190 932 193 948
rect 198 942 201 968
rect 214 962 217 1048
rect 270 1042 273 1068
rect 302 1052 305 1058
rect 246 1032 249 1038
rect 254 1032 257 1038
rect 310 1032 313 1118
rect 350 1102 353 1138
rect 374 1122 377 1128
rect 366 1112 369 1118
rect 322 1068 326 1071
rect 334 1042 337 1078
rect 358 1062 361 1108
rect 366 1052 369 1098
rect 374 1082 377 1118
rect 390 1072 393 1248
rect 406 1232 409 1298
rect 414 1242 417 1328
rect 526 1322 529 1328
rect 446 1272 449 1298
rect 458 1278 462 1281
rect 450 1268 454 1271
rect 426 1258 438 1261
rect 406 1142 409 1208
rect 422 1182 425 1218
rect 430 1212 433 1248
rect 462 1202 465 1268
rect 502 1262 505 1278
rect 486 1232 489 1248
rect 510 1232 513 1318
rect 534 1281 537 1358
rect 558 1352 561 1358
rect 530 1278 537 1281
rect 542 1282 545 1308
rect 558 1282 561 1318
rect 566 1282 569 1338
rect 574 1272 577 1368
rect 590 1342 593 1408
rect 622 1362 625 1368
rect 630 1352 633 1378
rect 650 1358 654 1361
rect 610 1348 622 1351
rect 582 1332 585 1338
rect 590 1321 593 1338
rect 582 1318 593 1321
rect 574 1262 577 1268
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 485 1203 488 1207
rect 430 1162 433 1198
rect 450 1158 454 1161
rect 450 1148 454 1151
rect 398 1072 401 1118
rect 406 1102 409 1138
rect 430 1122 433 1138
rect 446 1132 449 1148
rect 510 1142 513 1168
rect 534 1162 537 1218
rect 542 1162 545 1238
rect 550 1132 553 1198
rect 566 1142 569 1178
rect 574 1162 577 1258
rect 582 1252 585 1318
rect 590 1262 593 1268
rect 610 1258 614 1261
rect 622 1252 625 1328
rect 630 1272 633 1338
rect 638 1332 641 1358
rect 662 1342 665 1438
rect 694 1438 698 1442
rect 822 1438 826 1442
rect 862 1438 866 1442
rect 958 1438 962 1442
rect 1038 1438 1042 1442
rect 1062 1438 1066 1442
rect 1086 1438 1090 1442
rect 1182 1438 1186 1442
rect 1198 1438 1202 1442
rect 1214 1438 1218 1442
rect 1270 1438 1274 1442
rect 1302 1438 1306 1442
rect 1318 1438 1322 1442
rect 670 1368 678 1371
rect 670 1342 673 1368
rect 694 1362 697 1438
rect 774 1382 777 1398
rect 682 1348 686 1351
rect 650 1338 654 1341
rect 662 1322 665 1338
rect 694 1332 697 1358
rect 726 1352 729 1358
rect 742 1352 745 1378
rect 702 1322 705 1338
rect 714 1318 718 1321
rect 662 1282 665 1308
rect 670 1252 673 1278
rect 678 1252 681 1318
rect 690 1288 694 1291
rect 714 1278 718 1281
rect 582 1212 585 1248
rect 606 1232 609 1238
rect 482 1128 486 1131
rect 514 1128 518 1131
rect 422 1102 425 1118
rect 378 1068 382 1071
rect 402 1058 406 1061
rect 418 1058 422 1061
rect 370 1048 374 1051
rect 350 1042 353 1048
rect 430 1042 433 1048
rect 446 1042 449 1118
rect 454 1062 457 1068
rect 494 1062 497 1118
rect 518 1072 521 1118
rect 542 1092 545 1118
rect 550 1082 553 1128
rect 566 1082 569 1138
rect 582 1132 585 1138
rect 590 1132 593 1148
rect 598 1142 601 1218
rect 614 1172 617 1218
rect 622 1142 625 1248
rect 634 1238 638 1241
rect 710 1192 713 1228
rect 718 1192 721 1268
rect 682 1178 697 1181
rect 694 1171 697 1178
rect 726 1172 729 1328
rect 742 1282 745 1348
rect 766 1332 769 1368
rect 774 1362 777 1378
rect 774 1342 777 1348
rect 802 1338 806 1341
rect 822 1321 825 1438
rect 830 1332 833 1388
rect 842 1338 846 1341
rect 834 1328 838 1331
rect 822 1318 833 1321
rect 758 1272 761 1278
rect 734 1262 737 1268
rect 754 1258 758 1261
rect 746 1238 750 1241
rect 694 1168 702 1171
rect 654 1162 657 1168
rect 670 1162 673 1168
rect 690 1158 694 1161
rect 710 1152 713 1168
rect 654 1142 657 1148
rect 618 1128 622 1131
rect 574 1102 577 1118
rect 582 1092 585 1128
rect 678 1122 681 1148
rect 726 1142 729 1168
rect 766 1142 769 1248
rect 774 1152 777 1278
rect 782 1242 785 1318
rect 814 1272 817 1318
rect 790 1262 793 1268
rect 818 1258 822 1261
rect 830 1252 833 1318
rect 846 1281 849 1318
rect 862 1292 865 1438
rect 902 1362 905 1398
rect 958 1362 961 1438
rect 954 1358 958 1361
rect 986 1358 990 1361
rect 1018 1358 1022 1361
rect 890 1348 894 1351
rect 870 1342 873 1348
rect 870 1292 873 1328
rect 886 1292 889 1298
rect 846 1278 854 1281
rect 886 1272 889 1288
rect 894 1282 897 1338
rect 902 1332 905 1358
rect 1038 1352 1041 1438
rect 1050 1348 1054 1351
rect 930 1338 934 1341
rect 954 1338 958 1341
rect 994 1338 998 1341
rect 1006 1332 1009 1348
rect 1022 1342 1025 1348
rect 1062 1342 1065 1438
rect 946 1328 950 1331
rect 1050 1328 1054 1331
rect 1030 1322 1033 1328
rect 1062 1322 1065 1338
rect 1086 1332 1089 1438
rect 1182 1372 1185 1438
rect 1198 1412 1201 1438
rect 1214 1382 1217 1438
rect 1270 1392 1273 1438
rect 1302 1412 1305 1438
rect 1318 1402 1321 1438
rect 1190 1362 1193 1378
rect 1098 1358 1102 1361
rect 1146 1358 1150 1361
rect 1178 1358 1182 1361
rect 1106 1348 1110 1351
rect 1082 1328 1086 1331
rect 902 1282 905 1308
rect 790 1151 793 1218
rect 798 1172 801 1248
rect 814 1242 817 1248
rect 830 1242 833 1248
rect 846 1242 849 1268
rect 870 1262 873 1268
rect 858 1258 862 1261
rect 906 1248 910 1251
rect 822 1232 825 1238
rect 854 1172 857 1218
rect 826 1168 830 1171
rect 842 1168 846 1171
rect 862 1162 865 1248
rect 926 1242 929 1318
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 994 1278 998 1281
rect 966 1272 969 1278
rect 950 1262 953 1268
rect 938 1258 942 1261
rect 918 1232 921 1238
rect 942 1232 945 1248
rect 790 1148 801 1151
rect 810 1148 822 1151
rect 774 1142 777 1148
rect 790 1132 793 1138
rect 618 1118 622 1121
rect 538 1068 542 1071
rect 550 1062 553 1068
rect 534 1052 537 1058
rect 494 1042 497 1048
rect 518 1042 521 1048
rect 506 1038 510 1041
rect 574 1041 577 1088
rect 630 1082 633 1088
rect 670 1082 673 1108
rect 678 1082 681 1088
rect 630 1072 633 1078
rect 678 1072 681 1078
rect 686 1072 689 1128
rect 734 1072 737 1118
rect 742 1112 745 1128
rect 762 1118 766 1121
rect 798 1112 801 1148
rect 766 1102 769 1108
rect 742 1072 745 1088
rect 766 1082 769 1098
rect 794 1088 798 1091
rect 770 1078 774 1081
rect 782 1072 785 1078
rect 618 1068 622 1071
rect 606 1062 609 1068
rect 594 1058 598 1061
rect 602 1048 609 1051
rect 574 1038 582 1041
rect 414 1032 417 1038
rect 282 1028 286 1031
rect 358 1012 361 1018
rect 222 982 225 988
rect 234 968 238 971
rect 190 882 193 918
rect 214 882 217 958
rect 222 952 225 958
rect 246 952 249 998
rect 310 962 313 988
rect 318 962 321 998
rect 394 988 398 991
rect 330 968 334 971
rect 390 962 393 978
rect 334 952 337 958
rect 266 948 270 951
rect 290 938 294 941
rect 330 938 334 941
rect 246 872 249 908
rect 254 892 257 938
rect 262 932 265 938
rect 334 932 337 938
rect 358 932 361 938
rect 406 932 409 988
rect 422 981 425 1018
rect 454 981 457 1018
rect 494 1012 497 1038
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 485 1003 488 1007
rect 422 978 433 981
rect 454 978 465 981
rect 422 962 425 968
rect 430 952 433 978
rect 450 968 454 971
rect 438 942 441 958
rect 462 952 465 978
rect 498 968 502 971
rect 470 942 473 958
rect 510 952 513 1018
rect 558 972 561 978
rect 534 962 537 968
rect 518 942 521 958
rect 542 952 545 958
rect 550 942 553 958
rect 574 952 577 1018
rect 606 1012 609 1048
rect 686 1022 689 1068
rect 702 1062 705 1068
rect 714 1058 718 1061
rect 718 1031 721 1048
rect 742 1042 745 1048
rect 814 1042 817 1108
rect 822 1062 825 1108
rect 838 1082 841 1158
rect 858 1148 862 1151
rect 846 1112 849 1118
rect 862 1092 865 1138
rect 854 1072 857 1078
rect 854 1052 857 1058
rect 862 1052 865 1088
rect 870 1082 873 1158
rect 886 1152 889 1228
rect 898 1168 902 1171
rect 938 1168 942 1171
rect 954 1168 958 1171
rect 910 1151 913 1168
rect 966 1162 969 1228
rect 974 1202 977 1278
rect 1030 1272 1033 1318
rect 1070 1282 1073 1328
rect 1078 1312 1081 1318
rect 1090 1278 1094 1281
rect 1070 1272 1073 1278
rect 906 1148 913 1151
rect 938 1148 942 1151
rect 954 1148 958 1151
rect 918 1142 921 1148
rect 966 1142 969 1158
rect 970 1138 977 1141
rect 898 1118 902 1121
rect 910 1112 913 1128
rect 870 1052 873 1078
rect 878 1062 881 1068
rect 918 1062 921 1118
rect 958 1082 961 1108
rect 966 1082 969 1098
rect 958 1072 961 1078
rect 946 1068 950 1071
rect 934 1052 937 1058
rect 830 1042 833 1048
rect 846 1042 849 1048
rect 926 1042 929 1048
rect 730 1038 734 1041
rect 830 1032 833 1038
rect 878 1032 881 1038
rect 886 1032 889 1038
rect 718 1028 729 1031
rect 606 962 609 1008
rect 646 972 649 1018
rect 718 982 721 1018
rect 654 972 657 978
rect 618 968 622 971
rect 674 968 678 971
rect 598 952 601 958
rect 370 928 374 931
rect 186 868 190 871
rect 242 868 246 871
rect 150 848 158 851
rect 102 842 105 848
rect 166 842 169 858
rect 206 852 209 858
rect 214 852 217 858
rect 146 838 150 841
rect 110 832 113 838
rect 174 832 177 838
rect 222 832 225 858
rect 262 852 265 858
rect 270 852 273 878
rect 286 872 289 918
rect 302 862 305 918
rect 282 858 286 861
rect 314 858 318 861
rect 298 848 302 851
rect 326 841 329 898
rect 350 872 353 888
rect 358 882 361 928
rect 438 922 441 938
rect 382 902 385 918
rect 386 878 390 881
rect 390 862 393 868
rect 334 852 337 858
rect 366 852 369 858
rect 398 852 401 908
rect 410 858 414 861
rect 322 838 329 841
rect 166 822 169 828
rect 198 822 201 828
rect 230 822 233 838
rect 278 832 281 838
rect 286 832 289 838
rect 310 832 313 838
rect 218 818 222 821
rect 118 772 121 818
rect 134 761 137 818
rect 174 792 177 798
rect 134 758 145 761
rect 130 748 134 751
rect 94 742 97 747
rect 142 741 145 758
rect 138 738 145 741
rect 150 742 153 748
rect 170 738 174 741
rect 166 732 169 738
rect 94 722 97 728
rect 86 662 89 708
rect 94 682 97 718
rect 142 692 145 698
rect 150 692 153 728
rect 206 722 209 748
rect 214 741 217 808
rect 270 792 273 798
rect 298 788 302 791
rect 286 752 289 768
rect 390 762 393 848
rect 418 838 422 841
rect 430 841 433 918
rect 446 862 449 878
rect 462 852 465 918
rect 494 862 497 918
rect 510 872 513 938
rect 518 892 521 938
rect 526 872 529 918
rect 534 882 537 918
rect 550 912 553 938
rect 574 932 577 938
rect 566 882 569 928
rect 582 922 585 938
rect 562 878 566 881
rect 450 848 454 851
rect 430 838 438 841
rect 454 832 457 848
rect 486 842 489 848
rect 502 832 505 848
rect 406 822 409 828
rect 226 748 230 751
rect 214 738 225 741
rect 174 692 177 708
rect 222 692 225 738
rect 326 722 329 748
rect 350 722 353 748
rect 390 742 393 758
rect 430 752 433 818
rect 472 803 474 807
rect 478 803 481 807
rect 485 803 488 807
rect 150 682 153 688
rect 182 682 185 688
rect 214 682 217 688
rect 198 672 201 678
rect 270 672 273 718
rect 130 668 134 671
rect 162 668 166 671
rect 214 662 217 668
rect 374 662 377 738
rect 390 662 393 668
rect 186 658 190 661
rect 258 658 262 661
rect 126 652 129 658
rect 158 642 161 658
rect 374 652 377 658
rect 318 642 321 648
rect 38 542 41 568
rect 102 562 105 608
rect 126 592 129 638
rect 122 568 129 571
rect 62 532 65 538
rect 70 532 73 548
rect 30 512 33 528
rect 30 462 33 508
rect 46 462 49 468
rect 54 461 57 518
rect 54 458 62 461
rect 78 461 81 518
rect 94 512 97 538
rect 102 501 105 558
rect 114 548 118 551
rect 94 498 105 501
rect 70 458 81 461
rect 86 462 89 468
rect 42 448 46 451
rect 54 412 57 448
rect 70 442 73 458
rect 82 448 86 451
rect 86 392 89 418
rect 54 372 57 378
rect 74 368 78 371
rect 14 342 17 368
rect 30 352 33 358
rect 22 292 25 348
rect 46 322 49 368
rect 94 362 97 498
rect 126 492 129 568
rect 134 532 137 588
rect 398 581 401 718
rect 406 592 409 748
rect 414 742 417 748
rect 434 738 438 741
rect 434 728 438 731
rect 450 728 454 731
rect 466 718 470 721
rect 422 662 425 718
rect 470 662 473 688
rect 478 642 481 748
rect 494 742 497 818
rect 502 792 505 828
rect 510 812 513 868
rect 586 858 598 861
rect 606 852 609 958
rect 614 952 617 958
rect 630 952 633 958
rect 638 932 641 958
rect 646 952 649 958
rect 686 952 689 958
rect 614 872 617 888
rect 630 882 633 918
rect 638 912 641 928
rect 638 872 641 898
rect 594 848 598 851
rect 574 832 577 838
rect 534 822 537 828
rect 582 772 585 818
rect 606 792 609 848
rect 506 768 510 771
rect 622 762 625 788
rect 638 772 641 778
rect 646 762 649 918
rect 654 892 657 908
rect 662 852 665 928
rect 670 862 673 918
rect 678 842 681 888
rect 694 852 697 958
rect 702 932 705 938
rect 702 862 705 908
rect 690 848 694 851
rect 710 842 713 918
rect 726 872 729 1028
rect 734 932 737 988
rect 742 952 745 958
rect 790 952 793 998
rect 754 938 758 941
rect 766 932 769 938
rect 806 902 809 1018
rect 830 972 833 998
rect 846 962 849 1028
rect 854 962 857 968
rect 838 952 841 958
rect 846 932 849 958
rect 862 952 865 998
rect 870 972 873 1008
rect 890 948 894 951
rect 870 942 873 948
rect 814 892 817 918
rect 738 888 742 891
rect 774 872 777 878
rect 726 832 729 868
rect 742 862 745 868
rect 766 862 769 868
rect 802 858 814 861
rect 750 851 753 858
rect 746 848 753 851
rect 782 832 785 848
rect 798 832 801 838
rect 654 762 657 788
rect 630 752 633 758
rect 662 752 665 798
rect 670 772 673 818
rect 686 762 689 808
rect 694 782 697 788
rect 706 768 710 771
rect 718 771 721 818
rect 726 792 729 798
rect 734 772 737 778
rect 718 768 729 771
rect 694 752 697 768
rect 714 758 718 761
rect 726 752 729 768
rect 750 762 753 768
rect 766 752 769 758
rect 558 712 561 738
rect 566 722 569 747
rect 598 742 601 748
rect 746 738 750 741
rect 758 741 761 748
rect 782 742 785 828
rect 790 782 793 818
rect 822 772 825 918
rect 838 882 841 888
rect 878 882 881 888
rect 830 862 833 868
rect 838 862 841 878
rect 894 872 897 928
rect 902 891 905 1018
rect 910 1012 913 1038
rect 950 992 953 998
rect 914 958 918 961
rect 910 932 913 938
rect 942 932 945 988
rect 958 962 961 968
rect 974 962 977 1138
rect 982 1132 985 1178
rect 1022 1172 1025 1218
rect 1046 1192 1049 1268
rect 1086 1262 1089 1268
rect 1070 1252 1073 1258
rect 1086 1242 1089 1248
rect 1102 1212 1105 1268
rect 1110 1192 1113 1348
rect 1126 1342 1129 1358
rect 1166 1342 1169 1348
rect 1146 1338 1150 1341
rect 1166 1332 1169 1338
rect 1198 1332 1201 1368
rect 1230 1362 1233 1368
rect 1210 1358 1214 1361
rect 1242 1358 1246 1361
rect 1226 1348 1230 1351
rect 1118 1322 1121 1328
rect 1206 1322 1209 1328
rect 1138 1318 1142 1321
rect 1118 1272 1121 1278
rect 1142 1272 1145 1278
rect 1134 1242 1137 1258
rect 1142 1252 1145 1258
rect 1010 1168 1014 1171
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 1022 1082 1025 1138
rect 986 1048 990 1051
rect 970 948 974 951
rect 986 948 990 951
rect 998 932 1001 1078
rect 1006 1032 1009 1068
rect 1022 1062 1025 1068
rect 1030 1052 1033 1158
rect 1070 1132 1073 1178
rect 1134 1172 1137 1178
rect 1122 1168 1126 1171
rect 1078 1162 1081 1168
rect 1150 1161 1153 1248
rect 1158 1232 1161 1318
rect 1222 1292 1225 1348
rect 1258 1338 1262 1341
rect 1238 1332 1241 1338
rect 1270 1332 1273 1388
rect 1302 1342 1305 1348
rect 1310 1332 1313 1398
rect 1386 1368 1390 1371
rect 1418 1368 1422 1371
rect 1442 1358 1446 1361
rect 1398 1352 1401 1358
rect 1406 1352 1409 1358
rect 1362 1338 1366 1341
rect 1386 1338 1390 1341
rect 1346 1328 1350 1331
rect 1186 1278 1190 1281
rect 1166 1262 1169 1278
rect 1222 1272 1225 1288
rect 1254 1282 1257 1318
rect 1294 1312 1297 1318
rect 1318 1282 1321 1288
rect 1334 1282 1337 1318
rect 1358 1282 1361 1288
rect 1190 1252 1193 1258
rect 1238 1242 1241 1278
rect 1310 1262 1313 1268
rect 1282 1258 1294 1261
rect 1246 1252 1249 1258
rect 1258 1248 1262 1251
rect 1326 1251 1329 1278
rect 1366 1272 1369 1298
rect 1342 1262 1345 1268
rect 1374 1262 1377 1318
rect 1386 1258 1398 1261
rect 1406 1252 1409 1348
rect 1414 1342 1417 1348
rect 1326 1248 1337 1251
rect 1178 1238 1182 1241
rect 1218 1238 1222 1241
rect 1270 1232 1273 1238
rect 1286 1222 1289 1248
rect 1206 1162 1209 1168
rect 1146 1158 1153 1161
rect 1186 1158 1190 1161
rect 1114 1148 1118 1151
rect 1130 1148 1134 1151
rect 1094 1142 1097 1148
rect 1086 1132 1089 1138
rect 1142 1132 1145 1158
rect 1150 1132 1153 1148
rect 1206 1142 1209 1148
rect 1186 1138 1190 1141
rect 1062 1122 1065 1128
rect 1038 1062 1041 1068
rect 1030 1042 1033 1048
rect 1046 1042 1049 1118
rect 1086 1082 1089 1128
rect 1094 1072 1097 1128
rect 1182 1122 1185 1138
rect 1150 1082 1153 1118
rect 1174 1081 1177 1118
rect 1174 1078 1185 1081
rect 1154 1068 1158 1071
rect 1110 1062 1113 1068
rect 1174 1062 1177 1068
rect 1130 1058 1134 1061
rect 1078 1052 1081 1058
rect 1058 1048 1062 1051
rect 1146 1048 1150 1051
rect 1126 1042 1129 1048
rect 1182 1041 1185 1078
rect 1198 1072 1201 1078
rect 1214 1072 1217 1218
rect 1230 1192 1233 1208
rect 1246 1192 1249 1218
rect 1230 1152 1233 1188
rect 1278 1172 1281 1218
rect 1286 1172 1289 1178
rect 1242 1168 1246 1171
rect 1254 1152 1257 1158
rect 1246 1142 1249 1148
rect 1262 1142 1265 1158
rect 1286 1152 1289 1158
rect 1222 1132 1225 1138
rect 1294 1132 1297 1158
rect 1222 1092 1225 1128
rect 1194 1058 1198 1061
rect 1214 1052 1217 1068
rect 1254 1062 1257 1068
rect 1286 1062 1289 1068
rect 1294 1062 1297 1128
rect 1262 1052 1265 1058
rect 1294 1052 1297 1058
rect 1302 1052 1305 1248
rect 1334 1242 1337 1248
rect 1350 1232 1353 1248
rect 1310 1172 1313 1188
rect 1342 1172 1345 1218
rect 1318 1152 1321 1168
rect 1310 1082 1313 1118
rect 1182 1038 1190 1041
rect 1274 1038 1278 1041
rect 1006 1022 1009 1028
rect 1014 982 1017 1018
rect 1038 1012 1041 1018
rect 1062 992 1065 998
rect 1014 942 1017 978
rect 1054 962 1057 968
rect 1030 952 1033 958
rect 1062 952 1065 978
rect 1074 968 1078 971
rect 1086 942 1089 1038
rect 1134 1032 1137 1038
rect 1262 1031 1265 1038
rect 1262 1028 1273 1031
rect 1190 972 1193 978
rect 1254 972 1257 1018
rect 1202 968 1209 971
rect 1094 962 1097 968
rect 1106 958 1110 961
rect 1178 958 1182 961
rect 1134 952 1137 958
rect 1106 948 1110 951
rect 1194 948 1198 951
rect 1126 942 1129 948
rect 1150 942 1153 948
rect 1026 938 1030 941
rect 1050 938 1054 941
rect 1138 938 1142 941
rect 1018 928 1022 931
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 902 888 913 891
rect 902 872 905 878
rect 858 828 862 831
rect 814 742 817 748
rect 838 742 841 768
rect 846 742 849 748
rect 878 742 881 748
rect 758 738 766 741
rect 802 738 806 741
rect 862 738 870 741
rect 790 732 793 738
rect 818 728 822 731
rect 850 728 854 731
rect 882 728 886 731
rect 894 731 897 858
rect 902 842 905 848
rect 910 761 913 888
rect 934 882 937 888
rect 966 872 969 888
rect 1078 882 1081 908
rect 1174 902 1177 928
rect 1174 891 1177 898
rect 1170 888 1177 891
rect 1182 892 1185 918
rect 1150 882 1153 888
rect 1166 882 1169 888
rect 1002 878 1006 881
rect 1058 878 1062 881
rect 958 862 961 868
rect 934 852 937 858
rect 1014 852 1017 878
rect 1042 868 1046 871
rect 1030 862 1033 868
rect 1062 862 1065 868
rect 946 848 950 851
rect 1002 848 1006 851
rect 974 842 977 848
rect 1010 768 1014 771
rect 902 758 913 761
rect 902 742 905 758
rect 910 732 913 748
rect 1018 748 1022 751
rect 942 742 945 747
rect 894 728 905 731
rect 542 663 545 698
rect 558 672 561 708
rect 598 682 601 728
rect 802 718 806 721
rect 866 718 870 721
rect 614 682 617 688
rect 622 672 625 688
rect 630 672 633 718
rect 662 692 665 718
rect 830 702 833 718
rect 870 692 873 698
rect 846 682 849 688
rect 650 678 654 681
rect 722 678 726 681
rect 586 668 590 671
rect 598 662 601 668
rect 510 652 513 658
rect 438 632 441 638
rect 378 578 393 581
rect 398 578 409 581
rect 102 452 105 468
rect 114 458 118 461
rect 54 352 57 358
rect 62 282 65 358
rect 94 352 97 358
rect 70 292 73 338
rect 86 332 89 348
rect 102 342 105 448
rect 110 392 113 448
rect 126 392 129 478
rect 150 442 153 518
rect 174 512 177 538
rect 162 458 166 461
rect 170 458 174 461
rect 122 368 126 371
rect 134 362 137 388
rect 110 312 113 348
rect 118 292 121 318
rect 42 268 46 271
rect 38 262 41 268
rect 62 262 65 278
rect 94 272 97 278
rect 126 272 129 338
rect 134 282 137 358
rect 142 352 145 418
rect 166 412 169 448
rect 182 442 185 518
rect 190 472 193 568
rect 334 562 337 568
rect 282 558 286 561
rect 318 552 321 558
rect 342 552 345 578
rect 358 568 366 571
rect 390 571 393 578
rect 390 568 398 571
rect 350 552 353 558
rect 330 548 334 551
rect 306 538 310 541
rect 206 532 209 538
rect 246 532 249 538
rect 358 532 361 568
rect 406 562 409 578
rect 422 562 425 578
rect 454 572 457 618
rect 472 603 474 607
rect 478 603 481 607
rect 485 603 488 607
rect 514 568 518 571
rect 382 552 385 558
rect 370 548 374 551
rect 406 532 409 548
rect 254 522 257 528
rect 238 512 241 518
rect 198 482 201 508
rect 294 482 297 528
rect 422 502 425 548
rect 454 542 457 568
rect 430 512 433 518
rect 446 482 449 528
rect 454 492 457 528
rect 194 468 198 471
rect 262 462 265 468
rect 278 462 281 468
rect 218 458 222 461
rect 242 458 246 461
rect 166 392 169 408
rect 174 392 177 438
rect 162 368 166 371
rect 186 368 190 371
rect 150 292 153 368
rect 158 358 166 361
rect 130 268 134 271
rect 98 258 102 261
rect 6 162 9 258
rect 14 192 17 238
rect 22 222 25 258
rect 34 248 38 251
rect 70 231 73 258
rect 82 238 86 241
rect 70 228 81 231
rect 46 172 49 218
rect 78 192 81 228
rect 90 168 97 171
rect 14 142 17 148
rect 22 92 25 168
rect 70 162 73 168
rect 82 148 86 151
rect 58 138 62 141
rect 38 132 41 138
rect 58 128 62 131
rect 46 92 49 128
rect 94 92 97 168
rect 110 162 113 268
rect 158 262 161 358
rect 198 352 201 458
rect 286 452 289 478
rect 350 472 353 478
rect 382 472 385 478
rect 322 468 326 471
rect 338 468 342 471
rect 302 462 305 468
rect 350 452 353 468
rect 390 462 393 468
rect 410 458 422 461
rect 438 452 441 458
rect 226 448 230 451
rect 378 448 382 451
rect 242 438 246 441
rect 238 372 241 418
rect 294 392 297 448
rect 314 438 318 441
rect 246 362 249 388
rect 302 382 305 418
rect 222 352 225 358
rect 238 352 241 358
rect 178 348 182 351
rect 166 292 169 328
rect 198 272 201 348
rect 214 332 217 338
rect 206 292 209 308
rect 222 262 225 268
rect 154 258 158 261
rect 154 248 158 251
rect 126 232 129 248
rect 166 242 169 258
rect 190 252 193 258
rect 134 192 137 218
rect 102 152 105 158
rect 6 62 9 78
rect 46 72 49 88
rect 74 78 78 81
rect 102 72 105 78
rect 110 72 113 158
rect 122 138 126 141
rect 118 92 121 128
rect 126 82 129 128
rect 142 92 145 168
rect 158 162 161 168
rect 154 148 158 151
rect 166 142 169 148
rect 174 142 177 238
rect 198 222 201 258
rect 246 252 249 358
rect 286 352 289 358
rect 326 342 329 378
rect 254 332 257 338
rect 350 332 353 448
rect 358 442 361 448
rect 418 438 422 441
rect 430 432 433 438
rect 382 392 385 418
rect 370 368 374 371
rect 358 362 361 368
rect 394 358 398 361
rect 386 348 390 351
rect 402 348 406 351
rect 414 342 417 378
rect 446 352 449 478
rect 454 432 457 438
rect 462 422 465 458
rect 474 448 478 451
rect 472 403 474 407
rect 478 403 481 407
rect 485 403 488 407
rect 494 362 497 558
rect 502 552 505 568
rect 510 462 513 518
rect 518 452 521 548
rect 526 532 529 588
rect 554 568 558 571
rect 534 482 537 488
rect 534 462 537 468
rect 502 392 505 438
rect 510 372 513 418
rect 362 338 366 341
rect 422 332 425 338
rect 314 328 318 331
rect 286 322 289 328
rect 302 282 305 328
rect 326 322 329 328
rect 278 262 281 268
rect 302 262 305 268
rect 258 258 262 261
rect 310 252 313 288
rect 374 282 377 328
rect 422 292 425 328
rect 430 322 433 328
rect 462 292 465 338
rect 406 282 409 288
rect 378 278 382 281
rect 414 272 417 278
rect 326 262 329 268
rect 334 262 337 268
rect 374 262 377 268
rect 470 262 473 298
rect 478 292 481 358
rect 518 352 521 448
rect 534 442 537 448
rect 534 392 537 428
rect 526 372 529 378
rect 542 372 545 498
rect 550 482 553 498
rect 558 481 561 538
rect 566 522 569 528
rect 558 478 566 481
rect 550 442 553 468
rect 566 462 569 478
rect 558 392 561 448
rect 574 392 577 658
rect 582 552 585 558
rect 582 522 585 528
rect 582 452 585 508
rect 590 492 593 528
rect 598 451 601 638
rect 614 562 617 568
rect 622 552 625 558
rect 614 532 617 538
rect 606 462 609 468
rect 622 452 625 458
rect 598 448 609 451
rect 606 392 609 448
rect 582 372 585 378
rect 614 372 617 398
rect 542 362 545 368
rect 566 362 569 368
rect 598 362 601 368
rect 622 362 625 448
rect 630 432 633 658
rect 638 592 641 678
rect 682 668 686 671
rect 654 652 657 658
rect 690 648 694 651
rect 682 638 686 641
rect 702 632 705 638
rect 646 572 649 588
rect 638 542 641 568
rect 662 562 665 578
rect 718 572 721 678
rect 782 672 785 678
rect 726 622 729 668
rect 766 652 769 658
rect 742 642 745 648
rect 758 632 761 638
rect 734 572 737 588
rect 686 542 689 568
rect 742 562 745 578
rect 750 562 753 578
rect 766 572 769 618
rect 774 582 777 648
rect 790 622 793 668
rect 806 662 809 668
rect 826 658 830 661
rect 818 638 822 641
rect 830 632 833 648
rect 774 562 777 578
rect 798 572 801 578
rect 806 572 809 578
rect 814 562 817 628
rect 830 602 833 618
rect 838 592 841 638
rect 718 552 721 558
rect 738 548 742 551
rect 806 542 809 548
rect 698 538 702 541
rect 762 538 766 541
rect 786 538 790 541
rect 646 532 649 538
rect 658 518 662 521
rect 678 492 681 518
rect 734 502 737 518
rect 734 482 737 498
rect 742 482 745 508
rect 642 478 646 481
rect 642 468 646 471
rect 694 471 697 478
rect 694 468 702 471
rect 746 468 750 471
rect 662 462 665 468
rect 674 458 678 461
rect 666 448 670 451
rect 686 442 689 448
rect 670 392 673 398
rect 678 381 681 418
rect 694 392 697 468
rect 758 462 761 528
rect 790 482 793 508
rect 778 468 782 471
rect 806 462 809 478
rect 754 448 758 451
rect 778 448 782 451
rect 702 442 705 448
rect 742 392 745 438
rect 790 422 793 458
rect 782 392 785 398
rect 670 378 681 381
rect 638 372 641 378
rect 650 368 657 371
rect 510 342 513 348
rect 534 292 537 348
rect 550 342 553 348
rect 574 342 577 348
rect 606 342 609 348
rect 558 302 561 318
rect 558 282 561 288
rect 546 278 550 281
rect 514 268 518 271
rect 442 258 446 261
rect 238 248 246 251
rect 338 248 342 251
rect 206 192 209 238
rect 238 172 241 248
rect 266 238 270 241
rect 322 238 326 241
rect 194 158 198 161
rect 158 88 166 91
rect 134 72 137 78
rect 98 68 102 71
rect 62 12 65 58
rect 130 48 134 51
rect 86 -18 89 8
rect 158 -18 161 88
rect 166 82 169 88
rect 182 82 185 138
rect 190 122 193 128
rect 198 102 201 158
rect 206 92 209 168
rect 218 148 230 151
rect 246 151 249 238
rect 254 232 257 238
rect 270 192 273 218
rect 282 168 286 171
rect 262 162 265 168
rect 294 162 297 168
rect 326 162 329 168
rect 270 152 273 158
rect 246 148 254 151
rect 242 138 246 141
rect 198 72 201 78
rect 174 62 177 68
rect 214 52 217 108
rect 222 52 225 98
rect 230 92 233 138
rect 254 132 257 148
rect 294 142 297 148
rect 294 132 297 138
rect 326 132 329 148
rect 350 132 353 258
rect 398 252 401 258
rect 378 248 382 251
rect 450 238 454 241
rect 358 142 361 218
rect 382 192 385 228
rect 370 158 374 161
rect 382 132 385 148
rect 390 142 393 198
rect 438 192 441 238
rect 462 192 465 258
rect 470 252 473 258
rect 490 248 494 251
rect 534 242 537 258
rect 542 252 545 258
rect 554 238 561 241
rect 472 203 474 207
rect 478 203 481 207
rect 485 203 488 207
rect 558 192 561 238
rect 566 202 569 268
rect 582 252 585 278
rect 594 268 598 271
rect 606 262 609 278
rect 622 271 625 358
rect 630 352 633 358
rect 638 342 641 348
rect 654 341 657 368
rect 662 352 665 358
rect 670 352 673 378
rect 682 368 686 371
rect 654 338 665 341
rect 630 292 633 338
rect 614 268 625 271
rect 614 252 617 268
rect 630 262 633 268
rect 622 252 625 258
rect 578 238 598 241
rect 538 188 542 191
rect 422 168 430 171
rect 398 162 401 168
rect 414 132 417 158
rect 274 78 278 81
rect 258 68 262 71
rect 230 62 233 68
rect 242 38 246 41
rect 270 -18 273 68
rect 286 42 289 48
rect 318 32 321 78
rect 326 52 329 68
rect 342 62 345 78
rect 350 72 353 78
rect 358 72 361 128
rect 382 92 385 108
rect 422 92 425 168
rect 454 162 457 178
rect 474 168 481 171
rect 442 158 446 161
rect 442 148 449 151
rect 446 122 449 148
rect 438 112 441 118
rect 438 82 441 108
rect 462 92 465 148
rect 470 82 473 88
rect 370 68 374 71
rect 334 52 337 58
rect 374 42 377 48
rect 390 22 393 78
rect 398 62 401 78
rect 374 -18 377 8
rect 86 -22 90 -18
rect 158 -22 162 -18
rect 270 -22 274 -18
rect 374 -22 378 -18
rect 438 -19 441 78
rect 446 72 449 78
rect 478 52 481 168
rect 490 138 494 141
rect 502 82 505 128
rect 502 72 505 78
rect 518 62 521 178
rect 546 158 550 161
rect 542 132 545 138
rect 530 118 534 121
rect 542 82 545 88
rect 502 52 505 58
rect 514 48 518 51
rect 494 41 497 48
rect 494 38 502 41
rect 472 3 474 7
rect 478 3 481 7
rect 485 3 488 7
rect 534 -18 537 58
rect 446 -19 450 -18
rect 438 -22 450 -19
rect 534 -22 538 -18
rect 550 -19 553 158
rect 558 122 561 148
rect 566 92 569 168
rect 578 118 582 121
rect 590 82 593 198
rect 574 22 577 78
rect 598 72 601 218
rect 614 172 617 248
rect 622 192 625 238
rect 638 192 641 238
rect 606 142 609 168
rect 614 162 617 168
rect 614 148 622 151
rect 606 92 609 128
rect 614 92 617 148
rect 630 122 633 168
rect 646 152 649 328
rect 662 292 665 338
rect 678 282 681 288
rect 654 162 657 268
rect 694 262 697 268
rect 710 262 713 348
rect 718 322 721 328
rect 718 282 721 318
rect 742 292 745 368
rect 790 358 798 361
rect 782 352 785 358
rect 750 342 753 348
rect 774 332 777 348
rect 758 312 761 328
rect 754 278 758 281
rect 774 272 777 328
rect 790 292 793 358
rect 806 352 809 458
rect 814 382 817 558
rect 830 512 833 568
rect 838 552 841 568
rect 830 452 833 488
rect 846 481 849 618
rect 862 592 865 658
rect 886 652 889 658
rect 874 638 878 641
rect 886 631 889 638
rect 878 628 889 631
rect 878 592 881 628
rect 894 612 897 718
rect 902 652 905 728
rect 910 692 913 718
rect 926 712 929 738
rect 1030 732 1033 758
rect 1046 752 1049 858
rect 1062 762 1065 838
rect 1078 772 1081 878
rect 1158 872 1161 878
rect 1190 872 1193 938
rect 1206 892 1209 968
rect 1214 952 1217 958
rect 1226 938 1230 941
rect 1238 932 1241 948
rect 1230 882 1233 888
rect 1226 878 1230 881
rect 1238 872 1241 928
rect 1246 892 1249 958
rect 1258 948 1262 951
rect 1254 932 1257 938
rect 1262 882 1265 898
rect 1270 892 1273 1028
rect 1286 952 1289 1018
rect 1302 1002 1305 1048
rect 1310 1042 1313 1058
rect 1318 1042 1321 1048
rect 1298 968 1302 971
rect 1310 952 1313 1018
rect 1326 962 1329 1158
rect 1350 1152 1353 1188
rect 1358 1162 1361 1178
rect 1366 1162 1369 1228
rect 1390 1222 1393 1248
rect 1402 1238 1406 1241
rect 1386 1188 1390 1191
rect 1398 1172 1401 1218
rect 1358 1152 1361 1158
rect 1366 1142 1369 1158
rect 1386 1148 1390 1151
rect 1334 1052 1337 1138
rect 1414 1131 1417 1318
rect 1426 1258 1430 1261
rect 1422 1142 1425 1248
rect 1438 1242 1441 1278
rect 1446 1262 1449 1328
rect 1430 1172 1433 1218
rect 1434 1148 1438 1151
rect 1406 1128 1417 1131
rect 1374 1122 1377 1128
rect 1342 1092 1345 1118
rect 1390 1072 1393 1078
rect 1366 1062 1369 1068
rect 1346 1058 1350 1061
rect 1334 1012 1337 1048
rect 1354 1038 1358 1041
rect 1342 1032 1345 1038
rect 1382 1022 1385 1068
rect 1398 1002 1401 1078
rect 1406 1052 1409 1128
rect 1414 1092 1417 1118
rect 1438 1101 1441 1118
rect 1446 1112 1449 1258
rect 1454 1152 1457 1208
rect 1430 1098 1441 1101
rect 1398 992 1401 998
rect 1358 972 1361 978
rect 1346 968 1350 971
rect 1354 958 1358 961
rect 1278 928 1286 931
rect 1278 912 1281 928
rect 1286 872 1289 908
rect 1298 878 1302 881
rect 1106 868 1110 871
rect 1234 868 1238 871
rect 1258 868 1262 871
rect 1086 862 1089 868
rect 1122 858 1126 861
rect 1098 848 1102 851
rect 1170 848 1174 851
rect 1254 842 1257 848
rect 1278 832 1281 848
rect 1254 792 1257 798
rect 1118 772 1121 778
rect 1294 762 1297 818
rect 1310 792 1313 918
rect 1318 912 1321 958
rect 1366 952 1369 978
rect 1378 968 1385 971
rect 1394 968 1398 971
rect 1330 948 1334 951
rect 1322 858 1326 861
rect 1326 822 1329 828
rect 1094 752 1097 758
rect 1078 742 1081 748
rect 1126 742 1129 758
rect 1302 752 1305 758
rect 1178 748 1182 751
rect 1314 748 1318 751
rect 1262 742 1265 748
rect 1278 742 1281 748
rect 1286 742 1289 748
rect 1334 742 1337 918
rect 1350 872 1353 938
rect 1382 892 1385 968
rect 1414 942 1417 1088
rect 1430 1082 1433 1098
rect 1462 1092 1465 1338
rect 1438 1082 1441 1088
rect 1430 1072 1433 1078
rect 1426 1038 1430 1041
rect 1446 1032 1449 1068
rect 1430 962 1433 1008
rect 1442 978 1446 981
rect 1442 968 1446 971
rect 1394 938 1398 941
rect 1414 872 1417 938
rect 1422 932 1425 958
rect 1442 948 1446 951
rect 1422 892 1425 928
rect 1438 882 1441 898
rect 1370 868 1374 871
rect 1442 868 1446 871
rect 1350 862 1353 868
rect 1414 862 1417 868
rect 1398 852 1401 858
rect 1438 852 1441 858
rect 1362 848 1366 851
rect 1438 782 1441 788
rect 1350 751 1353 758
rect 1058 738 1062 741
rect 1090 738 1094 741
rect 1314 738 1318 741
rect 1134 732 1137 738
rect 1446 732 1449 868
rect 1462 842 1465 848
rect 1454 742 1457 808
rect 1470 792 1473 948
rect 1478 852 1481 868
rect 1066 728 1070 731
rect 1098 728 1102 731
rect 1258 728 1262 731
rect 1290 728 1294 731
rect 926 672 929 708
rect 942 692 945 728
rect 1166 722 1169 728
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 1022 672 1025 678
rect 1118 672 1121 678
rect 1166 672 1169 718
rect 1222 682 1225 688
rect 1246 672 1249 678
rect 1038 663 1041 668
rect 1138 659 1142 662
rect 910 592 913 658
rect 934 652 937 658
rect 942 652 945 658
rect 966 652 969 658
rect 974 652 977 658
rect 1102 652 1105 658
rect 930 648 934 651
rect 954 638 958 641
rect 986 638 990 641
rect 974 632 977 638
rect 1022 592 1025 638
rect 854 552 857 558
rect 862 542 865 548
rect 870 502 873 568
rect 886 552 889 568
rect 910 552 913 578
rect 942 572 945 578
rect 886 542 889 548
rect 842 478 849 481
rect 886 472 889 478
rect 838 452 841 468
rect 846 372 849 468
rect 862 462 865 468
rect 894 462 897 488
rect 874 458 878 461
rect 902 452 905 548
rect 910 492 913 538
rect 918 472 921 568
rect 934 492 937 558
rect 950 552 953 568
rect 942 542 945 548
rect 966 542 969 548
rect 978 538 982 541
rect 1006 541 1009 588
rect 1058 578 1062 581
rect 1014 562 1017 568
rect 1022 552 1025 578
rect 1058 568 1062 571
rect 1030 542 1033 568
rect 1042 558 1046 561
rect 1058 548 1062 551
rect 1006 538 1017 541
rect 942 492 945 498
rect 958 492 961 508
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 1006 492 1009 528
rect 986 478 990 481
rect 910 462 913 468
rect 934 462 937 468
rect 974 462 977 468
rect 1014 462 1017 538
rect 1038 482 1041 488
rect 1046 482 1049 488
rect 946 448 950 451
rect 874 438 878 441
rect 870 392 873 428
rect 902 412 905 448
rect 958 441 961 448
rect 950 438 961 441
rect 898 368 902 371
rect 846 342 849 348
rect 818 338 822 341
rect 834 338 838 341
rect 862 332 865 368
rect 910 362 913 438
rect 918 432 921 438
rect 934 392 937 438
rect 950 402 953 438
rect 922 368 926 371
rect 870 342 873 348
rect 818 328 822 331
rect 806 312 809 328
rect 822 292 825 318
rect 794 278 798 281
rect 830 272 833 328
rect 846 292 849 328
rect 730 268 734 271
rect 810 268 814 271
rect 730 258 734 261
rect 670 212 673 248
rect 678 162 681 198
rect 694 192 697 258
rect 710 162 713 218
rect 726 192 729 228
rect 734 182 737 258
rect 774 252 777 258
rect 750 212 753 248
rect 782 181 785 268
rect 794 248 798 251
rect 862 242 865 278
rect 870 272 873 278
rect 878 202 881 358
rect 894 322 897 348
rect 902 332 905 338
rect 894 292 897 298
rect 910 292 913 358
rect 942 351 945 368
rect 958 362 961 408
rect 966 362 969 368
rect 974 362 977 458
rect 1038 392 1041 418
rect 1062 362 1065 408
rect 1070 392 1073 648
rect 1078 552 1081 558
rect 1134 551 1137 608
rect 1166 552 1169 668
rect 1198 662 1201 668
rect 1206 652 1209 658
rect 1246 652 1249 658
rect 1254 652 1257 698
rect 1286 682 1289 728
rect 1350 722 1353 728
rect 1350 682 1353 718
rect 1310 672 1313 678
rect 1274 668 1278 671
rect 1298 668 1302 671
rect 1474 668 1478 671
rect 1262 662 1265 668
rect 1350 663 1353 668
rect 1418 658 1422 661
rect 1246 592 1249 638
rect 1254 592 1257 648
rect 1286 622 1289 628
rect 1318 612 1321 658
rect 1446 652 1449 658
rect 1414 642 1417 648
rect 1286 592 1289 608
rect 1222 572 1225 578
rect 1278 572 1281 578
rect 1258 568 1262 571
rect 1094 532 1097 538
rect 1094 492 1097 528
rect 1102 482 1105 528
rect 1158 492 1161 538
rect 1174 482 1177 508
rect 1190 492 1193 568
rect 1198 552 1201 568
rect 1214 532 1217 568
rect 1222 552 1225 558
rect 1238 542 1241 558
rect 1246 552 1249 558
rect 1238 492 1241 528
rect 1270 492 1273 568
rect 1294 562 1297 588
rect 1366 551 1369 618
rect 1398 552 1401 638
rect 1438 632 1441 638
rect 1286 542 1289 548
rect 1442 548 1446 551
rect 1478 542 1481 548
rect 1302 502 1305 538
rect 1286 482 1289 498
rect 1302 482 1305 498
rect 1138 478 1142 481
rect 1078 472 1081 478
rect 1206 472 1209 478
rect 1230 472 1233 478
rect 1090 468 1094 471
rect 1130 468 1134 471
rect 1306 468 1310 471
rect 1150 462 1153 468
rect 1262 462 1265 468
rect 1254 458 1262 461
rect 1078 442 1081 448
rect 1102 442 1105 458
rect 1110 452 1113 458
rect 1226 448 1230 451
rect 1090 438 1094 441
rect 1082 368 1086 371
rect 1022 358 1030 361
rect 938 348 945 351
rect 950 342 953 348
rect 1002 338 1006 341
rect 1014 332 1017 348
rect 918 282 921 328
rect 926 278 934 281
rect 942 272 945 278
rect 906 268 910 271
rect 930 268 934 271
rect 914 258 918 261
rect 798 192 801 198
rect 894 192 897 208
rect 934 202 937 268
rect 942 258 950 261
rect 782 178 793 181
rect 738 168 742 171
rect 778 168 782 171
rect 718 162 721 168
rect 790 162 793 178
rect 798 162 801 168
rect 646 132 649 148
rect 678 142 681 158
rect 714 148 726 151
rect 622 72 625 78
rect 598 22 601 68
rect 630 62 633 78
rect 582 -18 585 18
rect 598 -18 601 8
rect 622 -18 625 48
rect 638 42 641 48
rect 638 -18 641 18
rect 646 12 649 128
rect 694 122 697 138
rect 666 118 670 121
rect 734 92 737 158
rect 822 152 825 178
rect 878 162 881 168
rect 846 152 849 158
rect 810 148 814 151
rect 662 82 665 88
rect 658 68 662 71
rect 678 62 681 68
rect 702 62 705 78
rect 710 32 713 78
rect 742 52 745 128
rect 750 92 753 128
rect 758 92 761 148
rect 782 122 785 138
rect 766 72 769 118
rect 798 92 801 128
rect 838 122 841 128
rect 862 102 865 138
rect 894 132 897 148
rect 870 122 873 128
rect 910 92 913 178
rect 918 132 921 138
rect 926 82 929 198
rect 942 192 945 258
rect 958 252 961 258
rect 974 242 977 318
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 982 272 985 278
rect 982 252 985 258
rect 1006 252 1009 298
rect 1022 292 1025 358
rect 1142 352 1145 358
rect 1058 348 1062 351
rect 1106 348 1110 351
rect 1030 342 1033 348
rect 1030 282 1033 328
rect 1078 292 1081 348
rect 1122 338 1126 341
rect 1094 332 1097 338
rect 1114 328 1118 331
rect 1146 328 1150 331
rect 1030 272 1033 278
rect 1038 262 1041 278
rect 1014 242 1017 248
rect 958 192 961 208
rect 966 172 969 178
rect 994 168 998 171
rect 934 162 937 168
rect 954 158 958 161
rect 974 152 977 168
rect 982 162 985 168
rect 946 148 969 151
rect 966 141 969 148
rect 966 138 990 141
rect 950 92 953 128
rect 998 121 1001 148
rect 998 118 1009 121
rect 966 82 969 108
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 998 82 1001 88
rect 842 78 846 81
rect 774 72 777 78
rect 926 72 929 78
rect 754 68 758 71
rect 810 68 814 71
rect 834 68 838 71
rect 898 68 902 71
rect 862 62 865 68
rect 886 62 889 68
rect 934 62 937 68
rect 742 22 745 48
rect 814 12 817 58
rect 910 52 913 58
rect 886 42 889 48
rect 662 -18 665 8
rect 910 -18 913 8
rect 942 -18 945 78
rect 970 68 974 71
rect 1006 -18 1009 118
rect 558 -19 562 -18
rect 550 -22 562 -19
rect 582 -22 586 -18
rect 598 -22 602 -18
rect 622 -22 626 -18
rect 638 -22 642 -18
rect 662 -22 666 -18
rect 910 -22 914 -18
rect 942 -22 946 -18
rect 1006 -22 1010 -18
rect 1014 -19 1017 238
rect 1038 202 1041 258
rect 1046 212 1049 268
rect 1070 252 1073 288
rect 1142 282 1145 328
rect 1130 278 1134 281
rect 1102 262 1105 268
rect 1078 252 1081 258
rect 1058 248 1062 251
rect 1046 192 1049 208
rect 1046 172 1049 178
rect 1070 172 1073 248
rect 1086 242 1089 248
rect 1102 242 1105 248
rect 1150 212 1153 268
rect 1158 222 1161 338
rect 1166 312 1169 448
rect 1214 392 1217 448
rect 1238 432 1241 448
rect 1190 362 1193 368
rect 1206 362 1209 378
rect 1242 368 1246 371
rect 1254 362 1257 458
rect 1274 448 1278 451
rect 1290 448 1294 451
rect 1318 442 1321 518
rect 1334 512 1337 528
rect 1430 512 1433 518
rect 1382 482 1385 498
rect 1330 478 1334 481
rect 1342 462 1345 478
rect 1382 472 1385 478
rect 1462 472 1465 488
rect 1470 472 1473 478
rect 1334 452 1337 458
rect 1362 448 1366 451
rect 1278 392 1281 428
rect 1302 392 1305 438
rect 1350 432 1353 438
rect 1374 422 1377 428
rect 1310 372 1313 398
rect 1334 392 1337 418
rect 1342 372 1345 418
rect 1382 382 1385 468
rect 1390 462 1393 468
rect 1426 458 1430 461
rect 1446 452 1449 458
rect 1426 438 1430 441
rect 1270 362 1273 368
rect 1358 362 1361 368
rect 1366 362 1369 378
rect 1398 372 1401 418
rect 1374 362 1377 368
rect 1226 358 1230 361
rect 1298 358 1302 361
rect 1174 352 1177 358
rect 1194 348 1198 351
rect 1198 332 1201 338
rect 1190 292 1193 328
rect 1206 302 1209 358
rect 1242 348 1246 351
rect 1222 322 1225 328
rect 1166 252 1169 258
rect 1174 232 1177 278
rect 1206 262 1209 268
rect 1190 252 1193 258
rect 1182 222 1185 228
rect 1126 182 1129 188
rect 1110 172 1113 178
rect 1034 168 1038 171
rect 1130 168 1134 171
rect 1054 152 1057 168
rect 1062 162 1065 168
rect 1138 158 1142 161
rect 1022 142 1025 148
rect 1030 122 1033 128
rect 1022 91 1025 118
rect 1030 112 1033 118
rect 1022 88 1033 91
rect 1030 82 1033 88
rect 1042 78 1046 81
rect 1022 32 1025 78
rect 1062 62 1065 148
rect 1102 142 1105 158
rect 1158 152 1161 158
rect 1146 148 1150 151
rect 1086 132 1089 138
rect 1086 102 1089 128
rect 1094 122 1097 128
rect 1094 92 1097 108
rect 1118 92 1121 118
rect 1158 92 1161 128
rect 1166 122 1169 168
rect 1182 152 1185 198
rect 1214 192 1217 308
rect 1222 292 1225 318
rect 1230 272 1233 278
rect 1230 252 1233 258
rect 1238 252 1241 298
rect 1246 292 1249 328
rect 1174 92 1177 138
rect 1182 132 1185 148
rect 1190 132 1193 138
rect 1138 78 1142 81
rect 1082 68 1086 71
rect 1098 68 1102 71
rect 1122 68 1126 71
rect 1034 58 1038 61
rect 1050 58 1054 61
rect 1022 -19 1026 -18
rect 1014 -22 1026 -19
rect 1054 -19 1058 -18
rect 1062 -19 1065 58
rect 1086 52 1089 58
rect 1110 52 1113 58
rect 1054 -22 1065 -19
rect 1134 -18 1137 78
rect 1162 68 1166 71
rect 1174 32 1177 78
rect 1190 72 1193 108
rect 1198 92 1201 178
rect 1210 148 1214 151
rect 1222 132 1225 238
rect 1246 232 1249 248
rect 1254 192 1257 358
rect 1286 352 1289 358
rect 1262 272 1265 318
rect 1262 262 1265 268
rect 1270 252 1273 348
rect 1278 342 1281 348
rect 1302 332 1305 348
rect 1310 292 1313 338
rect 1278 262 1281 268
rect 1294 262 1297 268
rect 1306 258 1310 261
rect 1318 252 1321 358
rect 1326 352 1329 358
rect 1334 352 1337 358
rect 1370 348 1374 351
rect 1326 341 1329 348
rect 1390 342 1393 348
rect 1326 338 1337 341
rect 1334 292 1337 338
rect 1342 272 1345 308
rect 1358 292 1361 328
rect 1382 292 1385 318
rect 1358 262 1361 278
rect 1398 271 1401 368
rect 1406 342 1409 388
rect 1422 381 1425 418
rect 1430 392 1433 398
rect 1422 378 1433 381
rect 1414 332 1417 378
rect 1422 362 1425 368
rect 1430 352 1433 378
rect 1414 322 1417 328
rect 1422 292 1425 318
rect 1438 292 1441 368
rect 1446 358 1454 361
rect 1446 281 1449 358
rect 1454 342 1457 348
rect 1470 322 1473 338
rect 1438 278 1449 281
rect 1398 268 1409 271
rect 1398 242 1401 258
rect 1278 192 1281 238
rect 1310 222 1313 238
rect 1358 192 1361 228
rect 1366 192 1369 238
rect 1238 142 1241 148
rect 1186 68 1190 71
rect 1214 62 1217 78
rect 1222 72 1225 98
rect 1238 92 1241 98
rect 1190 52 1193 58
rect 1206 52 1209 58
rect 1150 -18 1153 8
rect 1174 -18 1177 28
rect 1222 -18 1225 68
rect 1246 62 1249 68
rect 1254 22 1257 158
rect 1270 122 1273 168
rect 1286 162 1289 188
rect 1358 162 1361 188
rect 1374 172 1377 178
rect 1394 168 1398 171
rect 1406 162 1409 268
rect 1430 232 1433 268
rect 1298 158 1302 161
rect 1278 152 1281 158
rect 1350 152 1353 158
rect 1362 148 1366 151
rect 1310 142 1313 148
rect 1318 112 1321 128
rect 1334 92 1337 138
rect 1350 92 1353 118
rect 1366 92 1369 108
rect 1262 62 1265 68
rect 1270 52 1273 78
rect 1358 72 1361 78
rect 1350 68 1358 71
rect 1298 58 1302 61
rect 1310 52 1313 68
rect 1334 62 1337 68
rect 1330 48 1334 51
rect 1262 21 1265 48
rect 1258 18 1265 21
rect 1254 -18 1257 18
rect 1270 -18 1273 48
rect 1318 42 1321 48
rect 1318 -18 1321 38
rect 1350 -18 1353 68
rect 1382 62 1385 158
rect 1402 148 1406 151
rect 1394 128 1398 131
rect 1406 82 1409 138
rect 1414 122 1417 168
rect 1422 162 1425 218
rect 1430 192 1433 218
rect 1430 162 1433 178
rect 1422 148 1430 151
rect 1422 132 1425 148
rect 1430 62 1433 118
rect 1438 92 1441 278
rect 1446 112 1449 248
rect 1462 82 1465 288
rect 1362 48 1366 51
rect 1414 42 1417 48
rect 1134 -22 1138 -18
rect 1150 -22 1154 -18
rect 1174 -22 1178 -18
rect 1222 -22 1226 -18
rect 1254 -22 1258 -18
rect 1270 -22 1274 -18
rect 1318 -22 1322 -18
rect 1350 -22 1354 -18
<< m3contact >>
rect 86 1358 90 1362
rect 54 1348 58 1352
rect 38 1338 42 1342
rect 86 1338 90 1342
rect 6 1328 10 1332
rect 6 1308 10 1312
rect 6 1248 10 1252
rect 14 1248 18 1252
rect 6 1228 10 1232
rect 166 1388 170 1392
rect 142 1358 146 1362
rect 294 1368 298 1372
rect 206 1358 210 1362
rect 238 1358 242 1362
rect 246 1358 250 1362
rect 438 1408 442 1412
rect 474 1403 478 1407
rect 481 1403 485 1407
rect 518 1388 522 1392
rect 358 1368 362 1372
rect 398 1368 402 1372
rect 454 1368 458 1372
rect 390 1358 394 1362
rect 406 1358 410 1362
rect 342 1348 346 1352
rect 182 1338 186 1342
rect 198 1338 202 1342
rect 222 1338 226 1342
rect 254 1338 258 1342
rect 334 1338 338 1342
rect 358 1338 362 1342
rect 366 1338 370 1342
rect 150 1328 154 1332
rect 38 1268 42 1272
rect 54 1268 58 1272
rect 70 1268 74 1272
rect 22 1238 26 1242
rect 102 1268 106 1272
rect 70 1258 74 1262
rect 86 1258 90 1262
rect 110 1258 114 1262
rect 78 1248 82 1252
rect 62 1238 66 1242
rect 46 1198 50 1202
rect 38 1188 42 1192
rect 70 1168 74 1172
rect 22 1138 26 1142
rect 70 1158 74 1162
rect 78 1138 82 1142
rect 62 1128 66 1132
rect 78 1118 82 1122
rect 6 1088 10 1092
rect 6 1078 10 1082
rect 62 1088 66 1092
rect 134 1298 138 1302
rect 158 1268 162 1272
rect 150 1258 154 1262
rect 142 1248 146 1252
rect 118 1238 122 1242
rect 126 1238 130 1242
rect 174 1238 178 1242
rect 102 1158 106 1162
rect 110 1158 114 1162
rect 94 1138 98 1142
rect 126 1178 130 1182
rect 238 1318 242 1322
rect 286 1328 290 1332
rect 326 1328 330 1332
rect 270 1278 274 1282
rect 198 1258 202 1262
rect 214 1258 218 1262
rect 206 1248 210 1252
rect 190 1238 194 1242
rect 182 1168 186 1172
rect 126 1158 130 1162
rect 198 1158 202 1162
rect 118 1148 122 1152
rect 142 1148 146 1152
rect 190 1148 194 1152
rect 94 1058 98 1062
rect 6 1048 10 1052
rect 46 1048 50 1052
rect 46 1038 50 1042
rect 54 1018 58 1022
rect 6 1008 10 1012
rect 6 998 10 1002
rect 14 988 18 992
rect 30 988 34 992
rect 30 968 34 972
rect 38 968 42 972
rect 38 958 42 962
rect 30 948 34 952
rect 78 1048 82 1052
rect 86 1028 90 1032
rect 94 1008 98 1012
rect 54 998 58 1002
rect 62 998 66 1002
rect 86 988 90 992
rect 70 968 74 972
rect 110 1058 114 1062
rect 166 1128 170 1132
rect 182 1128 186 1132
rect 190 1118 194 1122
rect 150 1108 154 1112
rect 166 1108 170 1112
rect 110 1028 114 1032
rect 110 1008 114 1012
rect 102 968 106 972
rect 182 1058 186 1062
rect 166 1038 170 1042
rect 150 1028 154 1032
rect 150 1008 154 1012
rect 126 978 130 982
rect 118 958 122 962
rect 142 958 146 962
rect 126 938 130 942
rect 46 928 50 932
rect 54 928 58 932
rect 110 928 114 932
rect 6 918 10 922
rect 30 878 34 882
rect 14 868 18 872
rect 70 858 74 862
rect 78 858 82 862
rect 94 858 98 862
rect 142 858 146 862
rect 54 848 58 852
rect 46 808 50 812
rect 22 798 26 802
rect 6 788 10 792
rect 6 748 10 752
rect 6 728 10 732
rect 6 678 10 682
rect 22 658 26 662
rect 6 608 10 612
rect 6 578 10 582
rect 6 488 10 492
rect 14 448 18 452
rect 102 848 106 852
rect 118 848 122 852
rect 238 1228 242 1232
rect 262 1218 266 1222
rect 246 1208 250 1212
rect 334 1288 338 1292
rect 342 1288 346 1292
rect 350 1288 354 1292
rect 294 1278 298 1282
rect 302 1278 306 1282
rect 310 1258 314 1262
rect 334 1258 338 1262
rect 454 1348 458 1352
rect 430 1338 434 1342
rect 502 1338 506 1342
rect 414 1328 418 1332
rect 574 1388 578 1392
rect 590 1408 594 1412
rect 614 1408 618 1412
rect 534 1358 538 1362
rect 542 1358 546 1362
rect 558 1358 562 1362
rect 526 1338 530 1342
rect 406 1318 410 1322
rect 398 1288 402 1292
rect 374 1278 378 1282
rect 302 1238 306 1242
rect 270 1198 274 1202
rect 326 1138 330 1142
rect 390 1248 394 1252
rect 382 1188 386 1192
rect 374 1138 378 1142
rect 230 1128 234 1132
rect 294 1128 298 1132
rect 302 1128 306 1132
rect 326 1128 330 1132
rect 342 1128 346 1132
rect 254 1118 258 1122
rect 230 1088 234 1092
rect 278 1108 282 1112
rect 222 1058 226 1062
rect 238 1058 242 1062
rect 262 1058 266 1062
rect 214 1048 218 1052
rect 230 1048 234 1052
rect 198 1028 202 1032
rect 190 1008 194 1012
rect 206 1008 210 1012
rect 182 968 186 972
rect 158 958 162 962
rect 158 948 162 952
rect 174 948 178 952
rect 302 1058 306 1062
rect 270 1038 274 1042
rect 374 1118 378 1122
rect 358 1108 362 1112
rect 366 1108 370 1112
rect 350 1098 354 1102
rect 318 1068 322 1072
rect 366 1098 370 1102
rect 526 1318 530 1322
rect 446 1298 450 1302
rect 454 1278 458 1282
rect 502 1278 506 1282
rect 446 1268 450 1272
rect 406 1228 410 1232
rect 406 1208 410 1212
rect 430 1208 434 1212
rect 566 1338 570 1342
rect 558 1318 562 1322
rect 542 1308 546 1312
rect 622 1358 626 1362
rect 654 1358 658 1362
rect 630 1348 634 1352
rect 582 1338 586 1342
rect 630 1338 634 1342
rect 622 1328 626 1332
rect 574 1258 578 1262
rect 486 1228 490 1232
rect 510 1228 514 1232
rect 474 1203 478 1207
rect 481 1203 485 1207
rect 430 1198 434 1202
rect 462 1198 466 1202
rect 422 1178 426 1182
rect 510 1168 514 1172
rect 454 1158 458 1162
rect 446 1148 450 1152
rect 550 1198 554 1202
rect 534 1158 538 1162
rect 566 1178 570 1182
rect 590 1268 594 1272
rect 606 1258 610 1262
rect 774 1398 778 1402
rect 742 1378 746 1382
rect 774 1378 778 1382
rect 678 1348 682 1352
rect 654 1338 658 1342
rect 670 1338 674 1342
rect 638 1328 642 1332
rect 766 1368 770 1372
rect 726 1348 730 1352
rect 694 1328 698 1332
rect 726 1328 730 1332
rect 662 1318 666 1322
rect 702 1318 706 1322
rect 710 1318 714 1322
rect 662 1308 666 1312
rect 694 1288 698 1292
rect 718 1278 722 1282
rect 582 1248 586 1252
rect 670 1248 674 1252
rect 678 1248 682 1252
rect 606 1228 610 1232
rect 598 1218 602 1222
rect 582 1208 586 1212
rect 574 1158 578 1162
rect 590 1148 594 1152
rect 566 1138 570 1142
rect 446 1128 450 1132
rect 486 1128 490 1132
rect 510 1128 514 1132
rect 430 1118 434 1122
rect 518 1118 522 1122
rect 406 1098 410 1102
rect 422 1098 426 1102
rect 374 1068 378 1072
rect 390 1068 394 1072
rect 398 1068 402 1072
rect 406 1058 410 1062
rect 414 1058 418 1062
rect 350 1048 354 1052
rect 374 1048 378 1052
rect 454 1068 458 1072
rect 542 1088 546 1092
rect 614 1168 618 1172
rect 638 1238 642 1242
rect 710 1228 714 1232
rect 718 1188 722 1192
rect 774 1348 778 1352
rect 806 1338 810 1342
rect 782 1318 786 1322
rect 830 1388 834 1392
rect 846 1338 850 1342
rect 838 1328 842 1332
rect 742 1278 746 1282
rect 774 1278 778 1282
rect 734 1268 738 1272
rect 758 1268 762 1272
rect 750 1258 754 1262
rect 742 1238 746 1242
rect 710 1168 714 1172
rect 726 1168 730 1172
rect 654 1158 658 1162
rect 670 1158 674 1162
rect 694 1158 698 1162
rect 654 1148 658 1152
rect 622 1138 626 1142
rect 582 1128 586 1132
rect 614 1128 618 1132
rect 574 1098 578 1102
rect 790 1268 794 1272
rect 814 1268 818 1272
rect 814 1258 818 1262
rect 902 1398 906 1402
rect 902 1358 906 1362
rect 950 1358 954 1362
rect 990 1358 994 1362
rect 1014 1358 1018 1362
rect 886 1348 890 1352
rect 870 1338 874 1342
rect 894 1338 898 1342
rect 886 1298 890 1302
rect 862 1288 866 1292
rect 870 1288 874 1292
rect 886 1288 890 1292
rect 854 1278 858 1282
rect 1038 1348 1042 1352
rect 1054 1348 1058 1352
rect 926 1338 930 1342
rect 958 1338 962 1342
rect 990 1338 994 1342
rect 1022 1338 1026 1342
rect 942 1328 946 1332
rect 1006 1328 1010 1332
rect 1030 1328 1034 1332
rect 1046 1328 1050 1332
rect 1198 1408 1202 1412
rect 1302 1408 1306 1412
rect 1310 1398 1314 1402
rect 1318 1398 1322 1402
rect 1270 1388 1274 1392
rect 1190 1378 1194 1382
rect 1214 1378 1218 1382
rect 1182 1368 1186 1372
rect 1198 1368 1202 1372
rect 1230 1368 1234 1372
rect 1102 1358 1106 1362
rect 1142 1358 1146 1362
rect 1182 1358 1186 1362
rect 1110 1348 1114 1352
rect 1070 1328 1074 1332
rect 1078 1328 1082 1332
rect 1062 1318 1066 1322
rect 902 1308 906 1312
rect 894 1278 898 1282
rect 846 1268 850 1272
rect 870 1268 874 1272
rect 814 1248 818 1252
rect 774 1148 778 1152
rect 862 1258 866 1262
rect 910 1248 914 1252
rect 830 1238 834 1242
rect 822 1228 826 1232
rect 798 1168 802 1172
rect 830 1168 834 1172
rect 846 1168 850 1172
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 966 1278 970 1282
rect 990 1278 994 1282
rect 950 1268 954 1272
rect 942 1258 946 1262
rect 918 1238 922 1242
rect 886 1228 890 1232
rect 942 1228 946 1232
rect 966 1228 970 1232
rect 838 1158 842 1162
rect 862 1158 866 1162
rect 766 1138 770 1142
rect 686 1128 690 1132
rect 790 1128 794 1132
rect 622 1118 626 1122
rect 678 1118 682 1122
rect 670 1108 674 1112
rect 574 1088 578 1092
rect 582 1088 586 1092
rect 630 1088 634 1092
rect 542 1068 546 1072
rect 534 1058 538 1062
rect 550 1058 554 1062
rect 334 1038 338 1042
rect 430 1038 434 1042
rect 494 1038 498 1042
rect 510 1038 514 1042
rect 518 1038 522 1042
rect 678 1088 682 1092
rect 758 1118 762 1122
rect 742 1108 746 1112
rect 766 1108 770 1112
rect 798 1108 802 1112
rect 814 1108 818 1112
rect 822 1108 826 1112
rect 766 1098 770 1102
rect 742 1088 746 1092
rect 798 1088 802 1092
rect 766 1078 770 1082
rect 782 1078 786 1082
rect 606 1068 610 1072
rect 614 1068 618 1072
rect 630 1068 634 1072
rect 678 1068 682 1072
rect 702 1068 706 1072
rect 734 1068 738 1072
rect 598 1058 602 1062
rect 246 1028 250 1032
rect 254 1028 258 1032
rect 286 1028 290 1032
rect 310 1028 314 1032
rect 414 1028 418 1032
rect 358 1008 362 1012
rect 246 998 250 1002
rect 318 998 322 1002
rect 222 978 226 982
rect 238 968 242 972
rect 214 958 218 962
rect 222 958 226 962
rect 198 938 202 942
rect 166 928 170 932
rect 190 928 194 932
rect 310 988 314 992
rect 390 988 394 992
rect 406 988 410 992
rect 390 978 394 982
rect 326 968 330 972
rect 334 958 338 962
rect 246 948 250 952
rect 262 948 266 952
rect 254 938 258 942
rect 286 938 290 942
rect 326 938 330 942
rect 246 908 250 912
rect 190 878 194 882
rect 214 878 218 882
rect 494 1008 498 1012
rect 474 1003 478 1007
rect 481 1003 485 1007
rect 422 958 426 962
rect 446 968 450 972
rect 494 968 498 972
rect 558 968 562 972
rect 534 958 538 962
rect 542 958 546 962
rect 710 1058 714 1062
rect 718 1048 722 1052
rect 854 1148 858 1152
rect 862 1138 866 1142
rect 846 1108 850 1112
rect 862 1088 866 1092
rect 838 1078 842 1082
rect 854 1068 858 1072
rect 902 1168 906 1172
rect 910 1168 914 1172
rect 934 1168 938 1172
rect 958 1168 962 1172
rect 902 1148 906 1152
rect 1078 1308 1082 1312
rect 1070 1278 1074 1282
rect 1086 1278 1090 1282
rect 974 1198 978 1202
rect 982 1178 986 1182
rect 918 1148 922 1152
rect 942 1148 946 1152
rect 950 1148 954 1152
rect 966 1138 970 1142
rect 894 1118 898 1122
rect 918 1118 922 1122
rect 910 1108 914 1112
rect 870 1078 874 1082
rect 878 1068 882 1072
rect 958 1108 962 1112
rect 966 1098 970 1102
rect 942 1068 946 1072
rect 958 1068 962 1072
rect 934 1058 938 1062
rect 846 1048 850 1052
rect 854 1048 858 1052
rect 734 1038 738 1042
rect 742 1038 746 1042
rect 830 1038 834 1042
rect 926 1038 930 1042
rect 830 1028 834 1032
rect 846 1028 850 1032
rect 878 1028 882 1032
rect 886 1028 890 1032
rect 686 1018 690 1022
rect 606 1008 610 1012
rect 654 978 658 982
rect 718 978 722 982
rect 614 968 618 972
rect 646 968 650 972
rect 670 968 674 972
rect 598 958 602 962
rect 614 958 618 962
rect 630 958 634 962
rect 646 958 650 962
rect 686 958 690 962
rect 574 948 578 952
rect 438 938 442 942
rect 470 938 474 942
rect 510 938 514 942
rect 518 938 522 942
rect 550 938 554 942
rect 574 938 578 942
rect 262 928 266 932
rect 334 928 338 932
rect 358 928 362 932
rect 374 928 378 932
rect 270 878 274 882
rect 182 868 186 872
rect 238 868 242 872
rect 206 858 210 862
rect 214 858 218 862
rect 262 858 266 862
rect 158 848 162 852
rect 150 838 154 842
rect 166 838 170 842
rect 286 868 290 872
rect 326 898 330 902
rect 286 858 290 862
rect 302 858 306 862
rect 318 858 322 862
rect 270 848 274 852
rect 294 848 298 852
rect 310 838 314 842
rect 350 888 354 892
rect 438 918 442 922
rect 398 908 402 912
rect 382 898 386 902
rect 358 878 362 882
rect 382 878 386 882
rect 390 858 394 862
rect 414 858 418 862
rect 334 848 338 852
rect 366 848 370 852
rect 390 848 394 852
rect 110 828 114 832
rect 174 828 178 832
rect 222 828 226 832
rect 278 828 282 832
rect 286 828 290 832
rect 166 818 170 822
rect 198 818 202 822
rect 214 818 218 822
rect 230 818 234 822
rect 86 788 90 792
rect 118 768 122 772
rect 214 808 218 812
rect 174 798 178 802
rect 134 748 138 752
rect 94 738 98 742
rect 150 748 154 752
rect 174 738 178 742
rect 166 728 170 732
rect 94 718 98 722
rect 86 708 90 712
rect 142 698 146 702
rect 270 798 274 802
rect 302 788 306 792
rect 286 768 290 772
rect 422 838 426 842
rect 446 878 450 882
rect 526 918 530 922
rect 550 908 554 912
rect 582 918 586 922
rect 534 878 538 882
rect 566 878 570 882
rect 446 848 450 852
rect 462 848 466 852
rect 486 848 490 852
rect 406 828 410 832
rect 454 828 458 832
rect 502 828 506 832
rect 390 758 394 762
rect 222 748 226 752
rect 206 718 210 722
rect 174 708 178 712
rect 474 803 478 807
rect 481 803 485 807
rect 414 748 418 752
rect 430 748 434 752
rect 270 718 274 722
rect 326 718 330 722
rect 350 718 354 722
rect 150 688 154 692
rect 182 688 186 692
rect 214 688 218 692
rect 198 678 202 682
rect 126 668 130 672
rect 158 668 162 672
rect 390 668 394 672
rect 182 658 186 662
rect 214 658 218 662
rect 254 658 258 662
rect 126 648 130 652
rect 318 648 322 652
rect 374 648 378 652
rect 126 638 130 642
rect 158 638 162 642
rect 62 608 66 612
rect 102 608 106 612
rect 38 568 42 572
rect 134 588 138 592
rect 70 548 74 552
rect 38 538 42 542
rect 62 528 66 532
rect 70 528 74 532
rect 30 508 34 512
rect 46 458 50 462
rect 94 508 98 512
rect 118 548 122 552
rect 86 458 90 462
rect 38 448 42 452
rect 78 448 82 452
rect 86 418 90 422
rect 54 408 58 412
rect 54 368 58 372
rect 70 368 74 372
rect 30 358 34 362
rect 14 338 18 342
rect 438 738 442 742
rect 438 728 442 732
rect 454 728 458 732
rect 470 718 474 722
rect 422 658 426 662
rect 638 928 642 932
rect 662 928 666 932
rect 630 918 634 922
rect 614 888 618 892
rect 638 908 642 912
rect 638 898 642 902
rect 598 848 602 852
rect 606 848 610 852
rect 574 828 578 832
rect 534 818 538 822
rect 510 808 514 812
rect 502 788 506 792
rect 622 788 626 792
rect 510 768 514 772
rect 582 768 586 772
rect 638 778 642 782
rect 654 908 658 912
rect 678 888 682 892
rect 702 928 706 932
rect 702 908 706 912
rect 686 848 690 852
rect 790 998 794 1002
rect 734 988 738 992
rect 742 958 746 962
rect 750 938 754 942
rect 766 928 770 932
rect 830 998 834 1002
rect 870 1008 874 1012
rect 862 998 866 1002
rect 854 968 858 972
rect 838 958 842 962
rect 870 948 874 952
rect 894 948 898 952
rect 846 928 850 932
rect 894 928 898 932
rect 806 898 810 902
rect 742 888 746 892
rect 814 888 818 892
rect 774 868 778 872
rect 742 858 746 862
rect 750 858 754 862
rect 766 858 770 862
rect 726 828 730 832
rect 782 828 786 832
rect 798 828 802 832
rect 662 798 666 802
rect 654 788 658 792
rect 630 758 634 762
rect 646 758 650 762
rect 686 808 690 812
rect 694 788 698 792
rect 694 768 698 772
rect 710 768 714 772
rect 726 798 730 802
rect 734 778 738 782
rect 750 768 754 772
rect 686 758 690 762
rect 710 758 714 762
rect 758 748 762 752
rect 766 748 770 752
rect 598 738 602 742
rect 742 738 746 742
rect 790 778 794 782
rect 838 888 842 892
rect 878 888 882 892
rect 910 1008 914 1012
rect 950 998 954 1002
rect 942 988 946 992
rect 918 958 922 962
rect 1086 1258 1090 1262
rect 1070 1248 1074 1252
rect 1086 1238 1090 1242
rect 1102 1208 1106 1212
rect 1166 1348 1170 1352
rect 1126 1338 1130 1342
rect 1150 1338 1154 1342
rect 1206 1358 1210 1362
rect 1238 1358 1242 1362
rect 1222 1348 1226 1352
rect 1166 1328 1170 1332
rect 1118 1318 1122 1322
rect 1142 1318 1146 1322
rect 1206 1318 1210 1322
rect 1118 1268 1122 1272
rect 1142 1268 1146 1272
rect 1134 1258 1138 1262
rect 1142 1248 1146 1252
rect 1046 1188 1050 1192
rect 1110 1188 1114 1192
rect 1070 1178 1074 1182
rect 1134 1178 1138 1182
rect 1006 1168 1010 1172
rect 1022 1168 1026 1172
rect 1030 1158 1034 1162
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 998 1078 1002 1082
rect 1022 1078 1026 1082
rect 990 1048 994 1052
rect 958 958 962 962
rect 974 958 978 962
rect 974 948 978 952
rect 982 948 986 952
rect 1022 1068 1026 1072
rect 1078 1168 1082 1172
rect 1118 1168 1122 1172
rect 1254 1338 1258 1342
rect 1302 1348 1306 1352
rect 1390 1368 1394 1372
rect 1414 1368 1418 1372
rect 1438 1358 1442 1362
rect 1398 1348 1402 1352
rect 1406 1348 1410 1352
rect 1366 1338 1370 1342
rect 1390 1338 1394 1342
rect 1238 1328 1242 1332
rect 1342 1328 1346 1332
rect 1222 1288 1226 1292
rect 1166 1278 1170 1282
rect 1182 1278 1186 1282
rect 1294 1308 1298 1312
rect 1318 1288 1322 1292
rect 1366 1298 1370 1302
rect 1358 1288 1362 1292
rect 1238 1278 1242 1282
rect 1254 1278 1258 1282
rect 1326 1278 1330 1282
rect 1334 1278 1338 1282
rect 1190 1248 1194 1252
rect 1310 1258 1314 1262
rect 1246 1248 1250 1252
rect 1262 1248 1266 1252
rect 1302 1248 1306 1252
rect 1342 1268 1346 1272
rect 1374 1258 1378 1262
rect 1414 1338 1418 1342
rect 1462 1338 1466 1342
rect 1182 1238 1186 1242
rect 1214 1238 1218 1242
rect 1158 1228 1162 1232
rect 1270 1228 1274 1232
rect 1214 1218 1218 1222
rect 1286 1218 1290 1222
rect 1206 1168 1210 1172
rect 1182 1158 1186 1162
rect 1094 1148 1098 1152
rect 1118 1148 1122 1152
rect 1126 1148 1130 1152
rect 1086 1138 1090 1142
rect 1150 1148 1154 1152
rect 1190 1138 1194 1142
rect 1206 1138 1210 1142
rect 1094 1128 1098 1132
rect 1142 1128 1146 1132
rect 1062 1118 1066 1122
rect 1038 1068 1042 1072
rect 1150 1118 1154 1122
rect 1182 1118 1186 1122
rect 1110 1068 1114 1072
rect 1150 1068 1154 1072
rect 1174 1068 1178 1072
rect 1126 1058 1130 1062
rect 1054 1048 1058 1052
rect 1078 1048 1082 1052
rect 1126 1048 1130 1052
rect 1150 1048 1154 1052
rect 1030 1038 1034 1042
rect 1086 1038 1090 1042
rect 1134 1038 1138 1042
rect 1230 1208 1234 1212
rect 1230 1188 1234 1192
rect 1246 1188 1250 1192
rect 1238 1168 1242 1172
rect 1286 1168 1290 1172
rect 1254 1158 1258 1162
rect 1286 1158 1290 1162
rect 1246 1148 1250 1152
rect 1222 1138 1226 1142
rect 1262 1138 1266 1142
rect 1222 1128 1226 1132
rect 1294 1128 1298 1132
rect 1198 1068 1202 1072
rect 1254 1068 1258 1072
rect 1286 1068 1290 1072
rect 1190 1058 1194 1062
rect 1262 1058 1266 1062
rect 1294 1058 1298 1062
rect 1350 1248 1354 1252
rect 1390 1248 1394 1252
rect 1406 1248 1410 1252
rect 1350 1228 1354 1232
rect 1366 1228 1370 1232
rect 1310 1188 1314 1192
rect 1350 1188 1354 1192
rect 1318 1168 1322 1172
rect 1326 1158 1330 1162
rect 1310 1078 1314 1082
rect 1214 1048 1218 1052
rect 1270 1038 1274 1042
rect 1006 1028 1010 1032
rect 1006 1018 1010 1022
rect 1014 1018 1018 1022
rect 1038 1008 1042 1012
rect 1062 998 1066 1002
rect 1014 978 1018 982
rect 1062 978 1066 982
rect 1054 968 1058 972
rect 1078 968 1082 972
rect 1030 948 1034 952
rect 1190 978 1194 982
rect 1254 968 1258 972
rect 1094 958 1098 962
rect 1110 958 1114 962
rect 1134 958 1138 962
rect 1174 958 1178 962
rect 1102 948 1106 952
rect 1126 948 1130 952
rect 1198 948 1202 952
rect 1022 938 1026 942
rect 1054 938 1058 942
rect 1086 938 1090 942
rect 1142 938 1146 942
rect 1150 938 1154 942
rect 1190 938 1194 942
rect 910 928 914 932
rect 998 928 1002 932
rect 1014 928 1018 932
rect 1078 908 1082 912
rect 986 903 990 907
rect 993 903 997 907
rect 902 878 906 882
rect 830 858 834 862
rect 838 858 842 862
rect 862 828 866 832
rect 822 768 826 772
rect 838 768 842 772
rect 782 738 786 742
rect 798 738 802 742
rect 814 738 818 742
rect 846 738 850 742
rect 870 738 874 742
rect 878 738 882 742
rect 598 728 602 732
rect 790 728 794 732
rect 814 728 818 732
rect 846 728 850 732
rect 878 728 882 732
rect 902 838 906 842
rect 934 888 938 892
rect 966 888 970 892
rect 1182 918 1186 922
rect 1174 898 1178 902
rect 1150 888 1154 892
rect 1166 888 1170 892
rect 998 878 1002 882
rect 1014 878 1018 882
rect 1062 878 1066 882
rect 958 868 962 872
rect 1030 868 1034 872
rect 1046 868 1050 872
rect 1062 868 1066 872
rect 1046 858 1050 862
rect 934 848 938 852
rect 950 848 954 852
rect 974 848 978 852
rect 1006 848 1010 852
rect 1014 768 1018 772
rect 1014 748 1018 752
rect 942 738 946 742
rect 910 728 914 732
rect 566 718 570 722
rect 558 708 562 712
rect 542 698 546 702
rect 806 718 810 722
rect 870 718 874 722
rect 614 688 618 692
rect 622 688 626 692
rect 830 698 834 702
rect 870 698 874 702
rect 662 688 666 692
rect 846 688 850 692
rect 638 678 642 682
rect 646 678 650 682
rect 726 678 730 682
rect 590 668 594 672
rect 630 668 634 672
rect 598 658 602 662
rect 510 648 514 652
rect 438 638 442 642
rect 478 638 482 642
rect 454 618 458 622
rect 190 568 194 572
rect 126 478 130 482
rect 110 458 114 462
rect 102 448 106 452
rect 54 358 58 362
rect 46 318 50 322
rect 94 348 98 352
rect 70 338 74 342
rect 174 508 178 512
rect 166 458 170 462
rect 110 388 114 392
rect 134 388 138 392
rect 126 368 130 372
rect 102 338 106 342
rect 86 328 90 332
rect 126 338 130 342
rect 118 318 122 322
rect 110 308 114 312
rect 62 278 66 282
rect 94 278 98 282
rect 46 268 50 272
rect 278 558 282 562
rect 318 558 322 562
rect 334 558 338 562
rect 326 548 330 552
rect 342 548 346 552
rect 350 548 354 552
rect 310 538 314 542
rect 422 578 426 582
rect 474 603 478 607
rect 481 603 485 607
rect 526 588 530 592
rect 454 568 458 572
rect 518 568 522 572
rect 366 548 370 552
rect 382 548 386 552
rect 206 528 210 532
rect 246 528 250 532
rect 294 528 298 532
rect 358 528 362 532
rect 406 528 410 532
rect 254 518 258 522
rect 198 508 202 512
rect 238 508 242 512
rect 494 558 498 562
rect 454 528 458 532
rect 430 508 434 512
rect 422 498 426 502
rect 294 478 298 482
rect 446 478 450 482
rect 190 468 194 472
rect 262 468 266 472
rect 198 458 202 462
rect 214 458 218 462
rect 246 458 250 462
rect 278 458 282 462
rect 174 438 178 442
rect 182 438 186 442
rect 166 408 170 412
rect 166 388 170 392
rect 158 368 162 372
rect 190 368 194 372
rect 134 278 138 282
rect 110 268 114 272
rect 126 268 130 272
rect 6 258 10 262
rect 38 258 42 262
rect 94 258 98 262
rect 38 248 42 252
rect 86 238 90 242
rect 22 218 26 222
rect 46 168 50 172
rect 70 168 74 172
rect 14 138 18 142
rect 78 148 82 152
rect 62 138 66 142
rect 38 128 42 132
rect 46 128 50 132
rect 54 128 58 132
rect 302 468 306 472
rect 318 468 322 472
rect 334 468 338 472
rect 382 468 386 472
rect 390 458 394 462
rect 438 458 442 462
rect 222 448 226 452
rect 286 448 290 452
rect 350 448 354 452
rect 382 448 386 452
rect 238 438 242 442
rect 318 438 322 442
rect 246 388 250 392
rect 294 388 298 392
rect 238 368 242 372
rect 302 378 306 382
rect 326 378 330 382
rect 222 358 226 362
rect 238 358 242 362
rect 182 348 186 352
rect 166 328 170 332
rect 214 328 218 332
rect 206 308 210 312
rect 198 268 202 272
rect 222 268 226 272
rect 158 258 162 262
rect 190 258 194 262
rect 158 248 162 252
rect 166 238 170 242
rect 126 228 130 232
rect 134 218 138 222
rect 158 168 162 172
rect 102 158 106 162
rect 110 158 114 162
rect 78 78 82 82
rect 102 78 106 82
rect 126 138 130 142
rect 118 128 122 132
rect 158 148 162 152
rect 286 348 290 352
rect 358 438 362 442
rect 414 438 418 442
rect 430 438 434 442
rect 382 418 386 422
rect 414 378 418 382
rect 358 368 362 372
rect 366 368 370 372
rect 398 358 402 362
rect 390 348 394 352
rect 406 348 410 352
rect 454 428 458 432
rect 478 448 482 452
rect 462 418 466 422
rect 474 403 478 407
rect 481 403 485 407
rect 518 548 522 552
rect 550 568 554 572
rect 542 498 546 502
rect 550 498 554 502
rect 534 488 538 492
rect 534 468 538 472
rect 510 368 514 372
rect 494 358 498 362
rect 366 338 370 342
rect 422 338 426 342
rect 462 338 466 342
rect 254 328 258 332
rect 302 328 306 332
rect 310 328 314 332
rect 350 328 354 332
rect 374 328 378 332
rect 286 318 290 322
rect 326 318 330 322
rect 310 288 314 292
rect 278 268 282 272
rect 262 258 266 262
rect 302 258 306 262
rect 430 318 434 322
rect 470 298 474 302
rect 382 278 386 282
rect 406 278 410 282
rect 414 278 418 282
rect 334 268 338 272
rect 534 438 538 442
rect 534 428 538 432
rect 526 378 530 382
rect 566 518 570 522
rect 566 478 570 482
rect 558 448 562 452
rect 550 438 554 442
rect 598 638 602 642
rect 582 558 586 562
rect 590 528 594 532
rect 582 518 586 522
rect 582 508 586 512
rect 614 568 618 572
rect 622 548 626 552
rect 614 528 618 532
rect 606 458 610 462
rect 622 458 626 462
rect 614 398 618 402
rect 582 378 586 382
rect 542 368 546 372
rect 566 368 570 372
rect 598 368 602 372
rect 678 668 682 672
rect 654 648 658 652
rect 686 648 690 652
rect 678 638 682 642
rect 702 638 706 642
rect 638 588 642 592
rect 646 588 650 592
rect 662 578 666 582
rect 638 568 642 572
rect 782 668 786 672
rect 806 668 810 672
rect 766 648 770 652
rect 742 638 746 642
rect 758 628 762 632
rect 726 618 730 622
rect 734 588 738 592
rect 750 578 754 582
rect 686 568 690 572
rect 718 568 722 572
rect 822 658 826 662
rect 814 638 818 642
rect 838 638 842 642
rect 814 628 818 632
rect 830 628 834 632
rect 790 618 794 622
rect 774 578 778 582
rect 798 578 802 582
rect 806 578 810 582
rect 766 568 770 572
rect 830 598 834 602
rect 838 568 842 572
rect 718 558 722 562
rect 742 558 746 562
rect 774 558 778 562
rect 734 548 738 552
rect 694 538 698 542
rect 758 538 762 542
rect 790 538 794 542
rect 806 538 810 542
rect 646 528 650 532
rect 758 528 762 532
rect 654 518 658 522
rect 734 518 738 522
rect 742 508 746 512
rect 734 498 738 502
rect 678 488 682 492
rect 646 478 650 482
rect 694 478 698 482
rect 638 468 642 472
rect 662 468 666 472
rect 750 468 754 472
rect 670 458 674 462
rect 662 448 666 452
rect 686 448 690 452
rect 630 428 634 432
rect 670 398 674 402
rect 638 378 642 382
rect 790 508 794 512
rect 806 478 810 482
rect 774 468 778 472
rect 758 458 762 462
rect 790 458 794 462
rect 750 448 754 452
rect 782 448 786 452
rect 702 438 706 442
rect 742 438 746 442
rect 790 418 794 422
rect 782 398 786 402
rect 622 358 626 362
rect 510 348 514 352
rect 518 348 522 352
rect 550 348 554 352
rect 574 338 578 342
rect 606 338 610 342
rect 558 298 562 302
rect 558 288 562 292
rect 542 278 546 282
rect 582 278 586 282
rect 606 278 610 282
rect 518 268 522 272
rect 566 268 570 272
rect 326 258 330 262
rect 350 258 354 262
rect 374 258 378 262
rect 446 258 450 262
rect 470 258 474 262
rect 542 258 546 262
rect 342 248 346 252
rect 198 218 202 222
rect 254 238 258 242
rect 270 238 274 242
rect 318 238 322 242
rect 238 168 242 172
rect 190 158 194 162
rect 166 138 170 142
rect 174 138 178 142
rect 166 88 170 92
rect 126 78 130 82
rect 134 78 138 82
rect 46 68 50 72
rect 94 68 98 72
rect 6 58 10 62
rect 134 48 138 52
rect 62 8 66 12
rect 86 8 90 12
rect 190 118 194 122
rect 198 98 202 102
rect 270 218 274 222
rect 262 168 266 172
rect 286 168 290 172
rect 294 168 298 172
rect 270 158 274 162
rect 326 158 330 162
rect 254 148 258 152
rect 294 148 298 152
rect 326 148 330 152
rect 230 138 234 142
rect 238 138 242 142
rect 214 108 218 112
rect 182 78 186 82
rect 198 78 202 82
rect 174 68 178 72
rect 222 98 226 102
rect 374 248 378 252
rect 398 248 402 252
rect 438 238 442 242
rect 446 238 450 242
rect 382 228 386 232
rect 358 218 362 222
rect 390 198 394 202
rect 374 158 378 162
rect 486 248 490 252
rect 534 238 538 242
rect 474 203 478 207
rect 481 203 485 207
rect 590 268 594 272
rect 630 348 634 352
rect 630 338 634 342
rect 638 338 642 342
rect 686 368 690 372
rect 742 368 746 372
rect 662 348 666 352
rect 646 328 650 332
rect 630 268 634 272
rect 622 258 626 262
rect 598 218 602 222
rect 566 198 570 202
rect 590 198 594 202
rect 542 188 546 192
rect 454 178 458 182
rect 518 178 522 182
rect 398 158 402 162
rect 294 128 298 132
rect 350 128 354 132
rect 382 128 386 132
rect 414 128 418 132
rect 270 78 274 82
rect 342 78 346 82
rect 350 78 354 82
rect 230 68 234 72
rect 262 68 266 72
rect 270 68 274 72
rect 246 38 250 42
rect 286 38 290 42
rect 326 68 330 72
rect 382 108 386 112
rect 438 158 442 162
rect 438 118 442 122
rect 446 118 450 122
rect 438 108 442 112
rect 470 88 474 92
rect 446 78 450 82
rect 366 68 370 72
rect 334 48 338 52
rect 374 48 378 52
rect 318 28 322 32
rect 398 58 402 62
rect 390 18 394 22
rect 374 8 378 12
rect 486 138 490 142
rect 502 78 506 82
rect 542 158 546 162
rect 542 138 546 142
rect 534 118 538 122
rect 542 88 546 92
rect 518 58 522 62
rect 534 58 538 62
rect 478 48 482 52
rect 494 48 498 52
rect 502 48 506 52
rect 510 48 514 52
rect 474 3 478 7
rect 481 3 485 7
rect 558 118 562 122
rect 574 118 578 122
rect 622 238 626 242
rect 638 188 642 192
rect 606 168 610 172
rect 614 168 618 172
rect 678 288 682 292
rect 654 268 658 272
rect 718 318 722 322
rect 782 358 786 362
rect 750 348 754 352
rect 774 348 778 352
rect 774 328 778 332
rect 758 308 762 312
rect 718 278 722 282
rect 750 278 754 282
rect 830 508 834 512
rect 830 488 834 492
rect 886 648 890 652
rect 870 638 874 642
rect 910 718 914 722
rect 1062 838 1066 842
rect 1214 958 1218 962
rect 1238 948 1242 952
rect 1222 938 1226 942
rect 1230 888 1234 892
rect 1222 878 1226 882
rect 1254 948 1258 952
rect 1254 928 1258 932
rect 1262 898 1266 902
rect 1318 1048 1322 1052
rect 1310 1038 1314 1042
rect 1302 998 1306 1002
rect 1294 968 1298 972
rect 1358 1178 1362 1182
rect 1398 1238 1402 1242
rect 1390 1218 1394 1222
rect 1382 1188 1386 1192
rect 1366 1158 1370 1162
rect 1358 1148 1362 1152
rect 1382 1148 1386 1152
rect 1334 1138 1338 1142
rect 1438 1278 1442 1282
rect 1422 1258 1426 1262
rect 1446 1258 1450 1262
rect 1430 1168 1434 1172
rect 1438 1148 1442 1152
rect 1422 1138 1426 1142
rect 1374 1118 1378 1122
rect 1342 1088 1346 1092
rect 1366 1068 1370 1072
rect 1390 1068 1394 1072
rect 1350 1058 1354 1062
rect 1342 1038 1346 1042
rect 1358 1038 1362 1042
rect 1382 1018 1386 1022
rect 1334 1008 1338 1012
rect 1454 1208 1458 1212
rect 1454 1148 1458 1152
rect 1446 1108 1450 1112
rect 1414 1088 1418 1092
rect 1406 1048 1410 1052
rect 1398 998 1402 1002
rect 1398 988 1402 992
rect 1358 978 1362 982
rect 1366 978 1370 982
rect 1350 968 1354 972
rect 1350 958 1354 962
rect 1286 948 1290 952
rect 1278 908 1282 912
rect 1286 908 1290 912
rect 1262 878 1266 882
rect 1294 878 1298 882
rect 1110 868 1114 872
rect 1158 868 1162 872
rect 1190 868 1194 872
rect 1230 868 1234 872
rect 1254 868 1258 872
rect 1086 858 1090 862
rect 1118 858 1122 862
rect 1094 848 1098 852
rect 1166 848 1170 852
rect 1254 838 1258 842
rect 1278 828 1282 832
rect 1254 798 1258 802
rect 1118 778 1122 782
rect 1078 768 1082 772
rect 1398 968 1402 972
rect 1326 948 1330 952
rect 1350 938 1354 942
rect 1318 908 1322 912
rect 1318 858 1322 862
rect 1326 818 1330 822
rect 1310 788 1314 792
rect 1126 758 1130 762
rect 1294 758 1298 762
rect 1302 758 1306 762
rect 1046 748 1050 752
rect 1078 748 1082 752
rect 1094 748 1098 752
rect 1182 748 1186 752
rect 1262 748 1266 752
rect 1278 748 1282 752
rect 1310 748 1314 752
rect 1438 1088 1442 1092
rect 1430 1078 1434 1082
rect 1446 1068 1450 1072
rect 1422 1038 1426 1042
rect 1446 1028 1450 1032
rect 1430 1008 1434 1012
rect 1446 978 1450 982
rect 1438 968 1442 972
rect 1422 958 1426 962
rect 1398 938 1402 942
rect 1414 938 1418 942
rect 1446 948 1450 952
rect 1470 948 1474 952
rect 1438 898 1442 902
rect 1422 888 1426 892
rect 1366 868 1370 872
rect 1414 868 1418 872
rect 1438 868 1442 872
rect 1350 858 1354 862
rect 1398 858 1402 862
rect 1438 858 1442 862
rect 1358 848 1362 852
rect 1438 788 1442 792
rect 1350 758 1354 762
rect 1062 738 1066 742
rect 1086 738 1090 742
rect 1134 738 1138 742
rect 1286 738 1290 742
rect 1318 738 1322 742
rect 1334 738 1338 742
rect 1462 838 1466 842
rect 1454 808 1458 812
rect 1478 868 1482 872
rect 1478 848 1482 852
rect 1454 738 1458 742
rect 942 728 946 732
rect 1030 728 1034 732
rect 1070 728 1074 732
rect 1102 728 1106 732
rect 1254 728 1258 732
rect 1286 728 1290 732
rect 926 708 930 712
rect 1166 718 1170 722
rect 986 703 990 707
rect 993 703 997 707
rect 1022 678 1026 682
rect 1118 678 1122 682
rect 1254 698 1258 702
rect 1222 678 1226 682
rect 926 668 930 672
rect 1038 668 1042 672
rect 1198 668 1202 672
rect 1246 668 1250 672
rect 934 658 938 662
rect 966 658 970 662
rect 1102 658 1106 662
rect 1142 659 1146 663
rect 902 648 906 652
rect 894 608 898 612
rect 926 648 930 652
rect 942 648 946 652
rect 974 648 978 652
rect 1070 648 1074 652
rect 958 638 962 642
rect 990 638 994 642
rect 1022 638 1026 642
rect 974 628 978 632
rect 862 588 866 592
rect 1006 588 1010 592
rect 910 578 914 582
rect 942 578 946 582
rect 886 568 890 572
rect 854 548 858 552
rect 862 538 866 542
rect 886 548 890 552
rect 870 498 874 502
rect 894 488 898 492
rect 862 468 866 472
rect 886 468 890 472
rect 838 448 842 452
rect 814 378 818 382
rect 870 458 874 462
rect 910 538 914 542
rect 934 558 938 562
rect 950 548 954 552
rect 966 548 970 552
rect 942 538 946 542
rect 974 538 978 542
rect 1022 578 1026 582
rect 1062 578 1066 582
rect 1014 568 1018 572
rect 1054 568 1058 572
rect 1038 558 1042 562
rect 1062 548 1066 552
rect 1030 538 1034 542
rect 958 508 962 512
rect 942 498 946 502
rect 986 503 990 507
rect 993 503 997 507
rect 934 488 938 492
rect 1006 488 1010 492
rect 982 478 986 482
rect 910 468 914 472
rect 918 468 922 472
rect 1038 488 1042 492
rect 1046 488 1050 492
rect 934 458 938 462
rect 974 458 978 462
rect 942 448 946 452
rect 870 438 874 442
rect 870 428 874 432
rect 934 438 938 442
rect 902 408 906 412
rect 846 368 850 372
rect 902 368 906 372
rect 806 348 810 352
rect 814 338 818 342
rect 838 338 842 342
rect 846 338 850 342
rect 918 428 922 432
rect 958 408 962 412
rect 950 398 954 402
rect 926 368 930 372
rect 878 358 882 362
rect 870 338 874 342
rect 814 328 818 332
rect 830 328 834 332
rect 846 328 850 332
rect 862 328 866 332
rect 822 318 826 322
rect 806 308 810 312
rect 790 278 794 282
rect 726 268 730 272
rect 782 268 786 272
rect 814 268 818 272
rect 830 268 834 272
rect 694 258 698 262
rect 710 258 714 262
rect 726 258 730 262
rect 774 258 778 262
rect 670 208 674 212
rect 678 198 682 202
rect 726 228 730 232
rect 694 188 698 192
rect 750 208 754 212
rect 734 178 738 182
rect 798 248 802 252
rect 870 268 874 272
rect 862 238 866 242
rect 902 338 906 342
rect 894 318 898 322
rect 894 298 898 302
rect 934 348 938 352
rect 966 368 970 372
rect 1038 418 1042 422
rect 1062 408 1066 412
rect 1134 608 1138 612
rect 1078 558 1082 562
rect 1350 718 1354 722
rect 1310 678 1314 682
rect 1262 668 1266 672
rect 1278 668 1282 672
rect 1302 668 1306 672
rect 1350 668 1354 672
rect 1478 668 1482 672
rect 1414 658 1418 662
rect 1206 648 1210 652
rect 1246 648 1250 652
rect 1286 628 1290 632
rect 1414 648 1418 652
rect 1446 648 1450 652
rect 1366 618 1370 622
rect 1286 608 1290 612
rect 1318 608 1322 612
rect 1254 588 1258 592
rect 1294 588 1298 592
rect 1222 578 1226 582
rect 1278 578 1282 582
rect 1190 568 1194 572
rect 1262 568 1266 572
rect 1270 568 1274 572
rect 1158 538 1162 542
rect 1094 528 1098 532
rect 1094 488 1098 492
rect 1174 508 1178 512
rect 1198 548 1202 552
rect 1222 558 1226 562
rect 1246 558 1250 562
rect 1238 538 1242 542
rect 1214 528 1218 532
rect 1238 528 1242 532
rect 1438 628 1442 632
rect 1446 548 1450 552
rect 1478 548 1482 552
rect 1286 538 1290 542
rect 1334 528 1338 532
rect 1286 498 1290 502
rect 1302 498 1306 502
rect 1078 478 1082 482
rect 1102 478 1106 482
rect 1134 478 1138 482
rect 1206 478 1210 482
rect 1230 478 1234 482
rect 1094 468 1098 472
rect 1126 468 1130 472
rect 1302 468 1306 472
rect 1110 458 1114 462
rect 1150 458 1154 462
rect 1262 458 1266 462
rect 1222 448 1226 452
rect 1078 438 1082 442
rect 1086 438 1090 442
rect 1086 368 1090 372
rect 974 358 978 362
rect 1142 358 1146 362
rect 950 338 954 342
rect 998 338 1002 342
rect 1014 328 1018 332
rect 910 288 914 292
rect 918 278 922 282
rect 934 278 938 282
rect 942 278 946 282
rect 910 268 914 272
rect 926 268 930 272
rect 918 258 922 262
rect 894 208 898 212
rect 798 198 802 202
rect 878 198 882 202
rect 950 258 954 262
rect 926 198 930 202
rect 934 198 938 202
rect 718 168 722 172
rect 742 168 746 172
rect 774 168 778 172
rect 822 178 826 182
rect 910 178 914 182
rect 654 158 658 162
rect 678 158 682 162
rect 710 158 714 162
rect 734 158 738 162
rect 798 158 802 162
rect 646 148 650 152
rect 630 118 634 122
rect 606 88 610 92
rect 622 78 626 82
rect 630 58 634 62
rect 622 48 626 52
rect 574 18 578 22
rect 582 18 586 22
rect 598 18 602 22
rect 598 8 602 12
rect 638 38 642 42
rect 638 18 642 22
rect 670 118 674 122
rect 694 118 698 122
rect 878 168 882 172
rect 846 158 850 162
rect 758 148 762 152
rect 814 148 818 152
rect 742 128 746 132
rect 662 78 666 82
rect 662 68 666 72
rect 678 68 682 72
rect 702 58 706 62
rect 798 128 802 132
rect 766 118 770 122
rect 782 118 786 122
rect 750 88 754 92
rect 838 118 842 122
rect 894 128 898 132
rect 870 118 874 122
rect 862 98 866 102
rect 918 138 922 142
rect 958 248 962 252
rect 986 303 990 307
rect 993 303 997 307
rect 1006 298 1010 302
rect 982 268 986 272
rect 1062 348 1066 352
rect 1102 348 1106 352
rect 1030 338 1034 342
rect 1030 328 1034 332
rect 1094 338 1098 342
rect 1118 338 1122 342
rect 1110 328 1114 332
rect 1142 328 1146 332
rect 1070 288 1074 292
rect 1030 278 1034 282
rect 1038 258 1042 262
rect 982 248 986 252
rect 1014 238 1018 242
rect 958 208 962 212
rect 966 178 970 182
rect 982 168 986 172
rect 998 168 1002 172
rect 934 158 938 162
rect 958 158 962 162
rect 950 128 954 132
rect 966 108 970 112
rect 986 103 990 107
rect 993 103 997 107
rect 846 78 850 82
rect 926 78 930 82
rect 942 78 946 82
rect 998 78 1002 82
rect 758 68 762 72
rect 766 68 770 72
rect 774 68 778 72
rect 814 68 818 72
rect 830 68 834 72
rect 862 68 866 72
rect 894 68 898 72
rect 886 58 890 62
rect 910 58 914 62
rect 934 58 938 62
rect 710 28 714 32
rect 742 18 746 22
rect 886 38 890 42
rect 646 8 650 12
rect 662 8 666 12
rect 814 8 818 12
rect 910 8 914 12
rect 966 68 970 72
rect 1126 278 1130 282
rect 1102 258 1106 262
rect 1054 248 1058 252
rect 1078 248 1082 252
rect 1086 248 1090 252
rect 1102 248 1106 252
rect 1046 208 1050 212
rect 1038 198 1042 202
rect 1046 188 1050 192
rect 1046 178 1050 182
rect 1238 428 1242 432
rect 1206 378 1210 382
rect 1246 368 1250 372
rect 1270 448 1274 452
rect 1294 448 1298 452
rect 1334 508 1338 512
rect 1430 508 1434 512
rect 1382 498 1386 502
rect 1462 488 1466 492
rect 1334 478 1338 482
rect 1342 478 1346 482
rect 1382 478 1386 482
rect 1470 468 1474 472
rect 1334 458 1338 462
rect 1358 448 1362 452
rect 1302 438 1306 442
rect 1318 438 1322 442
rect 1278 428 1282 432
rect 1350 428 1354 432
rect 1334 418 1338 422
rect 1374 418 1378 422
rect 1310 398 1314 402
rect 1390 458 1394 462
rect 1430 458 1434 462
rect 1446 448 1450 452
rect 1422 438 1426 442
rect 1382 378 1386 382
rect 1358 368 1362 372
rect 1406 388 1410 392
rect 1398 368 1402 372
rect 1174 358 1178 362
rect 1190 358 1194 362
rect 1230 358 1234 362
rect 1270 358 1274 362
rect 1302 358 1306 362
rect 1318 358 1322 362
rect 1334 358 1338 362
rect 1366 358 1370 362
rect 1374 358 1378 362
rect 1190 348 1194 352
rect 1198 338 1202 342
rect 1190 328 1194 332
rect 1166 308 1170 312
rect 1238 348 1242 352
rect 1246 328 1250 332
rect 1222 318 1226 322
rect 1214 308 1218 312
rect 1206 298 1210 302
rect 1166 258 1170 262
rect 1190 258 1194 262
rect 1206 258 1210 262
rect 1174 228 1178 232
rect 1158 218 1162 222
rect 1182 218 1186 222
rect 1150 208 1154 212
rect 1182 198 1186 202
rect 1110 178 1114 182
rect 1126 178 1130 182
rect 1030 168 1034 172
rect 1062 168 1066 172
rect 1070 168 1074 172
rect 1126 168 1130 172
rect 1166 168 1170 172
rect 1102 158 1106 162
rect 1134 158 1138 162
rect 1158 158 1162 162
rect 1022 148 1026 152
rect 1062 148 1066 152
rect 1022 118 1026 122
rect 1030 118 1034 122
rect 1030 108 1034 112
rect 1038 78 1042 82
rect 1150 148 1154 152
rect 1086 128 1090 132
rect 1158 128 1162 132
rect 1094 118 1098 122
rect 1118 118 1122 122
rect 1094 108 1098 112
rect 1086 98 1090 102
rect 1238 298 1242 302
rect 1222 288 1226 292
rect 1230 278 1234 282
rect 1230 248 1234 252
rect 1198 178 1202 182
rect 1182 148 1186 152
rect 1166 118 1170 122
rect 1190 138 1194 142
rect 1190 108 1194 112
rect 1174 88 1178 92
rect 1134 78 1138 82
rect 1078 68 1082 72
rect 1094 68 1098 72
rect 1118 68 1122 72
rect 1030 58 1034 62
rect 1054 58 1058 62
rect 1086 58 1090 62
rect 1110 58 1114 62
rect 1022 28 1026 32
rect 1158 68 1162 72
rect 1206 148 1210 152
rect 1246 228 1250 232
rect 1270 348 1274 352
rect 1286 348 1290 352
rect 1262 318 1266 322
rect 1262 258 1266 262
rect 1278 338 1282 342
rect 1310 338 1314 342
rect 1302 328 1306 332
rect 1278 268 1282 272
rect 1294 268 1298 272
rect 1302 258 1306 262
rect 1326 348 1330 352
rect 1374 348 1378 352
rect 1390 338 1394 342
rect 1358 328 1362 332
rect 1342 308 1346 312
rect 1382 318 1386 322
rect 1358 278 1362 282
rect 1414 378 1418 382
rect 1430 398 1434 402
rect 1406 338 1410 342
rect 1422 368 1426 372
rect 1414 318 1418 322
rect 1422 318 1426 322
rect 1454 348 1458 352
rect 1470 318 1474 322
rect 1462 288 1466 292
rect 1398 238 1402 242
rect 1358 228 1362 232
rect 1310 218 1314 222
rect 1254 188 1258 192
rect 1286 188 1290 192
rect 1358 188 1362 192
rect 1238 148 1242 152
rect 1222 128 1226 132
rect 1222 98 1226 102
rect 1238 98 1242 102
rect 1182 68 1186 72
rect 1190 58 1194 62
rect 1206 58 1210 62
rect 1214 58 1218 62
rect 1174 28 1178 32
rect 1150 8 1154 12
rect 1246 58 1250 62
rect 1374 178 1378 182
rect 1390 168 1394 172
rect 1430 228 1434 232
rect 1430 218 1434 222
rect 1278 158 1282 162
rect 1302 158 1306 162
rect 1350 158 1354 162
rect 1382 158 1386 162
rect 1310 148 1314 152
rect 1358 148 1362 152
rect 1270 118 1274 122
rect 1318 108 1322 112
rect 1350 118 1354 122
rect 1366 108 1370 112
rect 1334 88 1338 92
rect 1358 78 1362 82
rect 1262 68 1266 72
rect 1302 58 1306 62
rect 1334 58 1338 62
rect 1270 48 1274 52
rect 1310 48 1314 52
rect 1326 48 1330 52
rect 1254 18 1258 22
rect 1318 38 1322 42
rect 1398 148 1402 152
rect 1406 138 1410 142
rect 1390 128 1394 132
rect 1430 178 1434 182
rect 1422 158 1426 162
rect 1422 128 1426 132
rect 1414 118 1418 122
rect 1430 118 1434 122
rect 1446 108 1450 112
rect 1462 78 1466 82
rect 1382 58 1386 62
rect 1358 48 1362 52
rect 1414 48 1418 52
<< metal3 >>
rect 434 1408 438 1411
rect 594 1408 614 1411
rect 1194 1408 1198 1411
rect 1306 1408 1310 1411
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 486 1403 488 1407
rect 498 1398 774 1401
rect 906 1398 1310 1401
rect 1314 1398 1318 1401
rect 170 1388 518 1391
rect 834 1388 1270 1391
rect 358 1378 494 1381
rect 574 1381 577 1388
rect 574 1378 742 1381
rect 778 1378 1190 1381
rect 1194 1378 1214 1381
rect 358 1372 361 1378
rect 298 1368 358 1371
rect 402 1368 454 1371
rect 458 1368 502 1371
rect 522 1368 766 1371
rect 770 1368 1182 1371
rect 1186 1368 1198 1371
rect 1394 1368 1414 1371
rect 90 1358 142 1361
rect 210 1358 238 1361
rect 250 1358 390 1361
rect 410 1358 534 1361
rect 538 1358 542 1361
rect 546 1358 550 1361
rect 562 1358 590 1361
rect 626 1358 630 1361
rect 650 1358 654 1361
rect 738 1358 902 1361
rect 938 1358 950 1361
rect 994 1358 1014 1361
rect 1094 1358 1102 1361
rect 1106 1358 1142 1361
rect 1186 1358 1206 1361
rect 1230 1361 1233 1368
rect 1230 1358 1238 1361
rect 1398 1358 1438 1361
rect 1398 1352 1401 1358
rect -26 1351 -22 1352
rect -26 1348 54 1351
rect 58 1348 270 1351
rect 338 1348 342 1351
rect 458 1348 614 1351
rect 634 1348 678 1351
rect 730 1348 774 1351
rect 890 1348 894 1351
rect 1042 1348 1054 1351
rect 1058 1348 1110 1351
rect 1170 1348 1222 1351
rect 1502 1351 1506 1352
rect 1410 1348 1506 1351
rect 42 1338 86 1341
rect 90 1338 182 1341
rect 202 1338 222 1341
rect 226 1338 254 1341
rect 338 1338 358 1341
rect 362 1338 366 1341
rect 434 1338 502 1341
rect 506 1338 526 1341
rect 530 1338 566 1341
rect 570 1338 582 1341
rect 586 1338 630 1341
rect 658 1338 670 1341
rect 810 1338 846 1341
rect 850 1338 870 1341
rect 874 1338 894 1341
rect 898 1338 926 1341
rect 962 1338 990 1341
rect 1026 1338 1126 1341
rect 1154 1338 1254 1341
rect 1258 1338 1262 1341
rect 1302 1341 1305 1348
rect 1302 1338 1366 1341
rect 1370 1338 1382 1341
rect 1386 1338 1390 1341
rect 1418 1338 1462 1341
rect -26 1331 -22 1332
rect -26 1328 6 1331
rect 154 1328 286 1331
rect 290 1328 302 1331
rect 318 1328 326 1331
rect 330 1328 414 1331
rect 626 1328 638 1331
rect 698 1328 726 1331
rect 778 1328 838 1331
rect 850 1328 942 1331
rect 1010 1328 1030 1331
rect 1034 1328 1046 1331
rect 1050 1328 1070 1331
rect 1118 1328 1166 1331
rect 1206 1328 1238 1331
rect 1322 1328 1342 1331
rect 1502 1331 1506 1332
rect 1346 1328 1506 1331
rect 1078 1322 1081 1328
rect 1118 1322 1121 1328
rect 1206 1322 1209 1328
rect 242 1318 406 1321
rect 530 1318 558 1321
rect 562 1318 646 1321
rect 666 1318 694 1321
rect 698 1318 702 1321
rect 714 1318 782 1321
rect 922 1318 1062 1321
rect 1134 1318 1142 1321
rect 1146 1318 1198 1321
rect 10 1308 542 1311
rect 546 1308 662 1311
rect 666 1308 902 1311
rect 1082 1308 1222 1311
rect 1298 1308 1358 1311
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 138 1298 382 1301
rect 450 1298 886 1301
rect 1150 1298 1366 1301
rect 294 1288 334 1291
rect 354 1288 398 1291
rect 402 1288 518 1291
rect 626 1288 694 1291
rect 730 1288 862 1291
rect 866 1288 870 1291
rect 1150 1291 1153 1298
rect 890 1288 1153 1291
rect 1226 1288 1318 1291
rect 1322 1288 1358 1291
rect 294 1282 297 1288
rect 274 1278 294 1281
rect 342 1281 345 1288
rect 306 1278 345 1281
rect 378 1278 454 1281
rect 458 1278 502 1281
rect 722 1278 742 1281
rect 746 1278 774 1281
rect 850 1278 854 1281
rect 898 1278 966 1281
rect 994 1278 998 1281
rect 1074 1278 1086 1281
rect 1118 1278 1166 1281
rect 1186 1278 1190 1281
rect 1202 1278 1238 1281
rect 1258 1278 1326 1281
rect 1338 1278 1438 1281
rect 1118 1272 1121 1278
rect -26 1271 -22 1272
rect -26 1268 38 1271
rect 74 1268 102 1271
rect 274 1268 446 1271
rect 762 1268 790 1271
rect 818 1268 846 1271
rect 1146 1268 1342 1271
rect 54 1261 57 1268
rect 54 1258 70 1261
rect 90 1258 110 1261
rect 158 1261 161 1268
rect 154 1258 161 1261
rect 202 1258 206 1261
rect 218 1258 310 1261
rect 338 1258 574 1261
rect 590 1261 593 1268
rect 590 1258 606 1261
rect 734 1261 737 1268
rect 734 1258 750 1261
rect 802 1258 814 1261
rect 870 1261 873 1268
rect 866 1258 873 1261
rect 950 1261 953 1268
rect 946 1258 953 1261
rect 1090 1258 1134 1261
rect 1210 1258 1302 1261
rect 1306 1258 1310 1261
rect 1378 1258 1422 1261
rect 1502 1261 1506 1262
rect 1450 1258 1506 1261
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 18 1248 78 1251
rect 82 1248 142 1251
rect 146 1248 206 1251
rect 394 1248 582 1251
rect 590 1248 670 1251
rect 682 1248 814 1251
rect 914 1248 1065 1251
rect 1074 1248 1142 1251
rect 1194 1248 1246 1251
rect 1266 1248 1302 1251
rect 1306 1248 1350 1251
rect 1394 1248 1406 1251
rect 26 1238 62 1241
rect 122 1238 126 1241
rect 178 1238 190 1241
rect 590 1241 593 1248
rect 830 1242 833 1248
rect 306 1238 593 1241
rect 642 1238 742 1241
rect 1062 1241 1065 1248
rect 1062 1238 1086 1241
rect 1186 1238 1214 1241
rect 1362 1238 1398 1241
rect 10 1228 238 1231
rect 410 1228 486 1231
rect 514 1228 606 1231
rect 714 1228 798 1231
rect 826 1228 862 1231
rect 918 1231 921 1238
rect 890 1228 921 1231
rect 946 1228 966 1231
rect 1162 1228 1270 1231
rect 1354 1228 1366 1231
rect 266 1218 598 1221
rect 602 1218 1206 1221
rect 1218 1218 1262 1221
rect 1266 1218 1286 1221
rect 1290 1218 1390 1221
rect 74 1208 246 1211
rect 410 1208 430 1211
rect 586 1208 1102 1211
rect 1234 1208 1454 1211
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 486 1203 488 1207
rect 50 1198 270 1201
rect 434 1198 462 1201
rect 554 1198 734 1201
rect 746 1198 974 1201
rect 978 1198 1318 1201
rect 42 1188 382 1191
rect 386 1188 718 1191
rect 722 1188 1046 1191
rect 1114 1188 1230 1191
rect 1250 1188 1310 1191
rect 1354 1188 1382 1191
rect 1386 1188 1393 1191
rect 426 1178 502 1181
rect 570 1178 982 1181
rect 986 1178 1070 1181
rect 1138 1178 1286 1181
rect 1502 1181 1506 1182
rect 1362 1178 1506 1181
rect 126 1171 129 1178
rect 74 1168 129 1171
rect 186 1168 510 1171
rect 514 1168 598 1171
rect 618 1168 710 1171
rect 730 1168 798 1171
rect 802 1168 814 1171
rect 826 1168 830 1171
rect 838 1168 846 1171
rect 850 1168 902 1171
rect 914 1168 934 1171
rect 938 1168 945 1171
rect 962 1168 1006 1171
rect 1010 1168 1017 1171
rect 1026 1168 1062 1171
rect 1122 1168 1126 1171
rect 1210 1168 1238 1171
rect 1290 1168 1318 1171
rect 1330 1168 1430 1171
rect 114 1158 126 1161
rect 202 1158 206 1161
rect 458 1158 534 1161
rect 578 1158 622 1161
rect 658 1158 670 1161
rect 698 1158 702 1161
rect 706 1158 838 1161
rect 842 1158 862 1161
rect 866 1158 1030 1161
rect 1078 1161 1081 1168
rect 1078 1158 1182 1161
rect 1226 1158 1254 1161
rect 1282 1158 1286 1161
rect 1330 1158 1361 1161
rect 1502 1161 1506 1162
rect 1370 1158 1506 1161
rect 70 1152 73 1158
rect 102 1151 105 1158
rect 1358 1152 1361 1158
rect 102 1148 118 1151
rect 146 1148 190 1151
rect 450 1148 494 1151
rect 594 1148 654 1151
rect 658 1148 774 1151
rect 858 1148 902 1151
rect 914 1148 918 1151
rect 934 1148 942 1151
rect 946 1148 950 1151
rect 1090 1148 1094 1151
rect 1110 1148 1118 1151
rect 1122 1148 1126 1151
rect 1146 1148 1150 1151
rect 1250 1148 1342 1151
rect 1370 1148 1382 1151
rect 1442 1148 1454 1151
rect -26 1141 -22 1142
rect -26 1138 22 1141
rect 26 1138 30 1141
rect 34 1138 78 1141
rect 82 1138 94 1141
rect 330 1138 374 1141
rect 386 1138 566 1141
rect 626 1138 766 1141
rect 770 1138 862 1141
rect 866 1138 966 1141
rect 1090 1138 1190 1141
rect 1194 1138 1206 1141
rect 1226 1138 1262 1141
rect 1266 1138 1334 1141
rect 1338 1138 1422 1141
rect 66 1128 166 1131
rect 186 1128 230 1131
rect 234 1128 278 1131
rect 298 1128 302 1131
rect 338 1128 342 1131
rect 346 1128 446 1131
rect 490 1128 510 1131
rect 514 1128 582 1131
rect 610 1128 614 1131
rect 690 1128 790 1131
rect 794 1128 1094 1131
rect 1146 1128 1222 1131
rect 1298 1128 1377 1131
rect 82 1118 190 1121
rect 326 1121 329 1128
rect 1374 1122 1377 1128
rect 258 1118 374 1121
rect 378 1118 430 1121
rect 434 1118 518 1121
rect 614 1118 622 1121
rect 626 1118 678 1121
rect 762 1118 822 1121
rect 898 1118 918 1121
rect 962 1118 1062 1121
rect 1154 1118 1182 1121
rect 154 1108 166 1111
rect 282 1108 358 1111
rect 370 1108 406 1111
rect 418 1108 670 1111
rect 674 1108 726 1111
rect 746 1108 766 1111
rect 802 1108 814 1111
rect 826 1108 846 1111
rect 914 1108 958 1111
rect 1062 1111 1065 1118
rect 1062 1108 1446 1111
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 354 1098 366 1101
rect 370 1098 406 1101
rect 578 1098 614 1101
rect 770 1098 966 1101
rect 422 1092 425 1098
rect 10 1088 62 1091
rect 234 1088 414 1091
rect 546 1088 574 1091
rect 586 1088 630 1091
rect 682 1088 742 1091
rect 790 1088 798 1091
rect 802 1088 862 1091
rect 1282 1088 1342 1091
rect 1418 1088 1438 1091
rect -26 1081 -22 1082
rect -26 1078 6 1081
rect 10 1078 766 1081
rect 786 1078 838 1081
rect 846 1078 870 1081
rect 958 1078 998 1081
rect 1002 1078 1022 1081
rect 1274 1078 1310 1081
rect 1386 1078 1430 1081
rect 322 1068 374 1071
rect 378 1068 390 1071
rect 402 1068 454 1071
rect 466 1068 542 1071
rect 618 1068 622 1071
rect 634 1068 678 1071
rect 846 1071 849 1078
rect 958 1072 961 1078
rect 1390 1072 1393 1078
rect 738 1068 849 1071
rect 858 1068 878 1071
rect 946 1068 950 1071
rect 1154 1068 1158 1071
rect 1202 1068 1254 1071
rect 1290 1068 1326 1071
rect 1502 1071 1506 1072
rect 1450 1068 1506 1071
rect 98 1058 110 1061
rect 186 1058 222 1061
rect 242 1058 257 1061
rect 266 1058 302 1061
rect 398 1058 406 1061
rect 410 1058 414 1061
rect 538 1058 550 1061
rect 606 1061 609 1068
rect 602 1058 609 1061
rect 702 1061 705 1068
rect 702 1058 710 1061
rect 1022 1061 1025 1068
rect 1038 1061 1041 1068
rect 1022 1058 1041 1061
rect 1110 1061 1113 1068
rect 1110 1058 1126 1061
rect 1174 1061 1177 1068
rect 1174 1058 1190 1061
rect 1266 1058 1294 1061
rect 1366 1061 1369 1068
rect 1354 1058 1369 1061
rect -26 1051 -22 1052
rect -26 1048 6 1051
rect 50 1048 78 1051
rect 218 1048 230 1051
rect 254 1051 257 1058
rect 846 1052 849 1058
rect 254 1048 350 1051
rect 378 1048 718 1051
rect 934 1051 937 1058
rect 858 1048 937 1051
rect 994 1048 1054 1051
rect 1082 1048 1126 1051
rect 1154 1048 1214 1051
rect 1218 1048 1262 1051
rect 1322 1048 1406 1051
rect 1502 1051 1506 1052
rect 1482 1048 1506 1051
rect 50 1038 166 1041
rect 170 1038 270 1041
rect 274 1038 334 1041
rect 434 1038 494 1041
rect 514 1038 518 1041
rect 738 1038 742 1041
rect 834 1038 926 1041
rect 1034 1038 1086 1041
rect 1138 1038 1270 1041
rect 1314 1038 1342 1041
rect 1362 1038 1422 1041
rect 90 1028 110 1031
rect 154 1028 190 1031
rect 202 1028 246 1031
rect 258 1028 286 1031
rect 314 1028 414 1031
rect 834 1028 846 1031
rect 858 1028 878 1031
rect 890 1028 982 1031
rect 1010 1028 1446 1031
rect 58 1018 686 1021
rect 834 1018 1006 1021
rect 1018 1018 1382 1021
rect 1386 1018 1478 1021
rect 10 1008 94 1011
rect 98 1008 110 1011
rect 114 1008 150 1011
rect 154 1008 190 1011
rect 202 1008 206 1011
rect 362 1008 454 1011
rect 498 1008 606 1011
rect 874 1008 878 1011
rect 914 1008 961 1011
rect 978 1008 1038 1011
rect 1338 1008 1430 1011
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 486 1003 488 1007
rect -26 1001 -22 1002
rect -26 998 6 1001
rect 18 998 54 1001
rect 66 998 246 1001
rect 322 998 462 1001
rect 498 998 790 1001
rect 834 998 854 1001
rect 866 998 950 1001
rect 958 1001 961 1008
rect 958 998 1062 1001
rect 1306 998 1358 1001
rect 1502 1001 1506 1002
rect 1402 998 1506 1001
rect 18 988 30 991
rect 90 988 225 991
rect 314 988 390 991
rect 394 988 401 991
rect 410 988 734 991
rect 738 988 942 991
rect 946 988 1398 991
rect 222 982 225 988
rect -26 981 -22 982
rect -26 978 6 981
rect 10 978 126 981
rect 394 978 561 981
rect 658 978 718 981
rect 802 978 1014 981
rect 1066 978 1190 981
rect 1370 978 1446 981
rect 558 972 561 978
rect 42 968 70 971
rect 106 968 182 971
rect 242 968 326 971
rect 410 968 446 971
rect 498 968 502 971
rect 610 968 614 971
rect 650 968 670 971
rect 818 968 854 971
rect 858 968 1054 971
rect 1082 968 1097 971
rect 1258 968 1294 971
rect 1358 971 1361 978
rect 1354 968 1361 971
rect 1402 968 1438 971
rect 1502 968 1506 972
rect 30 962 33 968
rect 1094 962 1097 968
rect -26 961 -22 962
rect -26 958 14 961
rect 162 958 166 961
rect 174 958 214 961
rect 226 958 334 961
rect 426 958 430 961
rect 458 958 534 961
rect 922 958 958 961
rect 978 958 1038 961
rect 1106 958 1110 961
rect 1138 958 1142 961
rect 1162 958 1174 961
rect 1354 958 1358 961
rect 1502 961 1505 968
rect 1426 958 1505 961
rect 38 951 41 958
rect 34 948 41 951
rect 118 952 121 958
rect 142 951 145 958
rect 174 952 177 958
rect 142 948 158 951
rect 250 948 262 951
rect 542 951 545 958
rect 542 948 574 951
rect 598 951 601 958
rect 614 951 617 958
rect 598 948 617 951
rect 630 951 633 958
rect 646 951 649 958
rect 630 948 649 951
rect 686 951 689 958
rect 742 951 745 958
rect 686 948 745 951
rect 838 951 841 958
rect 894 952 897 958
rect 838 948 870 951
rect 978 948 982 951
rect 1034 948 1086 951
rect 1098 948 1102 951
rect 1130 948 1153 951
rect 1214 951 1217 958
rect 1202 948 1217 951
rect 1242 948 1254 951
rect 1290 948 1326 951
rect 1450 948 1470 951
rect 1502 951 1506 952
rect 1482 948 1506 951
rect 1150 942 1153 948
rect -26 941 -22 942
rect -26 938 126 941
rect 130 938 190 941
rect 202 938 254 941
rect 262 938 286 941
rect 290 938 326 941
rect 442 938 470 941
rect 474 938 510 941
rect 522 938 550 941
rect 578 938 742 941
rect 754 938 758 941
rect 762 938 950 941
rect 986 938 1022 941
rect 1058 938 1086 941
rect 1098 938 1142 941
rect 1154 938 1190 941
rect 1226 938 1230 941
rect 1354 938 1398 941
rect 1402 938 1414 941
rect 262 932 265 938
rect 50 928 54 931
rect 58 928 110 931
rect 170 928 190 931
rect 338 928 358 931
rect 366 928 374 931
rect 574 931 577 938
rect 378 928 577 931
rect 642 928 662 931
rect 706 928 766 931
rect 850 928 894 931
rect 914 928 998 931
rect 1002 928 1014 931
rect 1106 928 1254 931
rect 10 918 438 921
rect 530 918 582 921
rect 586 918 630 921
rect 702 921 705 928
rect 634 918 705 921
rect 1138 918 1182 921
rect 250 908 398 911
rect 554 908 638 911
rect 658 908 702 911
rect 1082 908 1278 911
rect 1290 908 1318 911
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 330 898 382 901
rect 402 898 638 901
rect 642 898 798 901
rect 1178 898 1262 901
rect 1278 901 1281 908
rect 1278 898 1438 901
rect 1442 898 1478 901
rect 806 892 809 898
rect -26 891 -22 892
rect -26 888 33 891
rect 354 888 614 891
rect 618 888 670 891
rect 682 888 742 891
rect 818 888 838 891
rect 882 888 934 891
rect 938 888 958 891
rect 970 888 1073 891
rect 1154 888 1166 891
rect 1234 888 1422 891
rect 1502 891 1506 892
rect 1462 888 1506 891
rect 30 882 33 888
rect 146 878 190 881
rect 218 878 270 881
rect 362 878 382 881
rect 450 878 534 881
rect 570 878 878 881
rect 914 878 998 881
rect 1018 878 1062 881
rect 1070 881 1073 888
rect 1070 878 1161 881
rect 1178 878 1222 881
rect 1266 878 1294 881
rect 1462 881 1465 888
rect 1298 878 1465 881
rect -26 871 -22 872
rect -26 868 14 871
rect 34 868 182 871
rect 186 868 238 871
rect 290 868 774 871
rect 902 871 905 878
rect 1158 872 1161 878
rect 778 868 958 871
rect 962 868 1030 871
rect 1050 868 1062 871
rect 1074 868 1110 871
rect 1194 868 1230 871
rect 1258 868 1262 871
rect 1266 868 1366 871
rect 1418 868 1438 871
rect 1502 871 1506 872
rect 1482 868 1506 871
rect -26 858 70 861
rect 82 858 94 861
rect 146 858 174 861
rect 202 858 206 861
rect 282 858 286 861
rect 298 858 302 861
rect 322 858 337 861
rect 354 858 369 861
rect 394 858 398 861
rect 418 858 742 861
rect 754 858 758 861
rect 770 858 830 861
rect 842 858 1046 861
rect 1050 858 1086 861
rect 1090 858 1118 861
rect 1322 858 1350 861
rect 1402 858 1438 861
rect -26 852 -23 858
rect -26 848 -22 852
rect 10 848 54 851
rect 58 848 102 851
rect 106 848 118 851
rect 214 851 217 858
rect 162 848 217 851
rect 262 852 265 858
rect 334 852 337 858
rect 366 852 369 858
rect 274 848 294 851
rect 394 848 446 851
rect 466 848 486 851
rect 602 848 606 851
rect 610 848 686 851
rect 706 848 934 851
rect 954 848 974 851
rect 1010 848 1094 851
rect 1098 848 1166 851
rect 1170 848 1358 851
rect 1362 848 1478 851
rect 1502 848 1506 852
rect 146 838 150 841
rect 170 838 310 841
rect 426 838 902 841
rect 1066 838 1254 841
rect 1258 838 1462 841
rect 1502 841 1505 848
rect 1466 838 1505 841
rect 114 828 169 831
rect 178 828 201 831
rect 226 828 278 831
rect 290 828 294 831
rect 458 828 502 831
rect 534 828 574 831
rect 730 828 782 831
rect 802 828 862 831
rect 1282 828 1329 831
rect 166 822 169 828
rect 198 822 201 828
rect 210 818 214 821
rect 218 818 225 821
rect 406 821 409 828
rect 234 818 409 821
rect 534 822 537 828
rect 1326 822 1329 828
rect 50 808 214 811
rect 514 808 686 811
rect 1234 808 1454 811
rect 472 803 474 807
rect 478 803 481 807
rect 486 803 488 807
rect -26 801 -22 802
rect -26 798 6 801
rect 26 798 174 801
rect 194 798 270 801
rect 666 798 726 801
rect 1502 801 1506 802
rect 1258 798 1506 801
rect 90 788 302 791
rect 506 788 622 791
rect 626 788 654 791
rect -26 781 -22 782
rect 6 781 9 788
rect -26 778 9 781
rect 694 781 697 788
rect 1310 782 1313 788
rect 642 778 697 781
rect 738 778 790 781
rect 1438 781 1441 788
rect 1502 781 1506 782
rect 1438 778 1506 781
rect 122 768 126 771
rect 290 768 510 771
rect 586 768 694 771
rect 714 768 750 771
rect 826 768 838 771
rect 1018 768 1030 771
rect 1082 768 1086 771
rect 1118 771 1121 778
rect 1118 768 1505 771
rect 1502 762 1505 768
rect -26 758 -22 762
rect 10 758 390 761
rect 634 758 646 761
rect 690 758 710 761
rect 758 758 1126 761
rect 1258 758 1294 761
rect 1306 758 1350 761
rect 1502 758 1506 762
rect -26 751 -23 758
rect 758 752 761 758
rect -26 748 6 751
rect 154 748 222 751
rect 418 748 430 751
rect 438 748 758 751
rect 770 748 1014 751
rect 1050 748 1078 751
rect 1098 748 1102 751
rect 1186 748 1262 751
rect 1314 748 1318 751
rect 94 742 97 748
rect 134 742 137 748
rect 438 742 441 748
rect 1278 742 1281 748
rect 1286 742 1289 748
rect -26 741 -22 742
rect -26 738 6 741
rect 178 738 438 741
rect 602 738 742 741
rect 746 738 782 741
rect 802 738 806 741
rect 818 738 838 741
rect 850 738 854 741
rect 866 738 870 741
rect 882 738 886 741
rect 938 738 942 741
rect 1066 738 1086 741
rect 1322 738 1334 741
rect 1502 741 1506 742
rect 1458 738 1506 741
rect 10 728 166 731
rect 442 728 454 731
rect 458 728 598 731
rect 794 728 814 731
rect 818 728 846 731
rect 850 728 878 731
rect 914 728 942 731
rect 1034 728 1070 731
rect 1090 728 1102 731
rect 1134 731 1137 738
rect 1134 728 1254 731
rect 1258 728 1286 731
rect -26 721 -22 722
rect -26 718 94 721
rect 98 718 206 721
rect 210 718 270 721
rect 274 718 326 721
rect 354 718 470 721
rect 570 718 806 721
rect 862 718 870 721
rect 882 718 910 721
rect 1170 718 1350 721
rect 90 708 174 711
rect 562 708 926 711
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 98 698 142 701
rect 546 698 830 701
rect 850 698 870 701
rect 1258 698 1262 701
rect -26 691 -22 692
rect -26 688 142 691
rect 154 688 182 691
rect 186 688 214 691
rect 626 688 662 691
rect 1502 691 1506 692
rect 1222 688 1506 691
rect 122 678 198 681
rect 614 681 617 688
rect 614 678 630 681
rect 642 678 646 681
rect 846 681 849 688
rect 1222 682 1225 688
rect 730 678 849 681
rect 1026 678 1118 681
rect -26 671 -22 672
rect 6 671 9 678
rect -26 668 9 671
rect 122 668 126 671
rect 162 668 166 671
rect 594 668 630 671
rect 674 668 678 671
rect 682 668 782 671
rect 1022 671 1025 678
rect 1302 672 1305 678
rect 1310 672 1313 678
rect 930 668 1025 671
rect 1250 668 1262 671
rect 1274 668 1278 671
rect 1346 668 1350 671
rect 1502 671 1506 672
rect 1482 668 1506 671
rect 26 658 129 661
rect 186 658 190 661
rect 218 658 254 661
rect 390 661 393 668
rect 390 658 422 661
rect 602 658 790 661
rect 806 661 809 668
rect 1038 662 1041 668
rect 806 658 822 661
rect 938 658 966 661
rect 1138 659 1142 661
rect 1198 661 1201 668
rect 1138 658 1145 659
rect 1198 658 1414 661
rect 126 652 129 658
rect 886 652 889 658
rect -26 651 -22 652
rect -26 648 6 651
rect 146 648 318 651
rect 378 648 510 651
rect 658 648 686 651
rect 742 648 766 651
rect 906 648 926 651
rect 978 648 1070 651
rect 1102 651 1105 658
rect 1102 648 1206 651
rect 1250 648 1254 651
rect 1418 648 1446 651
rect 1502 651 1506 652
rect 1494 648 1506 651
rect 742 642 745 648
rect 942 642 945 648
rect 130 638 158 641
rect 482 638 598 641
rect 682 638 686 641
rect 794 638 814 641
rect 842 638 870 641
rect 954 638 958 641
rect 994 638 1022 641
rect 1494 641 1497 648
rect 1438 638 1497 641
rect 438 631 441 638
rect 10 628 441 631
rect 702 631 705 638
rect 1438 632 1441 638
rect 702 628 758 631
rect 818 628 830 631
rect 842 628 974 631
rect 458 618 726 621
rect 730 618 790 621
rect 1286 621 1289 628
rect 1286 618 1366 621
rect -26 611 -22 612
rect -26 608 6 611
rect 66 608 102 611
rect 898 608 1134 611
rect 1290 608 1318 611
rect 472 603 474 607
rect 478 603 481 607
rect 486 603 488 607
rect 834 598 1222 601
rect -26 591 -22 592
rect -26 588 134 591
rect 138 588 526 591
rect 530 588 638 591
rect 650 588 734 591
rect 866 588 918 591
rect 922 588 1006 591
rect 1258 588 1278 591
rect 1282 588 1294 591
rect 10 578 422 581
rect 426 578 662 581
rect 754 578 774 581
rect 794 578 798 581
rect 810 578 902 581
rect 914 578 942 581
rect 1026 578 1062 581
rect 1226 578 1278 581
rect -26 571 -22 572
rect -26 568 38 571
rect 194 568 454 571
rect 522 568 550 571
rect 618 568 630 571
rect 642 568 686 571
rect 690 568 718 571
rect 770 568 838 571
rect 890 568 934 571
rect 938 568 1014 571
rect 1058 568 1190 571
rect 1266 568 1270 571
rect 282 558 286 561
rect 330 558 334 561
rect 350 558 494 561
rect 586 558 625 561
rect -26 551 -22 552
rect -26 548 70 551
rect 114 548 118 551
rect 318 551 321 558
rect 342 552 345 558
rect 350 552 353 558
rect 622 552 625 558
rect 746 558 769 561
rect 778 558 934 561
rect 938 558 1038 561
rect 1218 558 1222 561
rect 1242 558 1246 561
rect 318 548 326 551
rect 362 548 366 551
rect 386 548 518 551
rect 718 551 721 558
rect 718 548 734 551
rect 766 551 769 558
rect 766 548 849 551
rect 858 548 886 551
rect 954 548 958 551
rect 1078 551 1081 558
rect 1066 548 1081 551
rect 1202 548 1446 551
rect 1502 551 1506 552
rect 1482 548 1506 551
rect 42 538 310 541
rect 314 538 694 541
rect 698 538 758 541
rect 782 538 790 541
rect 794 538 806 541
rect 846 541 849 548
rect 846 538 862 541
rect 890 538 910 541
rect 966 541 969 548
rect 946 538 969 541
rect 978 538 982 541
rect 1034 538 1158 541
rect 1242 538 1254 541
rect 1290 538 1294 541
rect -26 531 -22 532
rect -26 528 62 531
rect 74 528 206 531
rect 210 528 238 531
rect 250 528 294 531
rect 362 528 366 531
rect 410 528 454 531
rect 474 528 590 531
rect 618 528 646 531
rect 650 528 678 531
rect 682 528 758 531
rect 890 528 1094 531
rect 1218 528 1238 531
rect 1502 531 1506 532
rect 1338 528 1506 531
rect 62 521 65 528
rect 62 518 254 521
rect 258 518 566 521
rect 570 518 582 521
rect 658 518 726 521
rect 738 518 1049 521
rect 34 508 94 511
rect 98 508 174 511
rect 178 508 198 511
rect 242 508 422 511
rect 434 508 582 511
rect 674 508 742 511
rect 746 508 790 511
rect 834 508 958 511
rect 1046 511 1049 518
rect 1430 512 1433 518
rect 1046 508 1174 511
rect 1178 508 1334 511
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 426 498 542 501
rect 554 498 734 501
rect 874 498 942 501
rect 1050 498 1286 501
rect 1306 498 1382 501
rect 1046 492 1049 498
rect -26 491 -22 492
rect -26 488 6 491
rect 10 488 534 491
rect 538 488 670 491
rect 682 488 830 491
rect 898 488 934 491
rect 1010 488 1038 491
rect 1098 488 1462 491
rect 1502 491 1506 492
rect 1466 488 1506 491
rect 130 478 134 481
rect 298 478 382 481
rect 450 478 566 481
rect 570 478 646 481
rect 650 478 694 481
rect 810 478 982 481
rect 1038 481 1041 488
rect 1038 478 1078 481
rect 1082 478 1102 481
rect 1106 478 1134 481
rect 1138 478 1206 481
rect 1210 478 1230 481
rect 1326 478 1334 481
rect 1338 478 1342 481
rect 1386 478 1473 481
rect 382 472 385 478
rect 1470 472 1473 478
rect -26 471 -22 472
rect -26 468 190 471
rect 306 468 318 471
rect 322 468 329 471
rect 338 468 374 471
rect 394 468 534 471
rect 642 468 646 471
rect 754 468 774 471
rect 890 468 910 471
rect 922 468 1094 471
rect 1130 468 1134 471
rect 1138 468 1302 471
rect 1306 468 1462 471
rect 50 458 81 461
rect 90 458 110 461
rect 170 458 177 461
rect 202 458 214 461
rect 262 461 265 468
rect 250 458 265 461
rect 282 458 390 461
rect 394 458 430 461
rect 442 458 510 461
rect 514 458 606 461
rect 662 461 665 468
rect 662 458 670 461
rect 762 458 790 461
rect 862 461 865 468
rect 862 458 870 461
rect 938 458 974 461
rect 978 458 1110 461
rect 1114 458 1150 461
rect 1266 458 1334 461
rect 1338 458 1390 461
rect 1434 458 1449 461
rect 78 452 81 458
rect 18 448 38 451
rect 106 448 222 451
rect 290 448 350 451
rect 386 448 390 451
rect 482 448 558 451
rect 622 451 625 458
rect 1446 452 1449 458
rect 622 448 662 451
rect 730 448 750 451
rect 774 448 782 451
rect 786 448 822 451
rect 842 448 942 451
rect 962 448 1222 451
rect 1266 448 1270 451
rect 1298 448 1358 451
rect 1502 451 1506 452
rect 1466 448 1506 451
rect 114 438 174 441
rect 186 438 238 441
rect 322 438 358 441
rect 418 438 422 441
rect 434 438 457 441
rect 538 438 550 441
rect 686 441 689 448
rect 686 438 702 441
rect 746 438 870 441
rect 938 438 942 441
rect 1082 438 1086 441
rect 1290 438 1302 441
rect 1322 438 1422 441
rect 454 432 457 438
rect 538 428 630 431
rect 874 428 918 431
rect 1090 428 1238 431
rect 1282 428 1294 431
rect 1354 428 1377 431
rect 1374 422 1377 428
rect 90 418 190 421
rect 386 418 462 421
rect 794 418 1038 421
rect 1250 418 1334 421
rect 58 408 166 411
rect 906 408 958 411
rect 962 408 1062 411
rect 472 403 474 407
rect 478 403 481 407
rect 486 403 488 407
rect 618 398 670 401
rect 786 398 950 401
rect 1314 398 1430 401
rect 114 388 134 391
rect 170 388 246 391
rect 250 388 294 391
rect 414 388 974 391
rect 978 388 1406 391
rect 414 382 417 388
rect 58 378 302 381
rect 330 378 414 381
rect 586 378 638 381
rect 818 378 1014 381
rect 1210 378 1361 381
rect 1386 378 1414 381
rect 58 368 70 371
rect 130 368 158 371
rect 194 368 238 371
rect 362 368 366 371
rect 526 371 529 378
rect 1358 372 1361 378
rect 514 368 529 371
rect 546 368 566 371
rect 570 368 598 371
rect 690 368 742 371
rect 842 368 846 371
rect 898 368 902 371
rect 930 368 966 371
rect 1082 368 1086 371
rect 1242 368 1246 371
rect 1362 368 1398 371
rect 1190 362 1193 368
rect 58 358 62 361
rect 402 358 454 361
rect 458 358 494 361
rect 498 358 622 361
rect 882 358 974 361
rect 1234 358 1270 361
rect 1282 358 1302 361
rect 1306 358 1318 361
rect 1338 358 1366 361
rect 1378 358 1401 361
rect 1422 361 1425 368
rect 1502 361 1506 362
rect 1410 358 1506 361
rect 30 351 33 358
rect 30 348 94 351
rect 222 351 225 358
rect 186 348 225 351
rect 238 351 241 358
rect 238 348 286 351
rect 394 348 406 351
rect 506 348 510 351
rect 522 348 550 351
rect 554 348 582 351
rect 586 348 630 351
rect 634 348 662 351
rect 754 348 774 351
rect 782 351 785 358
rect 778 348 806 351
rect 846 348 873 351
rect 938 348 942 351
rect 1058 348 1062 351
rect 1066 348 1102 351
rect 1142 351 1145 358
rect 1142 348 1158 351
rect 1174 351 1177 358
rect 1174 348 1190 351
rect 1242 348 1246 351
rect 1274 348 1286 351
rect 1290 348 1326 351
rect 1398 351 1401 358
rect 1378 348 1393 351
rect 1398 348 1454 351
rect 846 342 849 348
rect 870 342 873 348
rect 1390 342 1393 348
rect 18 338 70 341
rect 106 338 126 341
rect 214 338 257 341
rect 370 338 382 341
rect 386 338 422 341
rect 466 338 574 341
rect 610 338 630 341
rect 642 338 646 341
rect 818 338 825 341
rect 834 338 838 341
rect 906 338 950 341
rect 1002 338 1006 341
rect 1034 338 1086 341
rect 1122 338 1126 341
rect 1202 338 1278 341
rect 1314 338 1318 341
rect 1502 341 1506 342
rect 1410 338 1506 341
rect 214 332 217 338
rect 254 332 257 338
rect 90 328 166 331
rect 258 328 302 331
rect 306 328 310 331
rect 314 328 350 331
rect 378 328 433 331
rect 650 328 721 331
rect 778 328 814 331
rect 818 328 830 331
rect 850 328 862 331
rect 1018 328 1030 331
rect 1094 331 1097 338
rect 1190 332 1193 338
rect 1034 328 1110 331
rect 1114 328 1142 331
rect 1242 328 1246 331
rect 1306 328 1358 331
rect 430 322 433 328
rect 718 322 721 328
rect 50 318 118 321
rect 290 318 326 321
rect 330 318 382 321
rect 826 318 894 321
rect 1042 318 1222 321
rect 1266 318 1382 321
rect 1386 318 1414 321
rect 1426 318 1470 321
rect 114 308 206 311
rect 430 311 433 318
rect 430 308 758 311
rect 762 308 806 311
rect 1170 308 1214 311
rect 1258 308 1342 311
rect 1346 308 1406 311
rect 894 302 897 308
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 474 298 558 301
rect 1010 298 1014 301
rect 1018 298 1206 301
rect 1210 298 1238 301
rect 314 288 409 291
rect 406 282 409 288
rect 914 288 1070 291
rect 1226 288 1462 291
rect -26 281 -22 282
rect -26 278 62 281
rect 66 278 94 281
rect 98 278 134 281
rect 378 278 382 281
rect 418 278 542 281
rect 550 281 553 288
rect 546 278 553 281
rect 558 281 561 288
rect 558 278 582 281
rect 678 281 681 288
rect 610 278 681 281
rect 722 278 750 281
rect 794 278 798 281
rect 866 278 918 281
rect 930 278 934 281
rect 946 278 1030 281
rect 1130 278 1134 281
rect 1234 278 1358 281
rect 870 272 873 278
rect 50 268 110 271
rect 114 268 126 271
rect 178 268 198 271
rect 202 268 222 271
rect 290 268 334 271
rect 522 268 566 271
rect 594 268 630 271
rect 658 268 726 271
rect 730 268 782 271
rect 818 268 830 271
rect 914 268 926 271
rect 986 268 1278 271
rect -26 261 -22 262
rect -26 258 6 261
rect 10 258 38 261
rect 46 258 94 261
rect 98 258 158 261
rect 162 258 190 261
rect 278 261 281 268
rect 266 258 281 261
rect 306 258 310 261
rect 330 258 350 261
rect 354 258 374 261
rect 450 258 462 261
rect 474 258 542 261
rect 546 258 622 261
rect 690 258 694 261
rect 714 258 726 261
rect 778 258 902 261
rect 922 258 926 261
rect 946 258 950 261
rect 958 258 985 261
rect 1042 258 1102 261
rect 1186 258 1190 261
rect 1210 258 1262 261
rect 1294 261 1297 268
rect 1294 258 1302 261
rect 46 251 49 258
rect 958 252 961 258
rect 982 252 985 258
rect 42 248 49 251
rect 162 248 286 251
rect 346 248 374 251
rect 402 248 486 251
rect 490 248 798 251
rect 802 248 953 251
rect 1058 248 1078 251
rect 1090 248 1102 251
rect 1166 251 1169 258
rect 1166 248 1230 251
rect 90 238 110 241
rect 170 238 254 241
rect 274 238 318 241
rect 442 238 446 241
rect 538 238 622 241
rect 634 238 862 241
rect 950 241 953 248
rect 950 238 1014 241
rect 1058 238 1398 241
rect 130 228 382 231
rect 642 228 726 231
rect 862 231 865 238
rect 862 228 1174 231
rect 1182 228 1246 231
rect 1362 228 1430 231
rect 1182 222 1185 228
rect 26 218 134 221
rect 202 218 270 221
rect 362 218 598 221
rect 602 218 846 221
rect 850 218 1158 221
rect 1314 218 1430 221
rect 666 208 670 211
rect 754 208 894 211
rect 954 208 958 211
rect 1050 208 1142 211
rect 1146 208 1150 211
rect 472 203 474 207
rect 478 203 481 207
rect 486 203 488 207
rect 394 198 465 201
rect 570 198 590 201
rect 594 198 678 201
rect 686 198 798 201
rect 882 198 926 201
rect 938 198 1038 201
rect 1042 198 1182 201
rect 462 191 465 198
rect 462 188 542 191
rect 686 191 689 198
rect 642 188 689 191
rect 698 188 1046 191
rect 1082 188 1129 191
rect 1258 188 1286 191
rect 1290 188 1358 191
rect 454 182 457 188
rect 1126 182 1129 188
rect 466 178 518 181
rect 522 178 734 181
rect 738 178 822 181
rect 914 178 966 181
rect 1010 178 1046 181
rect 1202 178 1374 181
rect 1410 178 1430 181
rect 50 168 70 171
rect 74 168 158 171
rect 162 168 238 171
rect 242 168 262 171
rect 290 168 294 171
rect 466 168 606 171
rect 618 168 718 171
rect 746 168 774 171
rect 810 168 878 171
rect 938 168 982 171
rect 1002 168 1030 171
rect 1034 168 1041 171
rect 1066 168 1070 171
rect 1110 171 1113 178
rect 1074 168 1113 171
rect 1130 168 1134 171
rect 1170 168 1390 171
rect 114 158 190 161
rect 274 158 326 161
rect 378 158 398 161
rect 442 158 510 161
rect 514 158 542 161
rect 546 158 654 161
rect 682 158 710 161
rect 738 158 798 161
rect 930 158 934 161
rect 954 158 958 161
rect 962 158 1102 161
rect 1106 158 1134 161
rect 1282 158 1302 161
rect 1386 158 1422 161
rect -26 151 -22 152
rect -26 148 57 151
rect 102 151 105 158
rect 82 148 105 151
rect 162 148 169 151
rect 258 148 294 151
rect 330 148 646 151
rect 762 148 806 151
rect 846 151 849 158
rect 818 148 849 151
rect 874 148 1022 151
rect 1026 148 1038 151
rect 1058 148 1062 151
rect 1158 151 1161 158
rect 1154 148 1161 151
rect 1186 148 1206 151
rect 1210 148 1238 151
rect 1298 148 1310 151
rect 1350 151 1353 158
rect 1350 148 1358 151
rect 1402 148 1406 151
rect 1502 148 1506 152
rect 54 142 57 148
rect 166 142 169 148
rect 18 138 41 141
rect 58 138 62 141
rect 122 138 126 141
rect 178 138 230 141
rect 242 138 254 141
rect 274 138 486 141
rect 490 138 534 141
rect 546 138 918 141
rect 922 138 1190 141
rect 1194 138 1406 141
rect 1502 141 1505 148
rect 1410 138 1505 141
rect 38 132 41 138
rect 50 128 54 131
rect 114 128 118 131
rect 298 128 350 131
rect 354 128 382 131
rect 418 128 742 131
rect 802 128 830 131
rect 838 128 894 131
rect 954 128 1006 131
rect 1026 128 1086 131
rect 1162 128 1222 131
rect 1394 128 1422 131
rect 838 122 841 128
rect 870 122 873 128
rect 1430 122 1433 128
rect 194 118 438 121
rect 450 118 534 121
rect 562 118 574 121
rect 578 118 585 121
rect 634 118 670 121
rect 698 118 758 121
rect 770 118 782 121
rect 786 118 838 121
rect 966 118 1022 121
rect 1034 118 1094 121
rect 1122 118 1166 121
rect 1182 118 1270 121
rect 1354 118 1414 121
rect 966 112 969 118
rect 218 108 382 111
rect 442 108 798 111
rect 858 108 966 111
rect 1010 108 1030 111
rect 1182 111 1185 118
rect 1098 108 1185 111
rect 1194 108 1318 111
rect 1370 108 1446 111
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect -26 101 -22 102
rect -26 98 70 101
rect 202 98 222 101
rect 282 98 862 101
rect 1090 98 1222 101
rect 1242 98 1406 101
rect 170 88 470 91
rect 474 88 526 91
rect 546 88 606 91
rect 662 88 670 91
rect 682 88 750 91
rect 754 88 854 91
rect 862 91 865 98
rect 862 88 1174 91
rect 1178 88 1334 91
rect 74 78 78 81
rect 106 78 126 81
rect 130 78 134 81
rect 138 78 182 81
rect 202 78 270 81
rect 274 78 342 81
rect 354 78 377 81
rect 450 78 502 81
rect 542 81 545 88
rect 662 82 665 88
rect 506 78 545 81
rect 842 78 846 81
rect 930 78 942 81
rect 946 78 950 81
rect 1002 78 1030 81
rect 1130 78 1134 81
rect 1502 81 1506 82
rect 1466 78 1506 81
rect 50 68 94 71
rect 170 68 174 71
rect 234 68 262 71
rect 274 68 278 71
rect 330 68 366 71
rect 374 71 377 78
rect 622 71 625 78
rect 774 72 777 78
rect 1038 72 1041 78
rect 1358 72 1361 78
rect 374 68 625 71
rect 666 68 678 71
rect 682 68 758 71
rect 762 68 766 71
rect 818 68 830 71
rect 834 68 862 71
rect 866 68 894 71
rect 898 68 966 71
rect 970 68 1006 71
rect 1082 68 1094 71
rect 1098 68 1118 71
rect 1122 68 1158 71
rect 1162 68 1182 71
rect 1266 68 1342 71
rect 934 62 937 68
rect 10 58 398 61
rect 402 58 510 61
rect 522 58 534 61
rect 634 58 702 61
rect 706 58 838 61
rect 890 58 910 61
rect 1034 58 1038 61
rect 1058 58 1086 61
rect 1106 58 1110 61
rect 1194 58 1206 61
rect 1218 58 1246 61
rect 1250 58 1302 61
rect 1306 58 1334 61
rect 1338 58 1382 61
rect -26 51 -22 52
rect 6 51 9 58
rect -26 48 9 51
rect 138 48 334 51
rect 482 48 494 51
rect 506 48 510 51
rect 610 48 622 51
rect 838 51 841 58
rect 838 48 1270 51
rect 1314 48 1326 51
rect 1346 48 1358 51
rect 1502 51 1506 52
rect 1418 48 1506 51
rect 250 38 286 41
rect 374 41 377 48
rect 374 38 638 41
rect 642 38 886 41
rect 890 38 1318 41
rect 322 28 710 31
rect 714 28 1022 31
rect 1026 28 1174 31
rect 394 18 574 21
rect 586 18 590 21
rect 602 18 638 21
rect 746 18 1254 21
rect 374 12 377 18
rect 66 8 86 11
rect 90 8 166 11
rect 574 11 577 18
rect 574 8 598 11
rect 602 8 630 11
rect 650 8 662 11
rect 818 8 910 11
rect 914 8 918 11
rect 1146 8 1150 11
rect 472 3 474 7
rect 478 3 481 7
rect 486 3 488 7
<< m4contact >>
rect 430 1408 434 1412
rect 1190 1408 1194 1412
rect 1310 1408 1314 1412
rect 474 1403 478 1407
rect 482 1403 485 1407
rect 485 1403 486 1407
rect 494 1398 498 1402
rect 494 1378 498 1382
rect 502 1368 506 1372
rect 518 1368 522 1372
rect 550 1358 554 1362
rect 590 1358 594 1362
rect 630 1358 634 1362
rect 646 1358 650 1362
rect 734 1358 738 1362
rect 934 1358 938 1362
rect 270 1348 274 1352
rect 334 1348 338 1352
rect 614 1348 618 1352
rect 894 1348 898 1352
rect 1262 1338 1266 1342
rect 1382 1338 1386 1342
rect 302 1328 306 1332
rect 774 1328 778 1332
rect 846 1328 850 1332
rect 1318 1328 1322 1332
rect 646 1318 650 1322
rect 694 1318 698 1322
rect 918 1318 922 1322
rect 1078 1318 1082 1322
rect 1198 1318 1202 1322
rect 1222 1308 1226 1312
rect 1358 1308 1362 1312
rect 986 1303 990 1307
rect 994 1303 997 1307
rect 997 1303 998 1307
rect 382 1298 386 1302
rect 518 1288 522 1292
rect 622 1288 626 1292
rect 726 1288 730 1292
rect 846 1278 850 1282
rect 998 1278 1002 1282
rect 1190 1278 1194 1282
rect 1198 1278 1202 1282
rect 270 1268 274 1272
rect 206 1258 210 1262
rect 798 1258 802 1262
rect 1206 1258 1210 1262
rect 1302 1258 1306 1262
rect 670 1248 674 1252
rect 830 1248 834 1252
rect 1358 1238 1362 1242
rect 798 1228 802 1232
rect 862 1228 866 1232
rect 1206 1218 1210 1222
rect 1262 1218 1266 1222
rect 70 1208 74 1212
rect 430 1208 434 1212
rect 474 1203 478 1207
rect 482 1203 485 1207
rect 485 1203 486 1207
rect 734 1198 738 1202
rect 742 1198 746 1202
rect 1318 1198 1322 1202
rect 502 1178 506 1182
rect 1286 1178 1290 1182
rect 598 1168 602 1172
rect 814 1168 818 1172
rect 822 1168 826 1172
rect 1062 1168 1066 1172
rect 1126 1168 1130 1172
rect 1326 1168 1330 1172
rect 206 1158 210 1162
rect 622 1158 626 1162
rect 702 1158 706 1162
rect 1222 1158 1226 1162
rect 1278 1158 1282 1162
rect 70 1148 74 1152
rect 494 1148 498 1152
rect 910 1148 914 1152
rect 1086 1148 1090 1152
rect 1142 1148 1146 1152
rect 1342 1148 1346 1152
rect 1366 1148 1370 1152
rect 30 1138 34 1142
rect 382 1138 386 1142
rect 278 1128 282 1132
rect 334 1128 338 1132
rect 606 1128 610 1132
rect 822 1118 826 1122
rect 958 1118 962 1122
rect 406 1108 410 1112
rect 414 1108 418 1112
rect 726 1108 730 1112
rect 986 1103 990 1107
rect 994 1103 997 1107
rect 997 1103 998 1107
rect 614 1098 618 1102
rect 414 1088 418 1092
rect 422 1088 426 1092
rect 1278 1088 1282 1092
rect 1270 1078 1274 1082
rect 1382 1078 1386 1082
rect 462 1068 466 1072
rect 622 1068 626 1072
rect 950 1068 954 1072
rect 1158 1068 1162 1072
rect 1326 1068 1330 1072
rect 846 1058 850 1062
rect 1262 1048 1266 1052
rect 1478 1048 1482 1052
rect 830 1038 834 1042
rect 190 1028 194 1032
rect 854 1028 858 1032
rect 982 1028 986 1032
rect 830 1018 834 1022
rect 1478 1018 1482 1022
rect 198 1008 202 1012
rect 454 1008 458 1012
rect 878 1008 882 1012
rect 974 1008 978 1012
rect 474 1003 478 1007
rect 482 1003 485 1007
rect 485 1003 486 1007
rect 14 998 18 1002
rect 462 998 466 1002
rect 494 998 498 1002
rect 854 998 858 1002
rect 1358 998 1362 1002
rect 6 978 10 982
rect 798 978 802 982
rect 406 968 410 972
rect 502 968 506 972
rect 606 968 610 972
rect 814 968 818 972
rect 14 958 18 962
rect 30 958 34 962
rect 166 958 170 962
rect 430 958 434 962
rect 454 958 458 962
rect 894 958 898 962
rect 1038 958 1042 962
rect 1102 958 1106 962
rect 1142 958 1146 962
rect 1158 958 1162 962
rect 1358 958 1362 962
rect 118 948 122 952
rect 1086 948 1090 952
rect 1094 948 1098 952
rect 1478 948 1482 952
rect 190 938 194 942
rect 742 938 746 942
rect 758 938 762 942
rect 950 938 954 942
rect 982 938 986 942
rect 1094 938 1098 942
rect 1230 938 1234 942
rect 1102 928 1106 932
rect 1134 918 1138 922
rect 986 903 990 907
rect 994 903 997 907
rect 997 903 998 907
rect 398 898 402 902
rect 798 898 802 902
rect 1478 898 1482 902
rect 670 888 674 892
rect 806 888 810 892
rect 958 888 962 892
rect 142 878 146 882
rect 878 878 882 882
rect 910 878 914 882
rect 1174 878 1178 882
rect 30 868 34 872
rect 1070 868 1074 872
rect 1262 868 1266 872
rect 174 858 178 862
rect 198 858 202 862
rect 278 858 282 862
rect 294 858 298 862
rect 350 858 354 862
rect 398 858 402 862
rect 758 858 762 862
rect 830 858 834 862
rect 6 848 10 852
rect 262 848 266 852
rect 702 848 706 852
rect 142 838 146 842
rect 294 828 298 832
rect 206 818 210 822
rect 1230 808 1234 812
rect 474 803 478 807
rect 482 803 485 807
rect 485 803 486 807
rect 6 798 10 802
rect 190 798 194 802
rect 1310 778 1314 782
rect 126 768 130 772
rect 1030 768 1034 772
rect 1086 768 1090 772
rect 6 758 10 762
rect 1254 758 1258 762
rect 94 748 98 752
rect 1102 748 1106 752
rect 1286 748 1290 752
rect 1318 748 1322 752
rect 6 738 10 742
rect 134 738 138 742
rect 806 738 810 742
rect 838 738 842 742
rect 854 738 858 742
rect 862 738 866 742
rect 886 738 890 742
rect 934 738 938 742
rect 1278 738 1282 742
rect 1086 728 1090 732
rect 870 718 874 722
rect 878 718 882 722
rect 986 703 990 707
rect 994 703 997 707
rect 997 703 998 707
rect 94 698 98 702
rect 846 698 850 702
rect 1262 698 1266 702
rect 142 688 146 692
rect 118 678 122 682
rect 630 678 634 682
rect 1302 678 1306 682
rect 118 668 122 672
rect 166 668 170 672
rect 670 668 674 672
rect 1270 668 1274 672
rect 1310 668 1314 672
rect 1342 668 1346 672
rect 190 658 194 662
rect 790 658 794 662
rect 886 658 890 662
rect 1038 658 1042 662
rect 1134 658 1138 662
rect 6 648 10 652
rect 142 648 146 652
rect 1254 648 1258 652
rect 686 638 690 642
rect 790 638 794 642
rect 942 638 946 642
rect 950 638 954 642
rect 6 628 10 632
rect 838 628 842 632
rect 474 603 478 607
rect 482 603 485 607
rect 485 603 486 607
rect 1222 598 1226 602
rect 918 588 922 592
rect 1278 588 1282 592
rect 790 578 794 582
rect 902 578 906 582
rect 630 568 634 572
rect 934 568 938 572
rect 286 558 290 562
rect 326 558 330 562
rect 342 558 346 562
rect 110 548 114 552
rect 1214 558 1218 562
rect 1238 558 1242 562
rect 358 548 362 552
rect 958 548 962 552
rect 886 538 890 542
rect 982 538 986 542
rect 1254 538 1258 542
rect 1294 538 1298 542
rect 238 528 242 532
rect 366 528 370 532
rect 470 528 474 532
rect 678 528 682 532
rect 886 528 890 532
rect 726 518 730 522
rect 422 508 426 512
rect 670 508 674 512
rect 1430 518 1434 522
rect 986 503 990 507
rect 994 503 997 507
rect 997 503 998 507
rect 1046 498 1050 502
rect 670 488 674 492
rect 134 478 138 482
rect 382 478 386 482
rect 374 468 378 472
rect 390 468 394 472
rect 646 468 650 472
rect 1134 468 1138 472
rect 1462 468 1466 472
rect 430 458 434 462
rect 510 458 514 462
rect 390 448 394 452
rect 726 448 730 452
rect 822 448 826 452
rect 958 448 962 452
rect 1262 448 1266 452
rect 1462 448 1466 452
rect 110 438 114 442
rect 422 438 426 442
rect 942 438 946 442
rect 1286 438 1290 442
rect 1086 428 1090 432
rect 1294 428 1298 432
rect 190 418 194 422
rect 1246 418 1250 422
rect 474 403 478 407
rect 482 403 485 407
rect 485 403 486 407
rect 974 388 978 392
rect 54 378 58 382
rect 1014 378 1018 382
rect 838 368 842 372
rect 894 368 898 372
rect 1078 368 1082 372
rect 1190 368 1194 372
rect 1238 368 1242 372
rect 62 358 66 362
rect 454 358 458 362
rect 1278 358 1282 362
rect 1406 358 1410 362
rect 502 348 506 352
rect 582 348 586 352
rect 942 348 946 352
rect 1054 348 1058 352
rect 1158 348 1162 352
rect 1246 348 1250 352
rect 382 338 386 342
rect 646 338 650 342
rect 814 338 818 342
rect 830 338 834 342
rect 1006 338 1010 342
rect 1086 338 1090 342
rect 1126 338 1130 342
rect 1190 338 1194 342
rect 1318 338 1322 342
rect 1238 328 1242 332
rect 382 318 386 322
rect 1038 318 1042 322
rect 894 308 898 312
rect 1254 308 1258 312
rect 1406 308 1410 312
rect 986 303 990 307
rect 994 303 997 307
rect 997 303 998 307
rect 1014 298 1018 302
rect 550 288 554 292
rect 374 278 378 282
rect 798 278 802 282
rect 862 278 866 282
rect 926 278 930 282
rect 1134 278 1138 282
rect 174 268 178 272
rect 286 268 290 272
rect 310 258 314 262
rect 462 258 466 262
rect 686 258 690 262
rect 902 258 906 262
rect 926 258 930 262
rect 942 258 946 262
rect 1182 258 1186 262
rect 286 248 290 252
rect 110 238 114 242
rect 630 238 634 242
rect 1054 238 1058 242
rect 638 228 642 232
rect 846 218 850 222
rect 662 208 666 212
rect 950 208 954 212
rect 1142 208 1146 212
rect 474 203 478 207
rect 482 203 485 207
rect 485 203 486 207
rect 454 188 458 192
rect 1078 188 1082 192
rect 1358 188 1362 192
rect 462 178 466 182
rect 1006 178 1010 182
rect 1406 178 1410 182
rect 462 168 466 172
rect 606 168 610 172
rect 806 168 810 172
rect 934 168 938 172
rect 1134 168 1138 172
rect 510 158 514 162
rect 926 158 930 162
rect 950 158 954 162
rect 806 148 810 152
rect 870 148 874 152
rect 1038 148 1042 152
rect 1054 148 1058 152
rect 1294 148 1298 152
rect 1406 148 1410 152
rect 54 138 58 142
rect 118 138 122 142
rect 254 138 258 142
rect 270 138 274 142
rect 534 138 538 142
rect 110 128 114 132
rect 830 128 834 132
rect 1006 128 1010 132
rect 1022 128 1026 132
rect 1430 128 1434 132
rect 758 118 762 122
rect 798 108 802 112
rect 854 108 858 112
rect 1006 108 1010 112
rect 986 103 990 107
rect 994 103 997 107
rect 997 103 998 107
rect 70 98 74 102
rect 278 98 282 102
rect 1406 98 1410 102
rect 526 88 530 92
rect 670 88 674 92
rect 678 88 682 92
rect 854 88 858 92
rect 70 78 74 82
rect 774 78 778 82
rect 838 78 842 82
rect 950 78 954 82
rect 1030 78 1034 82
rect 1126 78 1130 82
rect 166 68 170 72
rect 278 68 282 72
rect 1006 68 1010 72
rect 1038 68 1042 72
rect 1342 68 1346 72
rect 1358 68 1362 72
rect 510 58 514 62
rect 838 58 842 62
rect 1038 58 1042 62
rect 1102 58 1106 62
rect 606 48 610 52
rect 1342 48 1346 52
rect 374 18 378 22
rect 590 18 594 22
rect 166 8 170 12
rect 630 8 634 12
rect 918 8 922 12
rect 1142 8 1146 12
rect 474 3 478 7
rect 482 3 485 7
rect 485 3 486 7
<< metal4 >>
rect 1302 1408 1310 1411
rect 270 1272 273 1348
rect 306 1328 310 1331
rect 70 1152 73 1208
rect 206 1162 209 1258
rect 6 852 9 978
rect 14 962 17 998
rect 30 962 33 1138
rect 334 1132 337 1348
rect 382 1142 385 1298
rect 430 1212 433 1408
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 486 1403 488 1407
rect 494 1382 497 1398
rect 506 1368 510 1371
rect 518 1292 521 1368
rect 934 1362 937 1368
rect 622 1358 630 1361
rect 642 1358 646 1361
rect 550 1342 553 1358
rect 590 1352 593 1358
rect 614 1352 617 1358
rect 622 1292 625 1358
rect 698 1318 705 1321
rect 646 1282 649 1318
rect 670 1252 673 1268
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 486 1203 488 1207
rect 282 1128 286 1131
rect 190 1021 193 1028
rect 190 1018 201 1021
rect 198 1012 201 1018
rect 406 972 409 1108
rect 414 1092 417 1108
rect 422 961 425 1088
rect 454 962 457 1008
rect 462 1002 465 1068
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 486 1003 488 1007
rect 494 1002 497 1148
rect 502 972 505 1178
rect 598 1162 601 1168
rect 702 1162 705 1318
rect 622 1142 625 1158
rect 726 1152 729 1288
rect 734 1202 737 1358
rect 890 1348 894 1351
rect 846 1332 849 1338
rect 770 1328 774 1331
rect 798 1232 801 1258
rect 610 1128 614 1131
rect 614 971 617 1098
rect 622 1072 625 1138
rect 726 1112 729 1148
rect 610 968 617 971
rect 422 958 430 961
rect 30 872 33 958
rect 10 798 14 801
rect 6 742 9 758
rect 94 702 97 748
rect 118 682 121 948
rect 142 842 145 878
rect 126 671 129 768
rect 122 668 129 671
rect 6 632 9 648
rect 110 442 113 548
rect 134 482 137 738
rect 142 652 145 688
rect 166 672 169 958
rect 742 942 745 1198
rect 194 938 198 941
rect 754 938 758 941
rect 206 861 209 868
rect 398 862 401 898
rect 670 892 673 928
rect 798 902 801 978
rect 814 972 817 1168
rect 822 1122 825 1168
rect 830 1042 833 1248
rect 846 1062 849 1278
rect 202 858 209 861
rect 282 858 286 861
rect 346 858 350 861
rect 754 858 758 861
rect 174 832 177 858
rect 266 848 270 851
rect 294 832 297 858
rect 698 848 702 851
rect 206 822 209 828
rect 472 803 474 807
rect 478 803 481 807
rect 486 803 488 807
rect 186 798 190 801
rect 806 742 809 888
rect 830 862 833 1018
rect 854 1002 857 1028
rect 862 742 865 1228
rect 874 1008 878 1011
rect 894 962 897 1348
rect 918 1162 921 1318
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 994 1278 998 1281
rect 1066 1168 1070 1171
rect 918 1151 921 1158
rect 914 1148 921 1151
rect 1078 1132 1081 1318
rect 1190 1282 1193 1408
rect 1198 1282 1201 1318
rect 1190 1272 1193 1278
rect 1206 1222 1209 1258
rect 1122 1168 1126 1171
rect 1222 1162 1225 1308
rect 1262 1222 1265 1338
rect 1302 1262 1305 1408
rect 1318 1202 1321 1328
rect 1358 1242 1361 1308
rect 1286 1161 1289 1178
rect 1282 1158 1289 1161
rect 1090 1148 1097 1151
rect 1146 1148 1150 1151
rect 1094 1142 1097 1148
rect 950 942 953 1068
rect 958 892 961 1118
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 1154 1068 1158 1071
rect 970 1008 974 1011
rect 982 942 985 1028
rect 1038 962 1041 968
rect 1158 962 1161 968
rect 1134 958 1142 961
rect 1094 952 1097 958
rect 1086 941 1089 948
rect 1086 938 1094 941
rect 1102 932 1105 958
rect 1134 922 1137 958
rect 1230 932 1233 938
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 874 878 878 881
rect 1170 878 1174 881
rect 910 872 913 878
rect 1070 862 1073 868
rect 1230 812 1233 928
rect 1262 872 1265 1048
rect 1030 752 1033 768
rect 846 738 854 741
rect 878 738 886 741
rect 938 738 942 741
rect 630 672 633 678
rect 674 668 681 671
rect 190 422 193 658
rect 472 603 474 607
rect 478 603 481 607
rect 486 603 488 607
rect 630 572 633 578
rect 290 558 294 561
rect 330 558 334 561
rect 342 552 345 558
rect 354 548 358 551
rect 678 532 681 668
rect 794 658 798 661
rect 690 638 694 641
rect 786 638 790 641
rect 838 632 841 738
rect 846 702 849 738
rect 870 722 873 738
rect 878 722 881 738
rect 1086 732 1089 768
rect 1098 748 1102 751
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 1254 701 1257 758
rect 1254 698 1262 701
rect 1270 672 1273 1078
rect 1278 742 1281 1088
rect 1326 1072 1329 1168
rect 1346 1148 1350 1151
rect 1362 1148 1366 1151
rect 1382 1082 1385 1338
rect 1478 1022 1481 1048
rect 1358 962 1361 998
rect 1478 902 1481 948
rect 1038 662 1041 668
rect 1130 658 1134 661
rect 794 578 798 581
rect 886 542 889 658
rect 1246 648 1254 651
rect 902 562 905 578
rect 362 528 366 531
rect 466 528 470 531
rect 238 492 241 528
rect 374 472 377 478
rect 54 361 57 378
rect 54 358 62 361
rect 382 342 385 478
rect 390 452 393 468
rect 422 442 425 508
rect 670 492 673 508
rect 646 472 649 478
rect 430 462 433 468
rect 472 403 474 407
rect 478 403 481 407
rect 486 403 488 407
rect 386 318 390 321
rect 58 138 62 141
rect 110 132 113 238
rect 118 132 121 138
rect 70 82 73 98
rect 74 78 78 81
rect 174 71 177 268
rect 286 252 289 268
rect 314 258 318 261
rect 254 142 257 168
rect 266 138 270 141
rect 170 68 177 71
rect 278 72 281 98
rect 166 12 169 68
rect 374 22 377 278
rect 454 192 457 358
rect 510 351 513 458
rect 726 452 729 518
rect 886 482 889 528
rect 826 448 830 451
rect 842 368 849 371
rect 506 348 513 351
rect 462 182 465 258
rect 472 203 474 207
rect 478 203 481 207
rect 486 203 488 207
rect 458 168 462 171
rect 510 162 513 348
rect 550 282 553 288
rect 534 142 537 148
rect 526 92 529 138
rect 510 62 513 68
rect 582 21 585 348
rect 638 338 646 341
rect 818 338 822 341
rect 606 172 609 198
rect 606 52 609 168
rect 582 18 590 21
rect 630 12 633 238
rect 638 232 641 338
rect 830 332 833 338
rect 798 272 801 278
rect 690 258 694 261
rect 666 208 673 211
rect 670 92 673 208
rect 758 122 761 128
rect 798 112 801 268
rect 830 202 833 328
rect 846 222 849 368
rect 894 312 897 368
rect 806 152 809 168
rect 830 132 833 158
rect 862 142 865 278
rect 906 258 910 261
rect 918 261 921 588
rect 926 272 929 278
rect 918 258 926 261
rect 874 148 878 151
rect 854 92 857 108
rect 678 82 681 88
rect 774 72 777 78
rect 838 62 841 78
rect 918 12 921 258
rect 934 172 937 568
rect 942 442 945 638
rect 942 262 945 348
rect 950 212 953 638
rect 1222 561 1225 598
rect 1218 558 1225 561
rect 1234 558 1238 561
rect 958 452 961 548
rect 974 538 982 541
rect 974 392 977 538
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 1046 492 1049 498
rect 1130 468 1134 471
rect 1002 338 1006 341
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 1014 302 1017 378
rect 1034 318 1038 321
rect 1054 242 1057 348
rect 930 158 934 161
rect 950 82 953 158
rect 1006 132 1009 178
rect 1054 152 1057 238
rect 1078 192 1081 368
rect 1086 342 1089 428
rect 1246 422 1249 648
rect 1162 348 1166 351
rect 1190 342 1193 368
rect 1126 332 1129 338
rect 1238 332 1241 368
rect 1246 352 1249 358
rect 1254 312 1257 538
rect 1266 448 1270 451
rect 1278 362 1281 588
rect 1286 442 1289 748
rect 1302 672 1305 678
rect 1310 672 1313 778
rect 1294 432 1297 538
rect 1318 342 1321 748
rect 1346 668 1350 671
rect 1406 312 1409 358
rect 1130 278 1134 281
rect 1042 148 1046 151
rect 1018 128 1022 131
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect 1006 72 1009 108
rect 1030 82 1033 88
rect 1126 82 1129 278
rect 1186 258 1190 261
rect 1134 92 1137 168
rect 1034 68 1038 71
rect 1042 58 1046 61
rect 1106 58 1110 61
rect 1142 12 1145 208
rect 1290 148 1294 151
rect 1358 72 1361 188
rect 1406 182 1409 308
rect 1406 102 1409 148
rect 1430 132 1433 518
rect 1462 452 1465 468
rect 1342 52 1345 68
rect 472 3 474 7
rect 478 3 481 7
rect 486 3 488 7
<< m5contact >>
rect 310 1328 314 1332
rect 474 1403 478 1407
rect 481 1403 482 1407
rect 482 1403 485 1407
rect 510 1368 514 1372
rect 934 1368 938 1372
rect 614 1358 618 1362
rect 638 1358 642 1362
rect 590 1348 594 1352
rect 550 1338 554 1342
rect 646 1278 650 1282
rect 670 1268 674 1272
rect 474 1203 478 1207
rect 481 1203 482 1207
rect 482 1203 485 1207
rect 286 1128 290 1132
rect 474 1003 478 1007
rect 481 1003 482 1007
rect 482 1003 485 1007
rect 598 1158 602 1162
rect 886 1348 890 1352
rect 846 1338 850 1342
rect 766 1328 770 1332
rect 726 1148 730 1152
rect 622 1138 626 1142
rect 614 1128 618 1132
rect 14 798 18 802
rect 198 938 202 942
rect 750 938 754 942
rect 670 928 674 932
rect 206 868 210 872
rect 286 858 290 862
rect 342 858 346 862
rect 750 858 754 862
rect 270 848 274 852
rect 694 848 698 852
rect 174 828 178 832
rect 206 828 210 832
rect 474 803 478 807
rect 481 803 482 807
rect 482 803 485 807
rect 182 798 186 802
rect 870 1008 874 1012
rect 986 1303 990 1307
rect 993 1303 994 1307
rect 994 1303 997 1307
rect 990 1278 994 1282
rect 1070 1168 1074 1172
rect 918 1158 922 1162
rect 1190 1268 1194 1272
rect 1118 1168 1122 1172
rect 1150 1148 1154 1152
rect 1094 1138 1098 1142
rect 1078 1128 1082 1132
rect 950 1068 954 1072
rect 894 958 898 962
rect 986 1103 990 1107
rect 993 1103 994 1107
rect 994 1103 997 1107
rect 1150 1068 1154 1072
rect 966 1008 970 1012
rect 1038 968 1042 972
rect 1158 968 1162 972
rect 1094 958 1098 962
rect 1230 928 1234 932
rect 986 903 990 907
rect 993 903 994 907
rect 994 903 997 907
rect 870 878 874 882
rect 1166 878 1170 882
rect 910 868 914 872
rect 1070 858 1074 862
rect 1030 748 1034 752
rect 870 738 874 742
rect 942 738 946 742
rect 630 668 634 672
rect 474 603 478 607
rect 481 603 482 607
rect 482 603 485 607
rect 630 578 634 582
rect 294 558 298 562
rect 334 558 338 562
rect 342 548 346 552
rect 350 548 354 552
rect 798 658 802 662
rect 694 638 698 642
rect 782 638 786 642
rect 1094 748 1098 752
rect 986 703 990 707
rect 993 703 994 707
rect 994 703 997 707
rect 1350 1148 1354 1152
rect 1358 1148 1362 1152
rect 1038 668 1042 672
rect 1126 658 1130 662
rect 798 578 802 582
rect 902 558 906 562
rect 358 528 362 532
rect 462 528 466 532
rect 238 488 242 492
rect 374 478 378 482
rect 646 478 650 482
rect 430 468 434 472
rect 474 403 478 407
rect 481 403 482 407
rect 482 403 485 407
rect 390 318 394 322
rect 62 138 66 142
rect 118 128 122 132
rect 78 78 82 82
rect 318 258 322 262
rect 254 168 258 172
rect 262 138 266 142
rect 886 478 890 482
rect 830 448 834 452
rect 474 203 478 207
rect 481 203 482 207
rect 482 203 485 207
rect 454 168 458 172
rect 550 278 554 282
rect 534 148 538 152
rect 526 138 530 142
rect 510 68 514 72
rect 822 338 826 342
rect 606 198 610 202
rect 830 328 834 332
rect 798 268 802 272
rect 694 258 698 262
rect 758 128 762 132
rect 830 198 834 202
rect 830 158 834 162
rect 910 258 914 262
rect 926 268 930 272
rect 878 148 882 152
rect 862 138 866 142
rect 678 78 682 82
rect 774 68 778 72
rect 1230 558 1234 562
rect 986 503 990 507
rect 993 503 994 507
rect 994 503 997 507
rect 1046 488 1050 492
rect 1126 468 1130 472
rect 998 338 1002 342
rect 986 303 990 307
rect 993 303 994 307
rect 994 303 997 307
rect 1030 318 1034 322
rect 934 158 938 162
rect 1166 348 1170 352
rect 1246 358 1250 362
rect 1126 328 1130 332
rect 1270 448 1274 452
rect 1302 668 1306 672
rect 1350 668 1354 672
rect 1126 278 1130 282
rect 1046 148 1050 152
rect 1014 128 1018 132
rect 986 103 990 107
rect 993 103 994 107
rect 994 103 997 107
rect 1030 88 1034 92
rect 1190 258 1194 262
rect 1134 88 1138 92
rect 1030 68 1034 72
rect 1046 58 1050 62
rect 1110 58 1114 62
rect 1286 148 1290 152
rect 474 3 478 7
rect 481 3 482 7
rect 482 3 485 7
<< metal5 >>
rect 478 1403 481 1407
rect 478 1402 482 1403
rect 514 1368 934 1371
rect 618 1358 638 1361
rect 594 1348 886 1351
rect 554 1338 846 1341
rect 314 1328 766 1331
rect 990 1303 993 1307
rect 990 1302 994 1303
rect 650 1278 990 1281
rect 674 1268 1190 1271
rect 478 1203 481 1207
rect 478 1202 482 1203
rect 1074 1168 1118 1171
rect 602 1158 918 1161
rect 730 1148 1150 1151
rect 1354 1148 1358 1151
rect 626 1138 1094 1141
rect 290 1128 614 1131
rect 618 1128 1078 1131
rect 990 1103 993 1107
rect 990 1102 994 1103
rect 954 1068 1150 1071
rect 874 1008 966 1011
rect 478 1003 481 1007
rect 478 1002 482 1003
rect 1042 968 1158 971
rect 898 958 1094 961
rect 202 938 750 941
rect 674 928 1230 931
rect 990 903 993 907
rect 990 902 994 903
rect 874 878 1166 881
rect 210 868 910 871
rect 290 858 342 861
rect 754 858 1070 861
rect 274 848 694 851
rect 178 828 206 831
rect 478 803 481 807
rect 478 802 482 803
rect 18 798 182 801
rect 1034 748 1094 751
rect 874 738 942 741
rect 990 703 993 707
rect 990 702 994 703
rect 634 668 1038 671
rect 1306 668 1350 671
rect 802 658 1126 661
rect 698 638 782 641
rect 478 603 481 607
rect 478 602 482 603
rect 634 578 798 581
rect 298 558 334 561
rect 906 558 1230 561
rect 346 548 350 551
rect 362 528 462 531
rect 990 503 993 507
rect 990 502 994 503
rect 242 488 1046 491
rect 378 478 646 481
rect 650 478 886 481
rect 434 468 1126 471
rect 834 448 1270 451
rect 478 403 481 407
rect 478 402 482 403
rect 1246 351 1249 358
rect 1170 348 1249 351
rect 826 338 998 341
rect 834 328 1126 331
rect 394 318 1030 321
rect 990 303 993 307
rect 990 302 994 303
rect 554 278 1126 281
rect 802 268 926 271
rect 322 258 694 261
rect 914 258 1190 261
rect 478 203 481 207
rect 478 202 482 203
rect 610 198 830 201
rect 258 168 454 171
rect 834 158 934 161
rect 538 148 878 151
rect 1050 148 1286 151
rect 66 138 262 141
rect 530 138 862 141
rect 122 128 758 131
rect 762 128 1014 131
rect 990 103 993 107
rect 990 102 994 103
rect 1034 88 1134 91
rect 82 78 678 81
rect 514 68 774 71
rect 778 68 1030 71
rect 1050 58 1110 61
rect 478 3 481 7
rect 478 2 482 3
<< m6contact >>
rect 472 1407 478 1408
rect 482 1407 488 1408
rect 472 1403 474 1407
rect 474 1403 478 1407
rect 482 1403 485 1407
rect 485 1403 488 1407
rect 472 1402 478 1403
rect 482 1402 488 1403
rect 984 1307 990 1308
rect 994 1307 1000 1308
rect 984 1303 986 1307
rect 986 1303 990 1307
rect 994 1303 997 1307
rect 997 1303 1000 1307
rect 984 1302 990 1303
rect 994 1302 1000 1303
rect 472 1207 478 1208
rect 482 1207 488 1208
rect 472 1203 474 1207
rect 474 1203 478 1207
rect 482 1203 485 1207
rect 485 1203 488 1207
rect 472 1202 478 1203
rect 482 1202 488 1203
rect 984 1107 990 1108
rect 994 1107 1000 1108
rect 984 1103 986 1107
rect 986 1103 990 1107
rect 994 1103 997 1107
rect 997 1103 1000 1107
rect 984 1102 990 1103
rect 994 1102 1000 1103
rect 472 1007 478 1008
rect 482 1007 488 1008
rect 472 1003 474 1007
rect 474 1003 478 1007
rect 482 1003 485 1007
rect 485 1003 488 1007
rect 472 1002 478 1003
rect 482 1002 488 1003
rect 984 907 990 908
rect 994 907 1000 908
rect 984 903 986 907
rect 986 903 990 907
rect 994 903 997 907
rect 997 903 1000 907
rect 984 902 990 903
rect 994 902 1000 903
rect 472 807 478 808
rect 482 807 488 808
rect 472 803 474 807
rect 474 803 478 807
rect 482 803 485 807
rect 485 803 488 807
rect 472 802 478 803
rect 482 802 488 803
rect 984 707 990 708
rect 994 707 1000 708
rect 984 703 986 707
rect 986 703 990 707
rect 994 703 997 707
rect 997 703 1000 707
rect 984 702 990 703
rect 994 702 1000 703
rect 472 607 478 608
rect 482 607 488 608
rect 472 603 474 607
rect 474 603 478 607
rect 482 603 485 607
rect 485 603 488 607
rect 472 602 478 603
rect 482 602 488 603
rect 984 507 990 508
rect 994 507 1000 508
rect 984 503 986 507
rect 986 503 990 507
rect 994 503 997 507
rect 997 503 1000 507
rect 984 502 990 503
rect 994 502 1000 503
rect 472 407 478 408
rect 482 407 488 408
rect 472 403 474 407
rect 474 403 478 407
rect 482 403 485 407
rect 485 403 488 407
rect 472 402 478 403
rect 482 402 488 403
rect 984 307 990 308
rect 994 307 1000 308
rect 984 303 986 307
rect 986 303 990 307
rect 994 303 997 307
rect 997 303 1000 307
rect 984 302 990 303
rect 994 302 1000 303
rect 472 207 478 208
rect 482 207 488 208
rect 472 203 474 207
rect 474 203 478 207
rect 482 203 485 207
rect 485 203 488 207
rect 472 202 478 203
rect 482 202 488 203
rect 984 107 990 108
rect 994 107 1000 108
rect 984 103 986 107
rect 986 103 990 107
rect 994 103 997 107
rect 997 103 1000 107
rect 984 102 990 103
rect 994 102 1000 103
rect 472 7 478 8
rect 482 7 488 8
rect 472 3 474 7
rect 474 3 478 7
rect 482 3 485 7
rect 485 3 488 7
rect 472 2 478 3
rect 482 2 488 3
<< metal6 >>
rect 472 1408 488 1440
rect 478 1402 482 1408
rect 472 1208 488 1402
rect 478 1202 482 1208
rect 472 1008 488 1202
rect 478 1002 482 1008
rect 472 808 488 1002
rect 478 802 482 808
rect 472 608 488 802
rect 478 602 482 608
rect 472 408 488 602
rect 478 402 482 408
rect 472 208 488 402
rect 478 202 482 208
rect 472 8 488 202
rect 478 2 482 8
rect 472 -30 488 2
rect 984 1308 1000 1440
rect 990 1302 994 1308
rect 984 1108 1000 1302
rect 990 1102 994 1108
rect 984 908 1000 1102
rect 990 902 994 908
rect 984 708 1000 902
rect 990 702 994 708
rect 984 508 1000 702
rect 990 502 994 508
rect 984 308 1000 502
rect 990 302 994 308
rect 984 108 1000 302
rect 990 102 994 108
rect 984 -30 1000 102
use INVX1  _1059_
timestamp 1560018123
transform 1 0 4 0 1 1305
box -2 -3 18 103
use NAND2X1  _1060_
timestamp 1560018123
transform -1 0 44 0 1 1305
box -2 -3 26 103
use OR2X2  _1055_
timestamp 1560018123
transform 1 0 44 0 1 1305
box -2 -3 34 103
use NAND2X1  _1054_
timestamp 1560018123
transform -1 0 100 0 1 1305
box -2 -3 26 103
use NAND2X1  _1051_
timestamp 1560018123
transform 1 0 100 0 1 1305
box -2 -3 26 103
use INVX1  _1050_
timestamp 1560018123
transform -1 0 140 0 1 1305
box -2 -3 18 103
use INVX1  _1053_
timestamp 1560018123
transform -1 0 156 0 1 1305
box -2 -3 18 103
use INVX1  _1128_
timestamp 1560018123
transform -1 0 172 0 1 1305
box -2 -3 18 103
use NAND2X1  _1129_
timestamp 1560018123
transform -1 0 196 0 1 1305
box -2 -3 26 103
use OAI21X1  _1142_
timestamp 1560018123
transform -1 0 228 0 1 1305
box -2 -3 34 103
use INVX1  _1140_
timestamp 1560018123
transform -1 0 244 0 1 1305
box -2 -3 18 103
use NAND2X1  _1141_
timestamp 1560018123
transform -1 0 268 0 1 1305
box -2 -3 26 103
use NAND2X1  _1063_
timestamp 1560018123
transform 1 0 268 0 1 1305
box -2 -3 26 103
use INVX1  _1219_
timestamp 1560018123
transform 1 0 292 0 1 1305
box -2 -3 18 103
use NAND2X1  _1220_
timestamp 1560018123
transform -1 0 332 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert35
timestamp 1560018123
transform 1 0 332 0 1 1305
box -2 -3 26 103
use NAND2X1  _1229_
timestamp 1560018123
transform -1 0 380 0 1 1305
box -2 -3 26 103
use NAND2X1  _1307_
timestamp 1560018123
transform 1 0 380 0 1 1305
box -2 -3 26 103
use INVX1  _808_
timestamp 1560018123
transform 1 0 404 0 1 1305
box -2 -3 18 103
use OAI21X1  _810_
timestamp 1560018123
transform 1 0 420 0 1 1305
box -2 -3 34 103
use NAND2X1  _809_
timestamp 1560018123
transform -1 0 476 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_0_0
timestamp 1560018123
transform 1 0 476 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1560018123
transform 1 0 484 0 1 1305
box -2 -3 10 103
use NAND2X1  _797_
timestamp 1560018123
transform 1 0 492 0 1 1305
box -2 -3 26 103
use INVX1  _796_
timestamp 1560018123
transform -1 0 532 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_insert24
timestamp 1560018123
transform -1 0 556 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert21
timestamp 1560018123
transform 1 0 556 0 1 1305
box -2 -3 26 103
use OR2X2  _804_
timestamp 1560018123
transform 1 0 580 0 1 1305
box -2 -3 34 103
use NAND3X1  _807_
timestamp 1560018123
transform -1 0 644 0 1 1305
box -2 -3 34 103
use NAND2X1  _811_
timestamp 1560018123
transform -1 0 668 0 1 1305
box -2 -3 26 103
use NAND3X1  _812_
timestamp 1560018123
transform -1 0 700 0 1 1305
box -2 -3 34 103
use NAND2X1  _733_
timestamp 1560018123
transform 1 0 700 0 1 1305
box -2 -3 26 103
use OAI21X1  _732_
timestamp 1560018123
transform -1 0 756 0 1 1305
box -2 -3 34 103
use INVX1  _730_
timestamp 1560018123
transform -1 0 772 0 1 1305
box -2 -3 18 103
use NAND2X1  _731_
timestamp 1560018123
transform -1 0 796 0 1 1305
box -2 -3 26 103
use NAND2X1  _722_
timestamp 1560018123
transform 1 0 796 0 1 1305
box -2 -3 26 103
use INVX1  _721_
timestamp 1560018123
transform -1 0 836 0 1 1305
box -2 -3 18 103
use NAND2X1  _767_
timestamp 1560018123
transform 1 0 836 0 1 1305
box -2 -3 26 103
use INVX1  _766_
timestamp 1560018123
transform -1 0 876 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_insert23
timestamp 1560018123
transform -1 0 900 0 1 1305
box -2 -3 26 103
use INVX1  _679_
timestamp 1560018123
transform 1 0 900 0 1 1305
box -2 -3 18 103
use NAND2X1  _680_
timestamp 1560018123
transform -1 0 940 0 1 1305
box -2 -3 26 103
use INVX1  _974_
timestamp 1560018123
transform -1 0 956 0 1 1305
box -2 -3 18 103
use NAND2X1  _975_
timestamp 1560018123
transform -1 0 980 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_1_0
timestamp 1560018123
transform 1 0 980 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1560018123
transform 1 0 988 0 1 1305
box -2 -3 10 103
use OAI21X1  _976_
timestamp 1560018123
transform 1 0 996 0 1 1305
box -2 -3 34 103
use BUFX2  BUFX2_insert11
timestamp 1560018123
transform -1 0 1052 0 1 1305
box -2 -3 26 103
use OR2X2  _883_
timestamp 1560018123
transform 1 0 1052 0 1 1305
box -2 -3 34 103
use INVX1  _965_
timestamp 1560018123
transform 1 0 1084 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_insert14
timestamp 1560018123
transform 1 0 1100 0 1 1305
box -2 -3 26 103
use NAND2X1  _977_
timestamp 1560018123
transform -1 0 1148 0 1 1305
box -2 -3 26 103
use NAND2X1  _966_
timestamp 1560018123
transform -1 0 1172 0 1 1305
box -2 -3 26 103
use NAND2X1  _897_
timestamp 1560018123
transform 1 0 1172 0 1 1305
box -2 -3 26 103
use INVX1  _896_
timestamp 1560018123
transform 1 0 1196 0 1 1305
box -2 -3 18 103
use OAI21X1  _898_
timestamp 1560018123
transform -1 0 1244 0 1 1305
box -2 -3 34 103
use NAND2X1  _899_
timestamp 1560018123
transform -1 0 1268 0 1 1305
box -2 -3 26 103
use INVX1  _887_
timestamp 1560018123
transform 1 0 1268 0 1 1305
box -2 -3 18 103
use NAND2X1  _888_
timestamp 1560018123
transform -1 0 1308 0 1 1305
box -2 -3 26 103
use INVX1  _845_
timestamp 1560018123
transform 1 0 1308 0 1 1305
box -2 -3 18 103
use NAND2X1  _846_
timestamp 1560018123
transform -1 0 1348 0 1 1305
box -2 -3 26 103
use OR2X2  _844_
timestamp 1560018123
transform 1 0 1348 0 1 1305
box -2 -3 34 103
use NAND2X1  _927_
timestamp 1560018123
transform 1 0 1380 0 1 1305
box -2 -3 26 103
use NAND3X1  _929_
timestamp 1560018123
transform 1 0 1404 0 1 1305
box -2 -3 34 103
use INVX1  _926_
timestamp 1560018123
transform -1 0 1452 0 1 1305
box -2 -3 18 103
use FILL  FILL_14_1
timestamp 1560018123
transform 1 0 1452 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1560018123
transform 1 0 1460 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_3
timestamp 1560018123
transform 1 0 1468 0 1 1305
box -2 -3 10 103
use BUFX2  BUFX2_insert9
timestamp 1560018123
transform 1 0 4 0 -1 1305
box -2 -3 26 103
use OR2X2  _1058_
timestamp 1560018123
transform 1 0 28 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1061_
timestamp 1560018123
transform -1 0 92 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1056_
timestamp 1560018123
transform 1 0 92 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1052_
timestamp 1560018123
transform -1 0 156 0 -1 1305
box -2 -3 34 103
use OR2X2  _1049_
timestamp 1560018123
transform -1 0 188 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1130_
timestamp 1560018123
transform -1 0 220 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_insert6
timestamp 1560018123
transform -1 0 244 0 -1 1305
box -2 -3 26 103
use OR2X2  _1133_
timestamp 1560018123
transform -1 0 276 0 -1 1305
box -2 -3 34 103
use OAI21X1  _1064_
timestamp 1560018123
transform -1 0 308 0 -1 1305
box -2 -3 34 103
use OR2X2  _1127_
timestamp 1560018123
transform -1 0 340 0 -1 1305
box -2 -3 34 103
use INVX1  _1062_
timestamp 1560018123
transform -1 0 356 0 -1 1305
box -2 -3 18 103
use OAI21X1  _1230_
timestamp 1560018123
transform -1 0 388 0 -1 1305
box -2 -3 34 103
use INVX1  _1228_
timestamp 1560018123
transform -1 0 404 0 -1 1305
box -2 -3 18 103
use NAND3X1  _1222_
timestamp 1560018123
transform -1 0 436 0 -1 1305
box -2 -3 34 103
use OR2X2  _1221_
timestamp 1560018123
transform -1 0 468 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1560018123
transform -1 0 476 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1560018123
transform -1 0 484 0 -1 1305
box -2 -3 10 103
use OAI21X1  _1308_
timestamp 1560018123
transform -1 0 516 0 -1 1305
box -2 -3 34 103
use INVX1  _1306_
timestamp 1560018123
transform -1 0 532 0 -1 1305
box -2 -3 18 103
use INVX1  _1225_
timestamp 1560018123
transform -1 0 548 0 -1 1305
box -2 -3 18 103
use INVX1  _1294_
timestamp 1560018123
transform -1 0 564 0 -1 1305
box -2 -3 18 103
use OR2X2  _795_
timestamp 1560018123
transform 1 0 564 0 -1 1305
box -2 -3 34 103
use NAND3X1  _798_
timestamp 1560018123
transform -1 0 628 0 -1 1305
box -2 -3 34 103
use NAND2X1  _728_
timestamp 1560018123
transform 1 0 628 0 -1 1305
box -2 -3 26 103
use INVX1  _727_
timestamp 1560018123
transform -1 0 668 0 -1 1305
box -2 -3 18 103
use INVX1  _805_
timestamp 1560018123
transform 1 0 668 0 -1 1305
box -2 -3 18 103
use NAND2X1  _806_
timestamp 1560018123
transform -1 0 708 0 -1 1305
box -2 -3 26 103
use OR2X2  _726_
timestamp 1560018123
transform 1 0 708 0 -1 1305
box -2 -3 34 103
use NAND3X1  _729_
timestamp 1560018123
transform -1 0 772 0 -1 1305
box -2 -3 34 103
use NAND3X1  _734_
timestamp 1560018123
transform -1 0 804 0 -1 1305
box -2 -3 34 103
use NAND3X1  _813_
timestamp 1560018123
transform -1 0 836 0 -1 1305
box -2 -3 34 103
use NAND3X1  _724_
timestamp 1560018123
transform -1 0 868 0 -1 1305
box -2 -3 34 103
use OR2X2  _723_
timestamp 1560018123
transform -1 0 900 0 -1 1305
box -2 -3 34 103
use INVX1  _893_
timestamp 1560018123
transform 1 0 900 0 -1 1305
box -2 -3 18 103
use NAND3X1  _681_
timestamp 1560018123
transform -1 0 948 0 -1 1305
box -2 -3 34 103
use OR2X2  _678_
timestamp 1560018123
transform -1 0 980 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1560018123
transform 1 0 980 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1560018123
transform 1 0 988 0 -1 1305
box -2 -3 10 103
use INVX1  _962_
timestamp 1560018123
transform 1 0 996 0 -1 1305
box -2 -3 18 103
use NAND2X1  _963_
timestamp 1560018123
transform -1 0 1036 0 -1 1305
box -2 -3 26 103
use OR2X2  _892_
timestamp 1560018123
transform 1 0 1036 0 -1 1305
box -2 -3 34 103
use NAND2X1  _894_
timestamp 1560018123
transform 1 0 1068 0 -1 1305
box -2 -3 26 103
use OR2X2  _970_
timestamp 1560018123
transform 1 0 1092 0 -1 1305
box -2 -3 34 103
use NAND3X1  _895_
timestamp 1560018123
transform -1 0 1156 0 -1 1305
box -2 -3 34 103
use NAND3X1  _973_
timestamp 1560018123
transform 1 0 1156 0 -1 1305
box -2 -3 34 103
use INVX1  _971_
timestamp 1560018123
transform 1 0 1188 0 -1 1305
box -2 -3 18 103
use NAND2X1  _972_
timestamp 1560018123
transform -1 0 1228 0 -1 1305
box -2 -3 26 103
use NAND3X1  _978_
timestamp 1560018123
transform -1 0 1260 0 -1 1305
box -2 -3 34 103
use NAND3X1  _968_
timestamp 1560018123
transform -1 0 1292 0 -1 1305
box -2 -3 34 103
use OR2X2  _967_
timestamp 1560018123
transform -1 0 1324 0 -1 1305
box -2 -3 34 103
use NAND3X1  _900_
timestamp 1560018123
transform -1 0 1356 0 -1 1305
box -2 -3 34 103
use OR2X2  _889_
timestamp 1560018123
transform 1 0 1356 0 -1 1305
box -2 -3 34 103
use NAND3X1  _890_
timestamp 1560018123
transform 1 0 1388 0 -1 1305
box -2 -3 34 103
use NAND3X1  _847_
timestamp 1560018123
transform 1 0 1420 0 -1 1305
box -2 -3 34 103
use FILL  FILL_13_1
timestamp 1560018123
transform -1 0 1460 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1560018123
transform -1 0 1468 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_3
timestamp 1560018123
transform -1 0 1476 0 -1 1305
box -2 -3 10 103
use INVX4  _1009_
timestamp 1560018123
transform -1 0 28 0 1 1105
box -2 -3 26 103
use NAND2X1  _1065_
timestamp 1560018123
transform 1 0 28 0 1 1105
box -2 -3 26 103
use NAND3X1  _1134_
timestamp 1560018123
transform -1 0 84 0 1 1105
box -2 -3 34 103
use NAND3X1  _1057_
timestamp 1560018123
transform -1 0 116 0 1 1105
box -2 -3 34 103
use NAND3X1  _1135_
timestamp 1560018123
transform -1 0 148 0 1 1105
box -2 -3 34 103
use NAND2X1  _1132_
timestamp 1560018123
transform 1 0 148 0 1 1105
box -2 -3 26 103
use INVX1  _1131_
timestamp 1560018123
transform -1 0 188 0 1 1105
box -2 -3 18 103
use NAND2X1  _1143_
timestamp 1560018123
transform 1 0 188 0 1 1105
box -2 -3 26 103
use INVX1  _1297_
timestamp 1560018123
transform -1 0 228 0 1 1105
box -2 -3 18 103
use NAND2X1  _1298_
timestamp 1560018123
transform -1 0 252 0 1 1105
box -2 -3 26 103
use OR2X2  _1299_
timestamp 1560018123
transform 1 0 252 0 1 1105
box -2 -3 34 103
use INVX1  _1303_
timestamp 1560018123
transform 1 0 284 0 1 1105
box -2 -3 18 103
use NAND2X1  _1304_
timestamp 1560018123
transform -1 0 324 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert37
timestamp 1560018123
transform -1 0 348 0 1 1105
box -2 -3 26 103
use NAND2X1  _1231_
timestamp 1560018123
transform 1 0 348 0 1 1105
box -2 -3 26 103
use OR2X2  _1224_
timestamp 1560018123
transform 1 0 372 0 1 1105
box -2 -3 34 103
use NAND2X1  _1309_
timestamp 1560018123
transform 1 0 404 0 1 1105
box -2 -3 26 103
use NAND2X1  _1226_
timestamp 1560018123
transform 1 0 428 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert36
timestamp 1560018123
transform 1 0 452 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_0_0
timestamp 1560018123
transform -1 0 484 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1560018123
transform -1 0 492 0 1 1105
box -2 -3 10 103
use OR2X2  _1215_
timestamp 1560018123
transform -1 0 524 0 1 1105
box -2 -3 34 103
use NAND2X1  _1295_
timestamp 1560018123
transform 1 0 524 0 1 1105
box -2 -3 26 103
use INVX1  _1177_
timestamp 1560018123
transform 1 0 548 0 1 1105
box -2 -3 18 103
use NAND2X1  _1178_
timestamp 1560018123
transform -1 0 588 0 1 1105
box -2 -3 26 103
use OR2X2  _801_
timestamp 1560018123
transform 1 0 588 0 1 1105
box -2 -3 34 103
use INVX1  _799_
timestamp 1560018123
transform 1 0 620 0 1 1105
box -2 -3 18 103
use NAND2X1  _800_
timestamp 1560018123
transform -1 0 660 0 1 1105
box -2 -3 26 103
use NAND3X1  _802_
timestamp 1560018123
transform -1 0 692 0 1 1105
box -2 -3 34 103
use NAND3X1  _803_
timestamp 1560018123
transform -1 0 724 0 1 1105
box -2 -3 34 103
use INVX2  _676_
timestamp 1560018123
transform 1 0 724 0 1 1105
box -2 -3 18 103
use INVX1  _682_
timestamp 1560018123
transform 1 0 740 0 1 1105
box -2 -3 18 103
use NAND2X1  _683_
timestamp 1560018123
transform -1 0 780 0 1 1105
box -2 -3 26 103
use OR2X2  _684_
timestamp 1560018123
transform 1 0 780 0 1 1105
box -2 -3 34 103
use NAND3X1  _685_
timestamp 1560018123
transform -1 0 844 0 1 1105
box -2 -3 34 103
use NAND3X1  _725_
timestamp 1560018123
transform -1 0 876 0 1 1105
box -2 -3 34 103
use NAND3X1  _686_
timestamp 1560018123
transform 1 0 876 0 1 1105
box -2 -3 34 103
use OR2X2  _717_
timestamp 1560018123
transform 1 0 908 0 1 1105
box -2 -3 34 103
use NAND3X1  _720_
timestamp 1560018123
transform -1 0 972 0 1 1105
box -2 -3 34 103
use INVX1  _718_
timestamp 1560018123
transform -1 0 988 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_1_0
timestamp 1560018123
transform -1 0 996 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1560018123
transform -1 0 1004 0 1 1105
box -2 -3 10 103
use NAND2X1  _719_
timestamp 1560018123
transform -1 0 1028 0 1 1105
box -2 -3 26 103
use NAND2X1  _761_
timestamp 1560018123
transform 1 0 1028 0 1 1105
box -2 -3 26 103
use INVX1  _760_
timestamp 1560018123
transform -1 0 1068 0 1 1105
box -2 -3 18 103
use INVX1  _884_
timestamp 1560018123
transform 1 0 1068 0 1 1105
box -2 -3 18 103
use OR2X2  _961_
timestamp 1560018123
transform 1 0 1084 0 1 1105
box -2 -3 34 103
use NAND3X1  _964_
timestamp 1560018123
transform -1 0 1148 0 1 1105
box -2 -3 34 103
use INVX1  _932_
timestamp 1560018123
transform 1 0 1148 0 1 1105
box -2 -3 18 103
use NAND2X1  _933_
timestamp 1560018123
transform -1 0 1188 0 1 1105
box -2 -3 26 103
use NAND2X1  _885_
timestamp 1560018123
transform -1 0 1212 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert12
timestamp 1560018123
transform -1 0 1236 0 1 1105
box -2 -3 26 103
use NAND3X1  _886_
timestamp 1560018123
transform -1 0 1268 0 1 1105
box -2 -3 34 103
use NAND3X1  _969_
timestamp 1560018123
transform -1 0 1300 0 1 1105
box -2 -3 34 103
use NAND3X1  _979_
timestamp 1560018123
transform -1 0 1332 0 1 1105
box -2 -3 34 103
use NAND3X1  _901_
timestamp 1560018123
transform -1 0 1364 0 1 1105
box -2 -3 34 103
use INVX2  _842_
timestamp 1560018123
transform 1 0 1364 0 1 1105
box -2 -3 18 103
use NAND3X1  _891_
timestamp 1560018123
transform 1 0 1380 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert10
timestamp 1560018123
transform -1 0 1436 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert13
timestamp 1560018123
transform -1 0 1460 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1560018123
transform 1 0 1460 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1560018123
transform 1 0 1468 0 1 1105
box -2 -3 10 103
use INVX1  _1014_
timestamp 1560018123
transform 1 0 4 0 -1 1105
box -2 -3 18 103
use NAND2X1  _1015_
timestamp 1560018123
transform -1 0 44 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert5
timestamp 1560018123
transform -1 0 68 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1066_
timestamp 1560018123
transform -1 0 100 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1067_
timestamp 1560018123
transform -1 0 132 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1145_
timestamp 1560018123
transform 1 0 132 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1099_
timestamp 1560018123
transform 1 0 164 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1144_
timestamp 1560018123
transform 1 0 188 0 -1 1105
box -2 -3 34 103
use INVX1  _1098_
timestamp 1560018123
transform -1 0 236 0 -1 1105
box -2 -3 18 103
use NAND3X1  _1139_
timestamp 1560018123
transform 1 0 236 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1138_
timestamp 1560018123
transform 1 0 268 0 -1 1105
box -2 -3 26 103
use INVX1  _1137_
timestamp 1560018123
transform -1 0 308 0 -1 1105
box -2 -3 18 103
use OR2X2  _1136_
timestamp 1560018123
transform -1 0 340 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1300_
timestamp 1560018123
transform -1 0 372 0 -1 1105
box -2 -3 34 103
use OR2X2  _1302_
timestamp 1560018123
transform 1 0 372 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1305_
timestamp 1560018123
transform -1 0 436 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1227_
timestamp 1560018123
transform -1 0 468 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1560018123
transform 1 0 468 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1560018123
transform 1 0 476 0 -1 1105
box -2 -3 10 103
use NAND3X1  _1218_
timestamp 1560018123
transform 1 0 484 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1217_
timestamp 1560018123
transform 1 0 516 0 -1 1105
box -2 -3 26 103
use INVX1  _1011_
timestamp 1560018123
transform -1 0 556 0 -1 1105
box -2 -3 18 103
use INVX1  _1216_
timestamp 1560018123
transform -1 0 572 0 -1 1105
box -2 -3 18 103
use NAND3X1  _1296_
timestamp 1560018123
transform -1 0 604 0 -1 1105
box -2 -3 34 103
use OR2X2  _1293_
timestamp 1560018123
transform -1 0 636 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1265_
timestamp 1560018123
transform 1 0 636 0 -1 1105
box -2 -3 26 103
use INVX1  _1264_
timestamp 1560018123
transform -1 0 676 0 -1 1105
box -2 -3 18 103
use OR2X2  _1182_
timestamp 1560018123
transform 1 0 676 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1183_
timestamp 1560018123
transform 1 0 708 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1181_
timestamp 1560018123
transform 1 0 740 0 -1 1105
box -2 -3 26 103
use INVX1  _1180_
timestamp 1560018123
transform -1 0 780 0 -1 1105
box -2 -3 18 103
use INVX4  _677_
timestamp 1560018123
transform 1 0 780 0 -1 1105
box -2 -3 26 103
use NAND3X1  _735_
timestamp 1560018123
transform -1 0 836 0 -1 1105
box -2 -3 34 103
use NAND3X1  _768_
timestamp 1560018123
transform -1 0 868 0 -1 1105
box -2 -3 34 103
use NAND3X1  _773_
timestamp 1560018123
transform 1 0 868 0 -1 1105
box -2 -3 34 103
use NAND3X1  _696_
timestamp 1560018123
transform -1 0 932 0 -1 1105
box -2 -3 34 103
use OR2X2  _765_
timestamp 1560018123
transform -1 0 964 0 -1 1105
box -2 -3 34 103
use INVX1  _848_
timestamp 1560018123
transform 1 0 964 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_1_0
timestamp 1560018123
transform 1 0 980 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1560018123
transform 1 0 988 0 -1 1105
box -2 -3 10 103
use OR2X2  _762_
timestamp 1560018123
transform 1 0 996 0 -1 1105
box -2 -3 34 103
use NAND3X1  _763_
timestamp 1560018123
transform 1 0 1028 0 -1 1105
box -2 -3 34 103
use NAND2X1  _849_
timestamp 1560018123
transform -1 0 1084 0 -1 1105
box -2 -3 26 103
use OR2X2  _850_
timestamp 1560018123
transform 1 0 1084 0 -1 1105
box -2 -3 34 103
use NAND3X1  _851_
timestamp 1560018123
transform -1 0 1148 0 -1 1105
box -2 -3 34 103
use OR2X2  _931_
timestamp 1560018123
transform 1 0 1148 0 -1 1105
box -2 -3 34 103
use NAND3X1  _934_
timestamp 1560018123
transform -1 0 1212 0 -1 1105
box -2 -3 34 103
use INVX4  _843_
timestamp 1560018123
transform 1 0 1212 0 -1 1105
box -2 -3 26 103
use NAND3X1  _939_
timestamp 1560018123
transform -1 0 1268 0 -1 1105
box -2 -3 34 103
use NAND3X1  _852_
timestamp 1560018123
transform -1 0 1300 0 -1 1105
box -2 -3 34 103
use NAND3X1  _930_
timestamp 1560018123
transform 1 0 1300 0 -1 1105
box -2 -3 34 103
use NAND3X1  _925_
timestamp 1560018123
transform 1 0 1332 0 -1 1105
box -2 -3 34 103
use OR2X2  _922_
timestamp 1560018123
transform -1 0 1396 0 -1 1105
box -2 -3 34 103
use INVX1  _923_
timestamp 1560018123
transform 1 0 1396 0 -1 1105
box -2 -3 18 103
use NAND2X1  _924_
timestamp 1560018123
transform -1 0 1436 0 -1 1105
box -2 -3 26 103
use OR2X2  _928_
timestamp 1560018123
transform 1 0 1436 0 -1 1105
box -2 -3 34 103
use FILL  FILL_11_1
timestamp 1560018123
transform -1 0 1476 0 -1 1105
box -2 -3 10 103
use NAND3X1  _1017_
timestamp 1560018123
transform -1 0 36 0 1 905
box -2 -3 34 103
use OR2X2  _1016_
timestamp 1560018123
transform -1 0 68 0 1 905
box -2 -3 34 103
use NAND3X1  _1018_
timestamp 1560018123
transform -1 0 100 0 1 905
box -2 -3 34 103
use INVX2  _1008_
timestamp 1560018123
transform -1 0 116 0 1 905
box -2 -3 18 103
use OR2X2  _1097_
timestamp 1560018123
transform 1 0 116 0 1 905
box -2 -3 34 103
use NAND3X1  _1100_
timestamp 1560018123
transform -1 0 180 0 1 905
box -2 -3 34 103
use NAND3X1  _1105_
timestamp 1560018123
transform 1 0 180 0 1 905
box -2 -3 34 103
use NAND3X1  _1013_
timestamp 1560018123
transform 1 0 212 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_insert8
timestamp 1560018123
transform 1 0 244 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_insert7
timestamp 1560018123
transform 1 0 268 0 1 905
box -2 -3 26 103
use NAND2X1  _1090_
timestamp 1560018123
transform 1 0 292 0 1 905
box -2 -3 26 103
use NAND2X1  _1012_
timestamp 1560018123
transform -1 0 340 0 1 905
box -2 -3 26 103
use OR2X2  _1010_
timestamp 1560018123
transform -1 0 372 0 1 905
box -2 -3 34 103
use NAND2X1  _1021_
timestamp 1560018123
transform 1 0 372 0 1 905
box -2 -3 26 103
use INVX1  _1089_
timestamp 1560018123
transform -1 0 412 0 1 905
box -2 -3 18 103
use NAND3X1  _1310_
timestamp 1560018123
transform -1 0 444 0 1 905
box -2 -3 34 103
use NAND3X1  _1232_
timestamp 1560018123
transform -1 0 476 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1560018123
transform -1 0 484 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1560018123
transform -1 0 492 0 1 905
box -2 -3 10 103
use NAND3X1  _1223_
timestamp 1560018123
transform -1 0 524 0 1 905
box -2 -3 34 103
use NAND3X1  _1301_
timestamp 1560018123
transform -1 0 556 0 1 905
box -2 -3 34 103
use INVX1  _1020_
timestamp 1560018123
transform -1 0 572 0 1 905
box -2 -3 18 103
use OR2X2  _1176_
timestamp 1560018123
transform 1 0 572 0 1 905
box -2 -3 34 103
use NAND3X1  _1179_
timestamp 1560018123
transform 1 0 604 0 1 905
box -2 -3 34 103
use NAND3X1  _1184_
timestamp 1560018123
transform 1 0 636 0 1 905
box -2 -3 34 103
use NAND3X1  _1266_
timestamp 1560018123
transform -1 0 700 0 1 905
box -2 -3 34 103
use NAND2X1  _1256_
timestamp 1560018123
transform 1 0 700 0 1 905
box -2 -3 26 103
use INVX1  _1255_
timestamp 1560018123
transform -1 0 740 0 1 905
box -2 -3 18 103
use OR2X2  _1263_
timestamp 1560018123
transform -1 0 772 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_insert39
timestamp 1560018123
transform -1 0 796 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_insert38
timestamp 1560018123
transform 1 0 796 0 1 905
box -2 -3 26 103
use NAND3X1  _774_
timestamp 1560018123
transform -1 0 852 0 1 905
box -2 -3 34 103
use NAND3X1  _764_
timestamp 1560018123
transform 1 0 852 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_insert20
timestamp 1560018123
transform 1 0 884 0 1 905
box -2 -3 26 103
use NAND2X1  _758_
timestamp 1560018123
transform 1 0 908 0 1 905
box -2 -3 26 103
use INVX1  _757_
timestamp 1560018123
transform -1 0 948 0 1 905
box -2 -3 18 103
use NAND3X1  _759_
timestamp 1560018123
transform -1 0 980 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1560018123
transform -1 0 988 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1560018123
transform -1 0 996 0 1 905
box -2 -3 10 103
use OR2X2  _756_
timestamp 1560018123
transform -1 0 1028 0 1 905
box -2 -3 34 103
use NAND2X1  _772_
timestamp 1560018123
transform -1 0 1052 0 1 905
box -2 -3 26 103
use NAND3X1  _695_
timestamp 1560018123
transform 1 0 1052 0 1 905
box -2 -3 34 103
use NAND2X1  _694_
timestamp 1560018123
transform 1 0 1084 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_insert22
timestamp 1560018123
transform 1 0 1108 0 1 905
box -2 -3 26 103
use OAI21X1  _771_
timestamp 1560018123
transform -1 0 1164 0 1 905
box -2 -3 34 103
use INVX1  _769_
timestamp 1560018123
transform -1 0 1180 0 1 905
box -2 -3 18 103
use NAND3X1  _690_
timestamp 1560018123
transform 1 0 1180 0 1 905
box -2 -3 34 103
use OR2X2  _687_
timestamp 1560018123
transform -1 0 1244 0 1 905
box -2 -3 34 103
use OAI21X1  _693_
timestamp 1560018123
transform -1 0 1276 0 1 905
box -2 -3 34 103
use INVX1  _691_
timestamp 1560018123
transform -1 0 1292 0 1 905
box -2 -3 18 103
use NAND3X1  _940_
timestamp 1560018123
transform -1 0 1324 0 1 905
box -2 -3 34 103
use NAND3X1  _862_
timestamp 1560018123
transform 1 0 1324 0 1 905
box -2 -3 34 103
use NAND3X1  _861_
timestamp 1560018123
transform 1 0 1356 0 1 905
box -2 -3 34 103
use NAND2X1  _855_
timestamp 1560018123
transform 1 0 1388 0 1 905
box -2 -3 26 103
use INVX1  _854_
timestamp 1560018123
transform -1 0 1428 0 1 905
box -2 -3 18 103
use NAND3X1  _856_
timestamp 1560018123
transform 1 0 1428 0 1 905
box -2 -3 34 103
use FILL  FILL_10_1
timestamp 1560018123
transform 1 0 1460 0 1 905
box -2 -3 10 103
use FILL  FILL_10_2
timestamp 1560018123
transform 1 0 1468 0 1 905
box -2 -3 10 103
use BUFX2  _647_
timestamp 1560018123
transform -1 0 28 0 -1 905
box -2 -3 26 103
use BUFX2  _646_
timestamp 1560018123
transform -1 0 52 0 -1 905
box -2 -3 26 103
use INVX2  _986_
timestamp 1560018123
transform 1 0 52 0 -1 905
box -2 -3 18 103
use BUFX2  _650_
timestamp 1560018123
transform -1 0 92 0 -1 905
box -2 -3 26 103
use NAND3X1  _1028_
timestamp 1560018123
transform 1 0 92 0 -1 905
box -2 -3 34 103
use NAND3X1  _1106_
timestamp 1560018123
transform 1 0 124 0 -1 905
box -2 -3 34 103
use NAND3X1  _1027_
timestamp 1560018123
transform 1 0 156 0 -1 905
box -2 -3 34 103
use NAND2X1  _1026_
timestamp 1560018123
transform 1 0 188 0 -1 905
box -2 -3 26 103
use NAND3X1  _1096_
timestamp 1560018123
transform 1 0 212 0 -1 905
box -2 -3 34 103
use NAND2X1  _1104_
timestamp 1560018123
transform 1 0 244 0 -1 905
box -2 -3 26 103
use NAND3X1  _1091_
timestamp 1560018123
transform 1 0 268 0 -1 905
box -2 -3 34 103
use NAND3X1  _1022_
timestamp 1560018123
transform 1 0 300 0 -1 905
box -2 -3 34 103
use OR2X2  _1019_
timestamp 1560018123
transform -1 0 364 0 -1 905
box -2 -3 34 103
use OR2X2  _1088_
timestamp 1560018123
transform -1 0 396 0 -1 905
box -2 -3 34 103
use NAND3X1  _1095_
timestamp 1560018123
transform 1 0 396 0 -1 905
box -2 -3 34 103
use NAND3X1  _1311_
timestamp 1560018123
transform -1 0 460 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1560018123
transform -1 0 468 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1560018123
transform -1 0 476 0 -1 905
box -2 -3 10 103
use NAND3X1  _1233_
timestamp 1560018123
transform -1 0 508 0 -1 905
box -2 -3 34 103
use INVX2  _1174_
timestamp 1560018123
transform 1 0 508 0 -1 905
box -2 -3 18 103
use NAND2X1  _1187_
timestamp 1560018123
transform 1 0 524 0 -1 905
box -2 -3 26 103
use INVX1  _1186_
timestamp 1560018123
transform -1 0 564 0 -1 905
box -2 -3 18 103
use NAND3X1  _1188_
timestamp 1560018123
transform -1 0 596 0 -1 905
box -2 -3 34 103
use OR2X2  _1185_
timestamp 1560018123
transform -1 0 628 0 -1 905
box -2 -3 34 103
use OR2X2  _1254_
timestamp 1560018123
transform 1 0 628 0 -1 905
box -2 -3 34 103
use NAND3X1  _1271_
timestamp 1560018123
transform 1 0 660 0 -1 905
box -2 -3 34 103
use NAND3X1  _1257_
timestamp 1560018123
transform 1 0 692 0 -1 905
box -2 -3 34 103
use NAND2X1  _1270_
timestamp 1560018123
transform 1 0 724 0 -1 905
box -2 -3 26 103
use OR2X2  _1094_
timestamp 1560018123
transform -1 0 780 0 -1 905
box -2 -3 34 103
use NAND3X1  _1261_
timestamp 1560018123
transform 1 0 780 0 -1 905
box -2 -3 34 103
use OR2X2  _1260_
timestamp 1560018123
transform -1 0 844 0 -1 905
box -2 -3 34 103
use NAND2X1  _1259_
timestamp 1560018123
transform 1 0 844 0 -1 905
box -2 -3 26 103
use INVX1  _1258_
timestamp 1560018123
transform -1 0 884 0 -1 905
box -2 -3 18 103
use INVX2  _654_
timestamp 1560018123
transform -1 0 900 0 -1 905
box -2 -3 18 103
use NAND2X1  _1093_
timestamp 1560018123
transform 1 0 900 0 -1 905
box -2 -3 26 103
use INVX1  _1092_
timestamp 1560018123
transform -1 0 940 0 -1 905
box -2 -3 18 103
use OAI21X1  _1103_
timestamp 1560018123
transform -1 0 972 0 -1 905
box -2 -3 34 103
use NAND2X1  _1102_
timestamp 1560018123
transform 1 0 972 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1560018123
transform -1 0 1004 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1560018123
transform -1 0 1012 0 -1 905
box -2 -3 10 103
use OAI21X1  _1025_
timestamp 1560018123
transform -1 0 1044 0 -1 905
box -2 -3 34 103
use NAND2X1  _1024_
timestamp 1560018123
transform 1 0 1044 0 -1 905
box -2 -3 26 103
use INVX1  _1023_
timestamp 1560018123
transform -1 0 1084 0 -1 905
box -2 -3 18 103
use NAND2X1  _1268_
timestamp 1560018123
transform 1 0 1084 0 -1 905
box -2 -3 26 103
use OAI21X1  _1269_
timestamp 1560018123
transform -1 0 1140 0 -1 905
box -2 -3 34 103
use INVX1  _1267_
timestamp 1560018123
transform -1 0 1156 0 -1 905
box -2 -3 18 103
use INVX1  _1101_
timestamp 1560018123
transform -1 0 1172 0 -1 905
box -2 -3 18 103
use NAND2X1  _770_
timestamp 1560018123
transform -1 0 1196 0 -1 905
box -2 -3 26 103
use NAND2X1  _689_
timestamp 1560018123
transform 1 0 1196 0 -1 905
box -2 -3 26 103
use INVX1  _688_
timestamp 1560018123
transform -1 0 1236 0 -1 905
box -2 -3 18 103
use NAND2X1  _692_
timestamp 1560018123
transform 1 0 1236 0 -1 905
box -2 -3 26 103
use NAND2X1  _938_
timestamp 1560018123
transform 1 0 1260 0 -1 905
box -2 -3 26 103
use INVX2  _820_
timestamp 1560018123
transform 1 0 1284 0 -1 905
box -2 -3 18 103
use INVX1  _935_
timestamp 1560018123
transform 1 0 1300 0 -1 905
box -2 -3 18 103
use OAI21X1  _937_
timestamp 1560018123
transform 1 0 1316 0 -1 905
box -2 -3 34 103
use NAND2X1  _936_
timestamp 1560018123
transform 1 0 1348 0 -1 905
box -2 -3 26 103
use NAND2X1  _860_
timestamp 1560018123
transform 1 0 1372 0 -1 905
box -2 -3 26 103
use OAI21X1  _859_
timestamp 1560018123
transform -1 0 1428 0 -1 905
box -2 -3 34 103
use INVX1  _857_
timestamp 1560018123
transform -1 0 1444 0 -1 905
box -2 -3 18 103
use NAND2X1  _858_
timestamp 1560018123
transform 1 0 1444 0 -1 905
box -2 -3 26 103
use FILL  FILL_9_1
timestamp 1560018123
transform -1 0 1476 0 -1 905
box -2 -3 10 103
use BUFX2  _645_
timestamp 1560018123
transform -1 0 28 0 1 705
box -2 -3 26 103
use DFFPOSX1  _1147_
timestamp 1560018123
transform -1 0 124 0 1 705
box -2 -3 98 103
use AOI21X1  _1107_
timestamp 1560018123
transform 1 0 124 0 1 705
box -2 -3 34 103
use INVX2  _985_
timestamp 1560018123
transform -1 0 172 0 1 705
box -2 -3 18 103
use DFFPOSX1  _1149_
timestamp 1560018123
transform -1 0 268 0 1 705
box -2 -3 98 103
use BUFX2  _638_
timestamp 1560018123
transform -1 0 292 0 1 705
box -2 -3 26 103
use DFFPOSX1  _1314_
timestamp 1560018123
transform -1 0 388 0 1 705
box -2 -3 98 103
use INVX2  _1152_
timestamp 1560018123
transform 1 0 388 0 1 705
box -2 -3 18 103
use AOI21X1  _1312_
timestamp 1560018123
transform 1 0 404 0 1 705
box -2 -3 34 103
use INVX2  _1151_
timestamp 1560018123
transform 1 0 436 0 1 705
box -2 -3 18 103
use AOI21X1  _1234_
timestamp 1560018123
transform -1 0 484 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1560018123
transform -1 0 492 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1560018123
transform -1 0 500 0 1 705
box -2 -3 10 103
use DFFPOSX1  _816_
timestamp 1560018123
transform -1 0 596 0 1 705
box -2 -3 98 103
use INVX4  _1175_
timestamp 1560018123
transform 1 0 596 0 1 705
box -2 -3 26 103
use NAND3X1  _1194_
timestamp 1560018123
transform 1 0 620 0 1 705
box -2 -3 34 103
use NAND3X1  _1272_
timestamp 1560018123
transform 1 0 652 0 1 705
box -2 -3 34 103
use NAND3X1  _1193_
timestamp 1560018123
transform 1 0 684 0 1 705
box -2 -3 34 103
use NAND3X1  _1262_
timestamp 1560018123
transform 1 0 716 0 1 705
box -2 -3 34 103
use NAND2X1  _1192_
timestamp 1560018123
transform 1 0 748 0 1 705
box -2 -3 26 103
use INVX2  _653_
timestamp 1560018123
transform 1 0 772 0 1 705
box -2 -3 18 103
use AOI21X1  _736_
timestamp 1560018123
transform -1 0 820 0 1 705
box -2 -3 34 103
use AOI21X1  _775_
timestamp 1560018123
transform -1 0 852 0 1 705
box -2 -3 34 103
use AOI21X1  _814_
timestamp 1560018123
transform -1 0 884 0 1 705
box -2 -3 34 103
use AOI21X1  _697_
timestamp 1560018123
transform -1 0 916 0 1 705
box -2 -3 34 103
use DFFPOSX1  _818_
timestamp 1560018123
transform 1 0 916 0 1 705
box -2 -3 98 103
use FILL  FILL_7_1_0
timestamp 1560018123
transform -1 0 1020 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1560018123
transform -1 0 1028 0 1 705
box -2 -3 10 103
use OAI21X1  _1191_
timestamp 1560018123
transform -1 0 1060 0 1 705
box -2 -3 34 103
use NAND2X1  _1190_
timestamp 1560018123
transform -1 0 1084 0 1 705
box -2 -3 26 103
use INVX1  _1189_
timestamp 1560018123
transform -1 0 1100 0 1 705
box -2 -3 18 103
use BUFX2  _640_
timestamp 1560018123
transform 1 0 1100 0 1 705
box -2 -3 26 103
use INVX2  _819_
timestamp 1560018123
transform 1 0 1124 0 1 705
box -2 -3 18 103
use DFFPOSX1  _982_
timestamp 1560018123
transform 1 0 1140 0 1 705
box -2 -3 98 103
use BUFX2  _642_
timestamp 1560018123
transform 1 0 1236 0 1 705
box -2 -3 26 103
use AOI21X1  _902_
timestamp 1560018123
transform -1 0 1292 0 1 705
box -2 -3 34 103
use AOI21X1  _863_
timestamp 1560018123
transform -1 0 1324 0 1 705
box -2 -3 34 103
use DFFPOSX1  _981_
timestamp 1560018123
transform 1 0 1324 0 1 705
box -2 -3 98 103
use BUFX2  _641_
timestamp 1560018123
transform 1 0 1420 0 1 705
box -2 -3 26 103
use OR2X2  _853_
timestamp 1560018123
transform 1 0 1444 0 1 705
box -2 -3 34 103
use BUFX2  _648_
timestamp 1560018123
transform -1 0 28 0 -1 705
box -2 -3 26 103
use DFFPOSX1  _1150_
timestamp 1560018123
transform -1 0 124 0 -1 705
box -2 -3 98 103
use AOI21X1  _1029_
timestamp 1560018123
transform 1 0 124 0 -1 705
box -2 -3 34 103
use AOI21X1  _1146_
timestamp 1560018123
transform 1 0 156 0 -1 705
box -2 -3 34 103
use AOI21X1  _1068_
timestamp 1560018123
transform 1 0 188 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1148_
timestamp 1560018123
transform -1 0 316 0 -1 705
box -2 -3 98 103
use BUFX2  _652_
timestamp 1560018123
transform -1 0 340 0 -1 705
box -2 -3 26 103
use DFFPOSX1  _1316_
timestamp 1560018123
transform -1 0 436 0 -1 705
box -2 -3 98 103
use BUFX2  _639_
timestamp 1560018123
transform -1 0 460 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_0_0
timestamp 1560018123
transform -1 0 468 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1560018123
transform -1 0 476 0 -1 705
box -2 -3 10 103
use DFFPOSX1  _817_
timestamp 1560018123
transform -1 0 572 0 -1 705
box -2 -3 98 103
use AOI21X1  _1195_
timestamp 1560018123
transform 1 0 572 0 -1 705
box -2 -3 34 103
use AOI21X1  _1273_
timestamp 1560018123
transform -1 0 636 0 -1 705
box -2 -3 34 103
use INVX1  _747_
timestamp 1560018123
transform 1 0 636 0 -1 705
box -2 -3 18 103
use INVX1  _913_
timestamp 1560018123
transform 1 0 652 0 -1 705
box -2 -3 18 103
use NAND2X1  _914_
timestamp 1560018123
transform -1 0 692 0 -1 705
box -2 -3 26 103
use NAND2X1  _748_
timestamp 1560018123
transform -1 0 716 0 -1 705
box -2 -3 26 103
use OR2X2  _746_
timestamp 1560018123
transform 1 0 716 0 -1 705
box -2 -3 34 103
use NAND3X1  _749_
timestamp 1560018123
transform -1 0 780 0 -1 705
box -2 -3 34 103
use OR2X2  _912_
timestamp 1560018123
transform 1 0 780 0 -1 705
box -2 -3 34 103
use NAND3X1  _915_
timestamp 1560018123
transform -1 0 844 0 -1 705
box -2 -3 34 103
use BUFX2  BUFX2_insert34
timestamp 1560018123
transform -1 0 868 0 -1 705
box -2 -3 26 103
use NAND3X1  _755_
timestamp 1560018123
transform -1 0 900 0 -1 705
box -2 -3 34 103
use NAND3X1  _794_
timestamp 1560018123
transform 1 0 900 0 -1 705
box -2 -3 34 103
use NAND3X1  _675_
timestamp 1560018123
transform 1 0 932 0 -1 705
box -2 -3 34 103
use NAND3X1  _716_
timestamp 1560018123
transform 1 0 964 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1560018123
transform 1 0 996 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1560018123
transform 1 0 1004 0 -1 705
box -2 -3 10 103
use DFFPOSX1  _1315_
timestamp 1560018123
transform 1 0 1012 0 -1 705
box -2 -3 98 103
use DFFPOSX1  _1313_
timestamp 1560018123
transform 1 0 1108 0 -1 705
box -2 -3 98 103
use BUFX2  _651_
timestamp 1560018123
transform 1 0 1204 0 -1 705
box -2 -3 26 103
use NAND3X1  _960_
timestamp 1560018123
transform -1 0 1260 0 -1 705
box -2 -3 34 103
use AOI21X1  _980_
timestamp 1560018123
transform 1 0 1260 0 -1 705
box -2 -3 34 103
use AOI21X1  _941_
timestamp 1560018123
transform -1 0 1324 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _983_
timestamp 1560018123
transform 1 0 1324 0 -1 705
box -2 -3 98 103
use BUFX2  _649_
timestamp 1560018123
transform 1 0 1420 0 -1 705
box -2 -3 26 103
use BUFX2  _643_
timestamp 1560018123
transform 1 0 1444 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1560018123
transform -1 0 1476 0 -1 705
box -2 -3 10 103
use NAND2X1  _1122_
timestamp 1560018123
transform -1 0 28 0 1 505
box -2 -3 26 103
use OR2X2  _1117_
timestamp 1560018123
transform 1 0 28 0 1 505
box -2 -3 34 103
use INVX1  _1118_
timestamp 1560018123
transform 1 0 60 0 1 505
box -2 -3 18 103
use NAND2X1  _1119_
timestamp 1560018123
transform -1 0 100 0 1 505
box -2 -3 26 103
use NAND3X1  _1126_
timestamp 1560018123
transform 1 0 100 0 1 505
box -2 -3 34 103
use INVX1  _1079_
timestamp 1560018123
transform 1 0 132 0 1 505
box -2 -3 18 103
use NAND2X1  _1080_
timestamp 1560018123
transform -1 0 172 0 1 505
box -2 -3 26 103
use NAND2X1  _1113_
timestamp 1560018123
transform 1 0 172 0 1 505
box -2 -3 26 103
use INVX1  _1112_
timestamp 1560018123
transform -1 0 212 0 1 505
box -2 -3 18 103
use INVX1  _1278_
timestamp 1560018123
transform 1 0 212 0 1 505
box -2 -3 18 103
use NAND2X1  _1279_
timestamp 1560018123
transform -1 0 252 0 1 505
box -2 -3 26 103
use INVX1  _1284_
timestamp 1560018123
transform 1 0 252 0 1 505
box -2 -3 18 103
use NAND2X1  _1285_
timestamp 1560018123
transform -1 0 292 0 1 505
box -2 -3 26 103
use OR2X2  _1283_
timestamp 1560018123
transform 1 0 292 0 1 505
box -2 -3 34 103
use NAND3X1  _1286_
timestamp 1560018123
transform -1 0 356 0 1 505
box -2 -3 34 103
use NAND3X1  _1291_
timestamp 1560018123
transform -1 0 388 0 1 505
box -2 -3 34 103
use NAND3X1  _1292_
timestamp 1560018123
transform -1 0 420 0 1 505
box -2 -3 34 103
use NAND2X1  _1288_
timestamp 1560018123
transform -1 0 444 0 1 505
box -2 -3 26 103
use OR2X2  _1244_
timestamp 1560018123
transform 1 0 444 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1560018123
transform 1 0 476 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1560018123
transform 1 0 484 0 1 505
box -2 -3 10 103
use NAND3X1  _1247_
timestamp 1560018123
transform 1 0 492 0 1 505
box -2 -3 34 103
use INVX1  _1245_
timestamp 1560018123
transform 1 0 524 0 1 505
box -2 -3 18 103
use NAND2X1  _1246_
timestamp 1560018123
transform -1 0 564 0 1 505
box -2 -3 26 103
use INVX1  _786_
timestamp 1560018123
transform 1 0 564 0 1 505
box -2 -3 18 103
use INVX1  _952_
timestamp 1560018123
transform 1 0 580 0 1 505
box -2 -3 18 103
use NAND2X1  _953_
timestamp 1560018123
transform -1 0 620 0 1 505
box -2 -3 26 103
use NAND2X1  _787_
timestamp 1560018123
transform -1 0 644 0 1 505
box -2 -3 26 103
use NAND2X1  _956_
timestamp 1560018123
transform 1 0 644 0 1 505
box -2 -3 26 103
use NAND2X1  _790_
timestamp 1560018123
transform -1 0 692 0 1 505
box -2 -3 26 103
use OR2X2  _785_
timestamp 1560018123
transform 1 0 692 0 1 505
box -2 -3 34 103
use NAND3X1  _788_
timestamp 1560018123
transform -1 0 756 0 1 505
box -2 -3 34 103
use OR2X2  _951_
timestamp 1560018123
transform 1 0 756 0 1 505
box -2 -3 34 103
use NAND3X1  _954_
timestamp 1560018123
transform -1 0 820 0 1 505
box -2 -3 34 103
use NAND3X1  _754_
timestamp 1560018123
transform -1 0 852 0 1 505
box -2 -3 34 103
use NAND3X1  _793_
timestamp 1560018123
transform 1 0 852 0 1 505
box -2 -3 34 103
use INVX2  _655_
timestamp 1560018123
transform 1 0 884 0 1 505
box -2 -3 18 103
use NAND3X1  _784_
timestamp 1560018123
transform 1 0 900 0 1 505
box -2 -3 34 103
use NAND3X1  _779_
timestamp 1560018123
transform 1 0 932 0 1 505
box -2 -3 34 103
use OR2X2  _776_
timestamp 1560018123
transform -1 0 996 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1560018123
transform 1 0 996 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1560018123
transform 1 0 1004 0 1 505
box -2 -3 10 103
use NAND3X1  _715_
timestamp 1560018123
transform 1 0 1012 0 1 505
box -2 -3 34 103
use NAND3X1  _710_
timestamp 1560018123
transform 1 0 1044 0 1 505
box -2 -3 34 103
use OR2X2  _707_
timestamp 1560018123
transform -1 0 1108 0 1 505
box -2 -3 34 103
use DFFPOSX1  _815_
timestamp 1560018123
transform 1 0 1108 0 1 505
box -2 -3 98 103
use NAND3X1  _920_
timestamp 1560018123
transform -1 0 1236 0 1 505
box -2 -3 34 103
use NAND3X1  _959_
timestamp 1560018123
transform 1 0 1236 0 1 505
box -2 -3 34 103
use NAND3X1  _921_
timestamp 1560018123
transform -1 0 1300 0 1 505
box -2 -3 34 103
use NAND2X1  _875_
timestamp 1560018123
transform 1 0 1300 0 1 505
box -2 -3 26 103
use INVX1  _874_
timestamp 1560018123
transform -1 0 1340 0 1 505
box -2 -3 18 103
use DFFPOSX1  _984_
timestamp 1560018123
transform 1 0 1340 0 1 505
box -2 -3 98 103
use BUFX2  _637_
timestamp 1560018123
transform 1 0 1436 0 1 505
box -2 -3 26 103
use FILL  FILL_6_1
timestamp 1560018123
transform 1 0 1460 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1560018123
transform 1 0 1468 0 1 505
box -2 -3 10 103
use INVX1  _1121_
timestamp 1560018123
transform 1 0 4 0 -1 505
box -2 -3 18 103
use OAI21X1  _1123_
timestamp 1560018123
transform 1 0 20 0 -1 505
box -2 -3 34 103
use NAND3X1  _1120_
timestamp 1560018123
transform 1 0 52 0 -1 505
box -2 -3 34 103
use NAND2X1  _1124_
timestamp 1560018123
transform -1 0 108 0 -1 505
box -2 -3 26 103
use NAND3X1  _1125_
timestamp 1560018123
transform 1 0 108 0 -1 505
box -2 -3 34 103
use NAND3X1  _1081_
timestamp 1560018123
transform -1 0 172 0 -1 505
box -2 -3 34 103
use OR2X2  _1078_
timestamp 1560018123
transform -1 0 204 0 -1 505
box -2 -3 34 103
use BUFX2  BUFX2_insert16
timestamp 1560018123
transform -1 0 228 0 -1 505
box -2 -3 26 103
use NAND3X1  _1115_
timestamp 1560018123
transform 1 0 228 0 -1 505
box -2 -3 34 103
use OR2X2  _1114_
timestamp 1560018123
transform -1 0 292 0 -1 505
box -2 -3 34 103
use NAND3X1  _1042_
timestamp 1560018123
transform 1 0 292 0 -1 505
box -2 -3 34 103
use OR2X2  _1039_
timestamp 1560018123
transform -1 0 356 0 -1 505
box -2 -3 34 103
use NAND2X1  _1041_
timestamp 1560018123
transform 1 0 356 0 -1 505
box -2 -3 26 103
use OR2X2  _1280_
timestamp 1560018123
transform 1 0 380 0 -1 505
box -2 -3 34 103
use NAND3X1  _1281_
timestamp 1560018123
transform -1 0 444 0 -1 505
box -2 -3 34 103
use NAND3X1  _1282_
timestamp 1560018123
transform -1 0 476 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1560018123
transform -1 0 484 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1560018123
transform -1 0 492 0 -1 505
box -2 -3 10 103
use NAND3X1  _1252_
timestamp 1560018123
transform -1 0 524 0 -1 505
box -2 -3 34 103
use INVX1  _1287_
timestamp 1560018123
transform -1 0 540 0 -1 505
box -2 -3 18 103
use INVX1  _1040_
timestamp 1560018123
transform -1 0 556 0 -1 505
box -2 -3 18 103
use OAI21X1  _1289_
timestamp 1560018123
transform 1 0 556 0 -1 505
box -2 -3 34 103
use NAND2X1  _1290_
timestamp 1560018123
transform -1 0 612 0 -1 505
box -2 -3 26 103
use INVX4  _1154_
timestamp 1560018123
transform 1 0 612 0 -1 505
box -2 -3 26 103
use OR2X2  _1205_
timestamp 1560018123
transform 1 0 636 0 -1 505
box -2 -3 34 103
use NAND3X1  _1208_
timestamp 1560018123
transform 1 0 668 0 -1 505
box -2 -3 34 103
use NAND2X1  _1207_
timestamp 1560018123
transform 1 0 700 0 -1 505
box -2 -3 26 103
use INVX1  _1206_
timestamp 1560018123
transform -1 0 740 0 -1 505
box -2 -3 18 103
use INVX1  _955_
timestamp 1560018123
transform 1 0 740 0 -1 505
box -2 -3 18 103
use OAI21X1  _957_
timestamp 1560018123
transform -1 0 788 0 -1 505
box -2 -3 34 103
use INVX1  _789_
timestamp 1560018123
transform 1 0 788 0 -1 505
box -2 -3 18 103
use OAI21X1  _791_
timestamp 1560018123
transform 1 0 804 0 -1 505
box -2 -3 34 103
use OR2X2  _737_
timestamp 1560018123
transform 1 0 836 0 -1 505
box -2 -3 34 103
use NAND3X1  _740_
timestamp 1560018123
transform -1 0 900 0 -1 505
box -2 -3 34 103
use NAND3X1  _745_
timestamp 1560018123
transform 1 0 900 0 -1 505
box -2 -3 34 103
use NAND2X1  _792_
timestamp 1560018123
transform 1 0 932 0 -1 505
box -2 -3 26 103
use NAND2X1  _753_
timestamp 1560018123
transform -1 0 980 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_1_0
timestamp 1560018123
transform -1 0 988 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1560018123
transform -1 0 996 0 -1 505
box -2 -3 10 103
use BUFX2  BUFX2_insert31
timestamp 1560018123
transform -1 0 1020 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_insert33
timestamp 1560018123
transform 1 0 1020 0 -1 505
box -2 -3 26 103
use INVX1  _780_
timestamp 1560018123
transform 1 0 1044 0 -1 505
box -2 -3 18 103
use NAND2X1  _781_
timestamp 1560018123
transform -1 0 1084 0 -1 505
box -2 -3 26 103
use NAND3X1  _783_
timestamp 1560018123
transform -1 0 1116 0 -1 505
box -2 -3 34 103
use OR2X2  _782_
timestamp 1560018123
transform -1 0 1148 0 -1 505
box -2 -3 34 103
use NAND2X1  _714_
timestamp 1560018123
transform 1 0 1148 0 -1 505
box -2 -3 26 103
use INVX1  _708_
timestamp 1560018123
transform 1 0 1172 0 -1 505
box -2 -3 18 103
use NAND2X1  _709_
timestamp 1560018123
transform -1 0 1212 0 -1 505
box -2 -3 26 103
use NAND2X1  _778_
timestamp 1560018123
transform -1 0 1236 0 -1 505
box -2 -3 26 103
use NAND2X1  _919_
timestamp 1560018123
transform -1 0 1260 0 -1 505
box -2 -3 26 103
use NAND2X1  _958_
timestamp 1560018123
transform 1 0 1260 0 -1 505
box -2 -3 26 103
use INVX1  _946_
timestamp 1560018123
transform 1 0 1284 0 -1 505
box -2 -3 18 103
use OR2X2  _948_
timestamp 1560018123
transform 1 0 1300 0 -1 505
box -2 -3 34 103
use NAND3X1  _949_
timestamp 1560018123
transform 1 0 1332 0 -1 505
box -2 -3 34 103
use NAND2X1  _947_
timestamp 1560018123
transform -1 0 1388 0 -1 505
box -2 -3 26 103
use INVX4  _822_
timestamp 1560018123
transform 1 0 1388 0 -1 505
box -2 -3 26 103
use NAND3X1  _876_
timestamp 1560018123
transform 1 0 1412 0 -1 505
box -2 -3 34 103
use OR2X2  _873_
timestamp 1560018123
transform -1 0 1476 0 -1 505
box -2 -3 34 103
use NAND3X1  _1007_
timestamp 1560018123
transform -1 0 36 0 1 305
box -2 -3 34 103
use NAND3X1  _1047_
timestamp 1560018123
transform -1 0 68 0 1 305
box -2 -3 34 103
use NAND3X1  _1048_
timestamp 1560018123
transform -1 0 100 0 1 305
box -2 -3 34 103
use NAND3X1  _1087_
timestamp 1560018123
transform 1 0 100 0 1 305
box -2 -3 34 103
use NAND3X1  _1086_
timestamp 1560018123
transform 1 0 132 0 1 305
box -2 -3 34 103
use NAND3X1  _1116_
timestamp 1560018123
transform 1 0 164 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert19
timestamp 1560018123
transform 1 0 196 0 1 305
box -2 -3 26 103
use NAND3X1  _1111_
timestamp 1560018123
transform -1 0 252 0 1 305
box -2 -3 34 103
use NAND2X1  _1110_
timestamp 1560018123
transform 1 0 252 0 1 305
box -2 -3 26 103
use INVX1  _1109_
timestamp 1560018123
transform -1 0 292 0 1 305
box -2 -3 18 103
use OR2X2  _1108_
timestamp 1560018123
transform -1 0 324 0 1 305
box -2 -3 34 103
use INVX1  _1275_
timestamp 1560018123
transform 1 0 324 0 1 305
box -2 -3 18 103
use NAND2X1  _1276_
timestamp 1560018123
transform -1 0 364 0 1 305
box -2 -3 26 103
use NAND3X1  _1277_
timestamp 1560018123
transform -1 0 396 0 1 305
box -2 -3 34 103
use OR2X2  _1274_
timestamp 1560018123
transform -1 0 428 0 1 305
box -2 -3 34 103
use INVX1  _1248_
timestamp 1560018123
transform 1 0 428 0 1 305
box -2 -3 18 103
use OAI21X1  _1250_
timestamp 1560018123
transform 1 0 444 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1560018123
transform -1 0 484 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1560018123
transform -1 0 492 0 1 305
box -2 -3 10 103
use NAND2X1  _1251_
timestamp 1560018123
transform -1 0 516 0 1 305
box -2 -3 26 103
use NAND3X1  _1253_
timestamp 1560018123
transform -1 0 548 0 1 305
box -2 -3 34 103
use INVX2  _1153_
timestamp 1560018123
transform 1 0 548 0 1 305
box -2 -3 18 103
use NAND3X1  _1173_
timestamp 1560018123
transform 1 0 564 0 1 305
box -2 -3 34 103
use NAND3X1  _1214_
timestamp 1560018123
transform 1 0 596 0 1 305
box -2 -3 34 103
use NAND3X1  _1172_
timestamp 1560018123
transform 1 0 628 0 1 305
box -2 -3 34 103
use NAND3X1  _1213_
timestamp 1560018123
transform 1 0 660 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert0
timestamp 1560018123
transform -1 0 716 0 1 305
box -2 -3 26 103
use INVX1  _738_
timestamp 1560018123
transform 1 0 716 0 1 305
box -2 -3 18 103
use NAND2X1  _739_
timestamp 1560018123
transform -1 0 756 0 1 305
box -2 -3 26 103
use INVX1  _750_
timestamp 1560018123
transform 1 0 756 0 1 305
box -2 -3 18 103
use OAI21X1  _752_
timestamp 1560018123
transform 1 0 772 0 1 305
box -2 -3 34 103
use INVX1  _916_
timestamp 1560018123
transform 1 0 804 0 1 305
box -2 -3 18 103
use OR2X2  _743_
timestamp 1560018123
transform 1 0 820 0 1 305
box -2 -3 34 103
use NAND3X1  _744_
timestamp 1560018123
transform -1 0 884 0 1 305
box -2 -3 34 103
use NAND3X1  _660_
timestamp 1560018123
transform -1 0 916 0 1 305
box -2 -3 34 103
use INVX1  _824_
timestamp 1560018123
transform 1 0 916 0 1 305
box -2 -3 18 103
use NAND3X1  _665_
timestamp 1560018123
transform -1 0 964 0 1 305
box -2 -3 34 103
use NAND2X1  _825_
timestamp 1560018123
transform -1 0 988 0 1 305
box -2 -3 26 103
use FILL  FILL_3_1_0
timestamp 1560018123
transform 1 0 988 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1560018123
transform 1 0 996 0 1 305
box -2 -3 10 103
use OAI21X1  _918_
timestamp 1560018123
transform 1 0 1004 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert27
timestamp 1560018123
transform -1 0 1060 0 1 305
box -2 -3 26 103
use NAND3X1  _706_
timestamp 1560018123
transform 1 0 1060 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert25
timestamp 1560018123
transform -1 0 1116 0 1 305
box -2 -3 26 103
use OR2X2  _909_
timestamp 1560018123
transform 1 0 1116 0 1 305
box -2 -3 34 103
use OR2X2  _903_
timestamp 1560018123
transform 1 0 1148 0 1 305
box -2 -3 34 103
use NAND3X1  _906_
timestamp 1560018123
transform -1 0 1212 0 1 305
box -2 -3 34 103
use INVX1  _777_
timestamp 1560018123
transform -1 0 1228 0 1 305
box -2 -3 18 103
use NAND3X1  _910_
timestamp 1560018123
transform -1 0 1260 0 1 305
box -2 -3 34 103
use NAND3X1  _911_
timestamp 1560018123
transform -1 0 1292 0 1 305
box -2 -3 34 103
use NAND3X1  _882_
timestamp 1560018123
transform 1 0 1292 0 1 305
box -2 -3 34 103
use NAND3X1  _950_
timestamp 1560018123
transform 1 0 1324 0 1 305
box -2 -3 34 103
use NAND3X1  _945_
timestamp 1560018123
transform 1 0 1356 0 1 305
box -2 -3 34 103
use OR2X2  _942_
timestamp 1560018123
transform -1 0 1420 0 1 305
box -2 -3 34 103
use NAND3X1  _881_
timestamp 1560018123
transform 1 0 1420 0 1 305
box -2 -3 34 103
use NAND2X1  _944_
timestamp 1560018123
transform -1 0 1476 0 1 305
box -2 -3 26 103
use NAND3X1  _997_
timestamp 1560018123
transform -1 0 36 0 -1 305
box -2 -3 34 103
use INVX4  _988_
timestamp 1560018123
transform 1 0 36 0 -1 305
box -2 -3 26 103
use NAND3X1  _1006_
timestamp 1560018123
transform 1 0 60 0 -1 305
box -2 -3 34 103
use INVX2  _987_
timestamp 1560018123
transform 1 0 92 0 -1 305
box -2 -3 18 103
use NAND2X1  _1046_
timestamp 1560018123
transform 1 0 108 0 -1 305
box -2 -3 26 103
use NAND2X1  _1085_
timestamp 1560018123
transform 1 0 132 0 -1 305
box -2 -3 26 103
use NAND3X1  _1038_
timestamp 1560018123
transform 1 0 156 0 -1 305
box -2 -3 34 103
use NAND3X1  _1077_
timestamp 1560018123
transform 1 0 188 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert15
timestamp 1560018123
transform 1 0 220 0 -1 305
box -2 -3 26 103
use NAND3X1  _1033_
timestamp 1560018123
transform 1 0 244 0 -1 305
box -2 -3 34 103
use OR2X2  _1030_
timestamp 1560018123
transform -1 0 308 0 -1 305
box -2 -3 34 103
use NAND2X1  _1032_
timestamp 1560018123
transform -1 0 332 0 -1 305
box -2 -3 26 103
use OAI21X1  _1084_
timestamp 1560018123
transform -1 0 364 0 -1 305
box -2 -3 34 103
use INVX1  _1082_
timestamp 1560018123
transform -1 0 380 0 -1 305
box -2 -3 18 103
use NAND2X1  _1083_
timestamp 1560018123
transform 1 0 380 0 -1 305
box -2 -3 26 103
use INVX1  _1031_
timestamp 1560018123
transform -1 0 420 0 -1 305
box -2 -3 18 103
use BUFX2  BUFX2_insert3
timestamp 1560018123
transform -1 0 444 0 -1 305
box -2 -3 26 103
use NAND3X1  _1163_
timestamp 1560018123
transform -1 0 476 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1560018123
transform -1 0 484 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1560018123
transform -1 0 492 0 -1 305
box -2 -3 10 103
use NAND2X1  _1249_
timestamp 1560018123
transform -1 0 516 0 -1 305
box -2 -3 26 103
use NAND3X1  _1243_
timestamp 1560018123
transform -1 0 548 0 -1 305
box -2 -3 34 103
use INVX1  _1197_
timestamp 1560018123
transform 1 0 548 0 -1 305
box -2 -3 18 103
use NAND2X1  _1198_
timestamp 1560018123
transform 1 0 564 0 -1 305
box -2 -3 26 103
use NAND3X1  _1199_
timestamp 1560018123
transform -1 0 620 0 -1 305
box -2 -3 34 103
use NAND3X1  _1204_
timestamp 1560018123
transform 1 0 620 0 -1 305
box -2 -3 34 103
use NAND2X1  _1171_
timestamp 1560018123
transform 1 0 652 0 -1 305
box -2 -3 26 103
use OR2X2  _1196_
timestamp 1560018123
transform -1 0 708 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert4
timestamp 1560018123
transform -1 0 732 0 -1 305
box -2 -3 26 103
use NAND2X1  _1212_
timestamp 1560018123
transform 1 0 732 0 -1 305
box -2 -3 26 103
use INVX1  _904_
timestamp 1560018123
transform 1 0 756 0 -1 305
box -2 -3 18 103
use NAND2X1  _751_
timestamp 1560018123
transform 1 0 772 0 -1 305
box -2 -3 26 103
use OR2X2  _657_
timestamp 1560018123
transform 1 0 796 0 -1 305
box -2 -3 34 103
use NAND2X1  _742_
timestamp 1560018123
transform 1 0 828 0 -1 305
box -2 -3 26 103
use INVX1  _741_
timestamp 1560018123
transform -1 0 868 0 -1 305
box -2 -3 18 103
use INVX1  _658_
timestamp 1560018123
transform 1 0 868 0 -1 305
box -2 -3 18 103
use NAND2X1  _659_
timestamp 1560018123
transform -1 0 908 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert32
timestamp 1560018123
transform 1 0 908 0 -1 305
box -2 -3 26 103
use OR2X2  _823_
timestamp 1560018123
transform 1 0 932 0 -1 305
box -2 -3 34 103
use NAND3X1  _826_
timestamp 1560018123
transform -1 0 996 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1560018123
transform -1 0 1004 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1560018123
transform -1 0 1012 0 -1 305
box -2 -3 10 103
use NAND2X1  _917_
timestamp 1560018123
transform -1 0 1036 0 -1 305
box -2 -3 26 103
use OR2X2  _698_
timestamp 1560018123
transform 1 0 1036 0 -1 305
box -2 -3 34 103
use NAND3X1  _701_
timestamp 1560018123
transform 1 0 1068 0 -1 305
box -2 -3 34 103
use NAND2X1  _700_
timestamp 1560018123
transform 1 0 1100 0 -1 305
box -2 -3 26 103
use INVX1  _699_
timestamp 1560018123
transform -1 0 1140 0 -1 305
box -2 -3 18 103
use OR2X2  _864_
timestamp 1560018123
transform 1 0 1140 0 -1 305
box -2 -3 34 103
use INVX1  _907_
timestamp 1560018123
transform 1 0 1172 0 -1 305
box -2 -3 18 103
use NAND2X1  _905_
timestamp 1560018123
transform -1 0 1212 0 -1 305
box -2 -3 26 103
use NAND3X1  _867_
timestamp 1560018123
transform -1 0 1244 0 -1 305
box -2 -3 34 103
use NAND2X1  _908_
timestamp 1560018123
transform -1 0 1268 0 -1 305
box -2 -3 26 103
use NAND3X1  _831_
timestamp 1560018123
transform 1 0 1268 0 -1 305
box -2 -3 34 103
use NAND3X1  _841_
timestamp 1560018123
transform -1 0 1332 0 -1 305
box -2 -3 34 103
use INVX2  _821_
timestamp 1560018123
transform -1 0 1348 0 -1 305
box -2 -3 18 103
use NAND3X1  _872_
timestamp 1560018123
transform 1 0 1348 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert26
timestamp 1560018123
transform -1 0 1404 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert28
timestamp 1560018123
transform 1 0 1404 0 -1 305
box -2 -3 26 103
use NAND2X1  _880_
timestamp 1560018123
transform 1 0 1428 0 -1 305
box -2 -3 26 103
use FILL  FILL_3_1
timestamp 1560018123
transform -1 0 1460 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1560018123
transform -1 0 1468 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_3
timestamp 1560018123
transform -1 0 1476 0 -1 305
box -2 -3 10 103
use NAND3X1  _996_
timestamp 1560018123
transform 1 0 4 0 1 105
box -2 -3 34 103
use OR2X2  _995_
timestamp 1560018123
transform -1 0 68 0 1 105
box -2 -3 34 103
use NAND3X1  _1001_
timestamp 1560018123
transform 1 0 68 0 1 105
box -2 -3 34 103
use OR2X2  _998_
timestamp 1560018123
transform -1 0 132 0 1 105
box -2 -3 34 103
use NAND3X1  _992_
timestamp 1560018123
transform -1 0 164 0 1 105
box -2 -3 34 103
use OR2X2  _989_
timestamp 1560018123
transform -1 0 196 0 1 105
box -2 -3 34 103
use NAND3X1  _1076_
timestamp 1560018123
transform 1 0 196 0 1 105
box -2 -3 34 103
use OR2X2  _1075_
timestamp 1560018123
transform -1 0 260 0 1 105
box -2 -3 34 103
use NAND3X1  _1072_
timestamp 1560018123
transform 1 0 260 0 1 105
box -2 -3 34 103
use NAND2X1  _1071_
timestamp 1560018123
transform 1 0 292 0 1 105
box -2 -3 26 103
use INVX1  _1070_
timestamp 1560018123
transform -1 0 332 0 1 105
box -2 -3 18 103
use OR2X2  _1069_
timestamp 1560018123
transform -1 0 364 0 1 105
box -2 -3 34 103
use OAI21X1  _1045_
timestamp 1560018123
transform -1 0 396 0 1 105
box -2 -3 34 103
use NAND2X1  _1044_
timestamp 1560018123
transform 1 0 396 0 1 105
box -2 -3 26 103
use NAND3X1  _1162_
timestamp 1560018123
transform -1 0 452 0 1 105
box -2 -3 34 103
use NAND3X1  _1158_
timestamp 1560018123
transform 1 0 452 0 1 105
box -2 -3 34 103
use FILL  FILL_1_0_0
timestamp 1560018123
transform 1 0 484 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1560018123
transform 1 0 492 0 1 105
box -2 -3 10 103
use OR2X2  _1161_
timestamp 1560018123
transform 1 0 500 0 1 105
box -2 -3 34 103
use INVX1  _1043_
timestamp 1560018123
transform -1 0 548 0 1 105
box -2 -3 18 103
use NAND3X1  _1242_
timestamp 1560018123
transform 1 0 548 0 1 105
box -2 -3 34 103
use OR2X2  _1241_
timestamp 1560018123
transform -1 0 612 0 1 105
box -2 -3 34 103
use NAND3X1  _1238_
timestamp 1560018123
transform 1 0 612 0 1 105
box -2 -3 34 103
use INVX1  _1236_
timestamp 1560018123
transform 1 0 644 0 1 105
box -2 -3 18 103
use NAND2X1  _1237_
timestamp 1560018123
transform -1 0 684 0 1 105
box -2 -3 26 103
use OR2X2  _1164_
timestamp 1560018123
transform 1 0 684 0 1 105
box -2 -3 34 103
use NAND3X1  _1167_
timestamp 1560018123
transform 1 0 716 0 1 105
box -2 -3 34 103
use INVX1  _1165_
timestamp 1560018123
transform 1 0 748 0 1 105
box -2 -3 18 103
use NAND2X1  _1166_
timestamp 1560018123
transform -1 0 788 0 1 105
box -2 -3 26 103
use NAND3X1  _1203_
timestamp 1560018123
transform 1 0 788 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert1
timestamp 1560018123
transform 1 0 820 0 1 105
box -2 -3 26 103
use OR2X2  _1202_
timestamp 1560018123
transform -1 0 876 0 1 105
box -2 -3 34 103
use OAI21X1  _1211_
timestamp 1560018123
transform -1 0 908 0 1 105
box -2 -3 34 103
use INVX1  _1209_
timestamp 1560018123
transform -1 0 924 0 1 105
box -2 -3 18 103
use NAND3X1  _664_
timestamp 1560018123
transform -1 0 956 0 1 105
box -2 -3 34 103
use NAND3X1  _674_
timestamp 1560018123
transform -1 0 988 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1560018123
transform -1 0 996 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1560018123
transform -1 0 1004 0 1 105
box -2 -3 10 103
use OR2X2  _663_
timestamp 1560018123
transform -1 0 1036 0 1 105
box -2 -3 34 103
use NAND3X1  _669_
timestamp 1560018123
transform -1 0 1068 0 1 105
box -2 -3 34 103
use OR2X2  _666_
timestamp 1560018123
transform -1 0 1100 0 1 105
box -2 -3 34 103
use INVX4  _656_
timestamp 1560018123
transform 1 0 1100 0 1 105
box -2 -3 26 103
use NAND3X1  _705_
timestamp 1560018123
transform -1 0 1156 0 1 105
box -2 -3 34 103
use OR2X2  _704_
timestamp 1560018123
transform -1 0 1188 0 1 105
box -2 -3 34 103
use INVX1  _711_
timestamp 1560018123
transform 1 0 1188 0 1 105
box -2 -3 18 103
use OAI21X1  _713_
timestamp 1560018123
transform 1 0 1204 0 1 105
box -2 -3 34 103
use NAND2X1  _712_
timestamp 1560018123
transform 1 0 1236 0 1 105
box -2 -3 26 103
use NAND3X1  _830_
timestamp 1560018123
transform -1 0 1292 0 1 105
box -2 -3 34 103
use OR2X2  _829_
timestamp 1560018123
transform -1 0 1324 0 1 105
box -2 -3 34 103
use OR2X2  _870_
timestamp 1560018123
transform 1 0 1324 0 1 105
box -2 -3 34 103
use NAND3X1  _871_
timestamp 1560018123
transform 1 0 1356 0 1 105
box -2 -3 34 103
use NAND3X1  _835_
timestamp 1560018123
transform -1 0 1420 0 1 105
box -2 -3 34 103
use NAND3X1  _840_
timestamp 1560018123
transform 1 0 1420 0 1 105
box -2 -3 34 103
use FILL  FILL_2_1
timestamp 1560018123
transform 1 0 1452 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1560018123
transform 1 0 1460 0 1 105
box -2 -3 10 103
use FILL  FILL_2_3
timestamp 1560018123
transform 1 0 1468 0 1 105
box -2 -3 10 103
use INVX1  _993_
timestamp 1560018123
transform 1 0 4 0 -1 105
box -2 -3 18 103
use NAND2X1  _994_
timestamp 1560018123
transform -1 0 44 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert17
timestamp 1560018123
transform -1 0 68 0 -1 105
box -2 -3 26 103
use INVX1  _999_
timestamp 1560018123
transform 1 0 68 0 -1 105
box -2 -3 18 103
use NAND2X1  _1000_
timestamp 1560018123
transform -1 0 108 0 -1 105
box -2 -3 26 103
use NAND2X1  _1005_
timestamp 1560018123
transform 1 0 108 0 -1 105
box -2 -3 26 103
use NAND2X1  _991_
timestamp 1560018123
transform 1 0 132 0 -1 105
box -2 -3 26 103
use INVX1  _990_
timestamp 1560018123
transform -1 0 172 0 -1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert18
timestamp 1560018123
transform 1 0 172 0 -1 105
box -2 -3 26 103
use NAND2X1  _1074_
timestamp 1560018123
transform 1 0 196 0 -1 105
box -2 -3 26 103
use NAND3X1  _1037_
timestamp 1560018123
transform 1 0 220 0 -1 105
box -2 -3 34 103
use OR2X2  _1036_
timestamp 1560018123
transform -1 0 284 0 -1 105
box -2 -3 34 103
use NAND2X1  _1035_
timestamp 1560018123
transform 1 0 284 0 -1 105
box -2 -3 26 103
use INVX1  _1034_
timestamp 1560018123
transform -1 0 324 0 -1 105
box -2 -3 18 103
use OAI21X1  _1004_
timestamp 1560018123
transform -1 0 356 0 -1 105
box -2 -3 34 103
use NAND2X1  _1003_
timestamp 1560018123
transform 1 0 356 0 -1 105
box -2 -3 26 103
use INVX1  _1073_
timestamp 1560018123
transform -1 0 396 0 -1 105
box -2 -3 18 103
use INVX1  _1159_
timestamp 1560018123
transform 1 0 396 0 -1 105
box -2 -3 18 103
use NAND2X1  _1160_
timestamp 1560018123
transform -1 0 436 0 -1 105
box -2 -3 26 103
use OR2X2  _1155_
timestamp 1560018123
transform 1 0 436 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_0_0
timestamp 1560018123
transform 1 0 468 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1560018123
transform 1 0 476 0 -1 105
box -2 -3 10 103
use INVX1  _1156_
timestamp 1560018123
transform 1 0 484 0 -1 105
box -2 -3 18 103
use NAND2X1  _1157_
timestamp 1560018123
transform 1 0 500 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert2
timestamp 1560018123
transform 1 0 524 0 -1 105
box -2 -3 26 103
use NAND2X1  _1240_
timestamp 1560018123
transform 1 0 548 0 -1 105
box -2 -3 26 103
use INVX1  _1239_
timestamp 1560018123
transform 1 0 572 0 -1 105
box -2 -3 18 103
use OR2X2  _1235_
timestamp 1560018123
transform 1 0 588 0 -1 105
box -2 -3 34 103
use INVX1  _1002_
timestamp 1560018123
transform -1 0 636 0 -1 105
box -2 -3 18 103
use NAND2X1  _1169_
timestamp 1560018123
transform -1 0 660 0 -1 105
box -2 -3 26 103
use OAI21X1  _1170_
timestamp 1560018123
transform -1 0 692 0 -1 105
box -2 -3 34 103
use INVX1  _1168_
timestamp 1560018123
transform -1 0 708 0 -1 105
box -2 -3 18 103
use INVX1  _1200_
timestamp 1560018123
transform 1 0 708 0 -1 105
box -2 -3 18 103
use NAND2X1  _1201_
timestamp 1560018123
transform -1 0 748 0 -1 105
box -2 -3 26 103
use NAND2X1  _1210_
timestamp 1560018123
transform -1 0 772 0 -1 105
box -2 -3 26 103
use INVX1  _661_
timestamp 1560018123
transform 1 0 772 0 -1 105
box -2 -3 18 103
use NAND2X1  _662_
timestamp 1560018123
transform -1 0 812 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert30
timestamp 1560018123
transform 1 0 812 0 -1 105
box -2 -3 26 103
use INVX1  _670_
timestamp 1560018123
transform 1 0 836 0 -1 105
box -2 -3 18 103
use OAI21X1  _672_
timestamp 1560018123
transform 1 0 852 0 -1 105
box -2 -3 34 103
use NAND2X1  _671_
timestamp 1560018123
transform -1 0 908 0 -1 105
box -2 -3 26 103
use NAND2X1  _673_
timestamp 1560018123
transform -1 0 932 0 -1 105
box -2 -3 26 103
use NAND2X1  _668_
timestamp 1560018123
transform 1 0 932 0 -1 105
box -2 -3 26 103
use INVX1  _667_
timestamp 1560018123
transform -1 0 972 0 -1 105
box -2 -3 18 103
use NAND2X1  _703_
timestamp 1560018123
transform 1 0 972 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_1_0
timestamp 1560018123
transform -1 0 1004 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1560018123
transform -1 0 1012 0 -1 105
box -2 -3 10 103
use INVX1  _702_
timestamp 1560018123
transform -1 0 1028 0 -1 105
box -2 -3 18 103
use INVX1  _833_
timestamp 1560018123
transform 1 0 1028 0 -1 105
box -2 -3 18 103
use INVX1  _827_
timestamp 1560018123
transform 1 0 1044 0 -1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert29
timestamp 1560018123
transform 1 0 1060 0 -1 105
box -2 -3 26 103
use NAND2X1  _828_
timestamp 1560018123
transform -1 0 1108 0 -1 105
box -2 -3 26 103
use NAND2X1  _834_
timestamp 1560018123
transform -1 0 1132 0 -1 105
box -2 -3 26 103
use INVX1  _865_
timestamp 1560018123
transform -1 0 1148 0 -1 105
box -2 -3 18 103
use NAND2X1  _866_
timestamp 1560018123
transform -1 0 1172 0 -1 105
box -2 -3 26 103
use INVX1  _868_
timestamp 1560018123
transform 1 0 1172 0 -1 105
box -2 -3 18 103
use NAND2X1  _869_
timestamp 1560018123
transform 1 0 1188 0 -1 105
box -2 -3 26 103
use OR2X2  _832_
timestamp 1560018123
transform 1 0 1212 0 -1 105
box -2 -3 34 103
use NAND2X1  _878_
timestamp 1560018123
transform 1 0 1244 0 -1 105
box -2 -3 26 103
use INVX1  _836_
timestamp 1560018123
transform 1 0 1268 0 -1 105
box -2 -3 18 103
use OAI21X1  _838_
timestamp 1560018123
transform 1 0 1284 0 -1 105
box -2 -3 34 103
use NAND2X1  _837_
timestamp 1560018123
transform -1 0 1340 0 -1 105
box -2 -3 26 103
use NAND2X1  _839_
timestamp 1560018123
transform -1 0 1364 0 -1 105
box -2 -3 26 103
use OAI21X1  _879_
timestamp 1560018123
transform -1 0 1396 0 -1 105
box -2 -3 34 103
use INVX1  _877_
timestamp 1560018123
transform -1 0 1412 0 -1 105
box -2 -3 18 103
use BUFX2  _644_
timestamp 1560018123
transform -1 0 1436 0 -1 105
box -2 -3 26 103
use INVX1  _943_
timestamp 1560018123
transform -1 0 1452 0 -1 105
box -2 -3 18 103
use FILL  FILL_1_1
timestamp 1560018123
transform -1 0 1460 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1560018123
transform -1 0 1468 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_3
timestamp 1560018123
transform -1 0 1476 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 472 -30 488 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 984 -30 1000 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 718 -22 722 7 FreeSans 24 0 0 0 CLK
port 2 nsew
flabel metal3 s -26 608 -22 612 7 FreeSans 24 0 0 0 DATA_A[31]
port 3 nsew
flabel metal2 s 1022 -22 1026 -18 7 FreeSans 24 270 0 0 DATA_A[30]
port 4 nsew
flabel metal2 s 1254 -22 1258 -18 7 FreeSans 24 270 0 0 DATA_A[29]
port 5 nsew
flabel metal2 s 1318 -22 1322 -18 7 FreeSans 24 270 0 0 DATA_A[28]
port 6 nsew
flabel metal3 s -26 548 -22 552 7 FreeSans 24 0 0 0 DATA_A[27]
port 7 nsew
flabel metal2 s 598 -22 602 -18 7 FreeSans 24 270 0 0 DATA_A[26]
port 8 nsew
flabel metal2 s 1174 -22 1178 -18 7 FreeSans 24 270 0 0 DATA_A[25]
port 9 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 DATA_A[24]
port 10 nsew
flabel metal3 s -26 528 -22 532 7 FreeSans 24 0 0 0 DATA_A[23]
port 11 nsew
flabel metal3 s -26 588 -22 592 7 FreeSans 24 0 0 0 DATA_A[22]
port 12 nsew
flabel metal3 s 1502 528 1506 532 3 FreeSans 24 0 0 0 DATA_A[21]
port 13 nsew
flabel metal3 s -26 98 -22 102 7 FreeSans 24 0 0 0 DATA_A[20]
port 14 nsew
flabel metal3 s 1502 78 1506 82 3 FreeSans 24 0 0 0 DATA_A[19]
port 15 nsew
flabel metal2 s 662 -22 666 -18 7 FreeSans 24 270 0 0 DATA_A[18]
port 16 nsew
flabel metal2 s 1134 -22 1138 -18 7 FreeSans 24 270 0 0 DATA_A[17]
port 17 nsew
flabel metal2 s 158 -22 162 -18 7 FreeSans 24 270 0 0 DATA_A[16]
port 18 nsew
flabel metal3 s -26 488 -22 492 7 FreeSans 24 0 0 0 DATA_A[15]
port 19 nsew
flabel metal2 s 374 -22 378 -18 7 FreeSans 24 270 0 0 DATA_A[14]
port 20 nsew
flabel metal3 s 1502 148 1506 152 3 FreeSans 24 0 0 0 DATA_A[13]
port 21 nsew
flabel metal2 s 1270 -22 1274 -18 7 FreeSans 24 270 0 0 DATA_A[12]
port 22 nsew
flabel metal3 s 1502 448 1506 452 3 FreeSans 24 0 0 0 DATA_A[11]
port 23 nsew
flabel metal2 s 622 -22 626 -18 7 FreeSans 24 270 0 0 DATA_A[10]
port 24 nsew
flabel metal2 s 270 -22 274 -18 7 FreeSans 24 270 0 0 DATA_A[9]
port 25 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 DATA_A[8]
port 26 nsew
flabel metal3 s -26 568 -22 572 7 FreeSans 24 0 0 0 DATA_A[7]
port 27 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 DATA_A[6]
port 28 nsew
flabel metal3 s 1502 488 1506 492 3 FreeSans 24 0 0 0 DATA_A[5]
port 29 nsew
flabel metal2 s 1222 -22 1226 -18 7 FreeSans 24 270 0 0 DATA_A[4]
port 30 nsew
flabel metal3 s 1502 338 1506 342 3 FreeSans 24 0 0 0 DATA_A[3]
port 31 nsew
flabel metal2 s 638 -22 642 -18 7 FreeSans 24 270 0 0 DATA_A[2]
port 32 nsew
flabel metal2 s 1150 -22 1154 -18 7 FreeSans 24 270 0 0 DATA_A[1]
port 33 nsew
flabel metal2 s 446 -22 450 -18 7 FreeSans 24 270 0 0 DATA_A[0]
port 34 nsew
flabel metal2 s 958 1438 962 1442 3 FreeSans 24 90 0 0 DATA_B[31]
port 35 nsew
flabel metal3 s 1502 1258 1506 1262 3 FreeSans 24 0 0 0 DATA_B[30]
port 36 nsew
flabel metal2 s 1214 1438 1218 1442 3 FreeSans 24 90 0 0 DATA_B[29]
port 37 nsew
flabel metal3 s 1502 848 1506 852 3 FreeSans 24 0 0 0 DATA_B[28]
port 38 nsew
flabel metal2 s 1086 1438 1090 1442 3 FreeSans 24 90 0 0 DATA_B[27]
port 39 nsew
flabel metal3 s 1502 868 1506 872 3 FreeSans 24 0 0 0 DATA_B[26]
port 40 nsew
flabel metal2 s 1270 1438 1274 1442 3 FreeSans 24 90 0 0 DATA_B[25]
port 41 nsew
flabel metal3 s -26 1078 -22 1082 7 FreeSans 24 0 0 0 DATA_B[24]
port 42 nsew
flabel metal2 s 1198 1438 1202 1442 3 FreeSans 24 90 0 0 DATA_B[23]
port 43 nsew
flabel metal3 s 1502 998 1506 1002 3 FreeSans 24 0 0 0 DATA_B[22]
port 44 nsew
flabel metal3 s -26 1328 -22 1332 7 FreeSans 24 0 0 0 DATA_B[21]
port 45 nsew
flabel metal3 s 1502 968 1506 972 3 FreeSans 24 0 0 0 DATA_B[20]
port 46 nsew
flabel metal2 s 518 1438 522 1442 3 FreeSans 24 90 0 0 DATA_B[19]
port 47 nsew
flabel metal2 s 862 1438 866 1442 3 FreeSans 24 90 0 0 DATA_B[18]
port 48 nsew
flabel metal2 s 142 1438 146 1442 3 FreeSans 24 90 0 0 DATA_B[17]
port 49 nsew
flabel metal2 s 1318 1438 1322 1442 3 FreeSans 24 90 0 0 DATA_B[16]
port 50 nsew
flabel metal2 s 542 1438 546 1442 3 FreeSans 24 90 0 0 DATA_B[15]
port 51 nsew
flabel metal3 s 1502 1068 1506 1072 3 FreeSans 24 0 0 0 DATA_B[14]
port 52 nsew
flabel metal2 s 1182 1438 1186 1442 3 FreeSans 24 90 0 0 DATA_B[13]
port 53 nsew
flabel metal3 s 1502 948 1506 952 3 FreeSans 24 0 0 0 DATA_B[12]
port 54 nsew
flabel metal2 s 1302 1438 1306 1442 3 FreeSans 24 90 0 0 DATA_B[11]
port 55 nsew
flabel metal3 s 1502 888 1506 892 3 FreeSans 24 0 0 0 DATA_B[10]
port 56 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 90 0 0 DATA_B[9]
port 57 nsew
flabel metal3 s -26 958 -22 962 7 FreeSans 24 0 0 0 DATA_B[8]
port 58 nsew
flabel metal2 s 614 1438 618 1442 3 FreeSans 24 90 0 0 DATA_B[7]
port 59 nsew
flabel metal3 s 1502 1048 1506 1052 3 FreeSans 24 0 0 0 DATA_B[6]
port 60 nsew
flabel metal3 s -26 1268 -22 1272 7 FreeSans 24 0 0 0 DATA_B[5]
port 61 nsew
flabel metal3 s 1502 738 1506 742 3 FreeSans 24 0 0 0 DATA_B[4]
port 62 nsew
flabel metal2 s 590 1438 594 1442 3 FreeSans 24 90 0 0 DATA_B[3]
port 63 nsew
flabel metal3 s -26 938 -22 942 7 FreeSans 24 0 0 0 DATA_B[2]
port 64 nsew
flabel metal2 s 1062 1438 1066 1442 3 FreeSans 24 90 0 0 DATA_B[1]
port 65 nsew
flabel metal3 s 1502 1328 1506 1332 3 FreeSans 24 0 0 0 DATA_B[0]
port 66 nsew
flabel metal3 s -26 688 -22 692 7 FreeSans 24 0 0 0 NIBBLE_OUT[15]
port 67 nsew
flabel metal3 s 1502 688 1506 692 3 FreeSans 24 0 0 0 NIBBLE_OUT[14]
port 68 nsew
flabel metal3 s -26 848 -22 852 7 FreeSans 24 0 0 0 NIBBLE_OUT[13]
port 69 nsew
flabel metal3 s 1502 648 1506 652 3 FreeSans 24 0 0 0 NIBBLE_OUT[12]
port 70 nsew
flabel metal3 s -26 668 -22 672 7 FreeSans 24 0 0 0 NIBBLE_OUT[11]
port 71 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 NIBBLE_OUT[10]
port 72 nsew
flabel metal3 s -26 888 -22 892 7 FreeSans 24 0 0 0 NIBBLE_OUT[9]
port 73 nsew
flabel metal3 s -26 778 -22 782 7 FreeSans 24 0 0 0 NIBBLE_OUT[8]
port 74 nsew
flabel metal3 s 1502 48 1506 52 3 FreeSans 24 270 0 0 NIBBLE_OUT[7]
port 75 nsew
flabel metal3 s 1502 668 1506 672 3 FreeSans 24 0 0 0 NIBBLE_OUT[6]
port 76 nsew
flabel metal3 s 1502 798 1506 802 3 FreeSans 24 0 0 0 NIBBLE_OUT[5]
port 77 nsew
flabel metal3 s 1502 778 1506 782 3 FreeSans 24 0 0 0 NIBBLE_OUT[4]
port 78 nsew
flabel metal3 s 1502 758 1506 762 3 FreeSans 24 0 0 0 NIBBLE_OUT[3]
port 79 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 NIBBLE_OUT[2]
port 80 nsew
flabel metal3 s -26 798 -22 802 7 FreeSans 24 0 0 0 NIBBLE_OUT[1]
port 81 nsew
flabel metal3 s 1502 548 1506 552 3 FreeSans 24 0 0 0 NIBBLE_OUT[0]
port 82 nsew
flabel metal3 s -26 758 -22 762 7 FreeSans 24 0 0 0 RESET_L
port 83 nsew
flabel metal3 s -26 738 -22 742 7 FreeSans 24 0 0 0 SEL[3]
port 84 nsew
flabel metal3 s -26 978 -22 982 7 FreeSans 24 0 0 0 SEL[2]
port 85 nsew
flabel metal3 s 1502 1178 1506 1182 3 FreeSans 24 0 0 0 SEL[1]
port 86 nsew
flabel metal2 s 822 1438 826 1442 3 FreeSans 24 90 0 0 SEL[0]
port 87 nsew
flabel metal2 s 534 -22 538 -18 7 FreeSans 24 270 0 0 sel_A[11]
port 88 nsew
flabel metal2 s 558 -22 562 -18 7 FreeSans 24 270 0 0 sel_A[10]
port 89 nsew
flabel metal2 s 582 -22 586 -18 7 FreeSans 24 270 0 0 sel_A[9]
port 90 nsew
flabel metal2 s 86 -22 90 -18 7 FreeSans 24 270 0 0 sel_A[8]
port 91 nsew
flabel metal3 s -26 258 -22 262 7 FreeSans 24 0 0 0 sel_A[7]
port 92 nsew
flabel metal3 s -26 278 -22 282 7 FreeSans 24 0 0 0 sel_A[6]
port 93 nsew
flabel metal2 s 1054 -22 1058 -18 7 FreeSans 24 270 0 0 sel_A[5]
port 94 nsew
flabel metal2 s 1350 -22 1354 -18 7 FreeSans 24 270 0 0 sel_A[4]
port 95 nsew
flabel metal3 s 1502 358 1506 362 3 FreeSans 24 0 0 0 sel_A[3]
port 96 nsew
flabel metal2 s 910 -22 914 -18 7 FreeSans 24 270 0 0 sel_A[2]
port 97 nsew
flabel metal2 s 942 -22 946 -18 7 FreeSans 24 270 0 0 sel_A[1]
port 98 nsew
flabel metal2 s 1006 -22 1010 -18 7 FreeSans 24 270 0 0 sel_A[0]
port 99 nsew
flabel metal2 s 342 1438 346 1442 3 FreeSans 24 90 0 0 sel_B[11]
port 100 nsew
flabel metal2 s 438 1438 442 1442 3 FreeSans 24 90 0 0 sel_B[10]
port 101 nsew
flabel metal3 s -26 998 -22 1002 7 FreeSans 24 0 0 0 sel_B[9]
port 102 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 sel_B[8]
port 103 nsew
flabel metal3 s -26 1138 -22 1142 7 FreeSans 24 0 0 0 sel_B[7]
port 104 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 sel_B[6]
port 105 nsew
flabel metal2 s 1038 1438 1042 1442 3 FreeSans 24 90 0 0 sel_B[5]
port 106 nsew
flabel metal3 s 1502 1348 1506 1352 3 FreeSans 24 90 0 0 sel_B[4]
port 107 nsew
flabel metal3 s 1502 1158 1506 1162 3 FreeSans 24 0 0 0 sel_B[3]
port 108 nsew
flabel metal2 s 566 1438 570 1442 3 FreeSans 24 90 0 0 sel_B[2]
port 109 nsew
flabel metal2 s 654 1438 658 1442 3 FreeSans 24 90 0 0 sel_B[1]
port 110 nsew
flabel metal2 s 694 1438 698 1442 3 FreeSans 24 90 0 0 sel_B[0]
port 111 nsew
<< end >>
