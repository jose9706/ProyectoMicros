/* Verilog module written by DEF2Verilog (qflow) */
module nibble_top (
    input CLK,
    input [31:0] DATA_A,
    input [31:0] DATA_B,
    output [3:0] DATA_OUT,
    input RESET_L,
    input [11:0] SEL_A,
    input [3:0] SEL_AB,
    input [11:0] SEL_B
);

wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire [3:0] _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _773_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire [1:1] _638_ ;
wire _218_ ;
wire _391_ ;
wire SEL_B_5_bF$buf0 ;
wire SEL_B_5_bF$buf1 ;
wire SEL_B_5_bF$buf2 ;
wire SEL_B_5_bF$buf3 ;
wire SEL_B_5_bF$buf4 ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire _197_ ;
wire [3:0] SEL_AB ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [3:0] _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire _285_ ;
wire [3:0] _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _761_ ;
wire _341_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire SEL_B_11_bF$buf0 ;
wire SEL_B_11_bF$buf1 ;
wire SEL_B_11_bF$buf2 ;
wire SEL_B_11_bF$buf3 ;
wire SEL_B_11_bF$buf4 ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire CLK_bF$buf0 ;
wire CLK_bF$buf1 ;
wire CLK_bF$buf2 ;
wire CLK_bF$buf3 ;
wire CLK_bF$buf4 ;
wire CLK_bF$buf5 ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire [3:0] DATA_OUT ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire SEL_B_2_bF$buf0 ;
wire SEL_B_2_bF$buf1 ;
wire SEL_B_2_bF$buf2 ;
wire SEL_B_2_bF$buf3 ;
wire SEL_B_2_bF$buf4 ;
wire [3:0] \nibble_mayor.nibble_D  ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire [3:0] \nibble_mayor.nibble_A  ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire [3:0] _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire [3:0] _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire [3:0] _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _772_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire [3:0] _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire RESET_L_bF$buf0 ;
wire RESET_L_bF$buf1 ;
wire RESET_L_bF$buf2 ;
wire RESET_L_bF$buf3 ;
wire RESET_L_bF$buf4 ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire [3:0] _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire [3:0] \nibble_mayor.nibble_C  ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire RESET_L ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire CLK ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire [3:0] _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire [3:0] _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _771_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire SEL_A_8_bF$buf0 ;
wire SEL_A_8_bF$buf1 ;
wire SEL_A_8_bF$buf2 ;
wire SEL_A_8_bF$buf3 ;
wire SEL_A_8_bF$buf4 ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire [31:0] DATA_A ;
wire [31:0] DATA_B ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _765_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire gnd = 1'b0 ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire [3:0] _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _762_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire SEL_B_8_bF$buf0 ;
wire SEL_B_8_bF$buf1 ;
wire SEL_B_8_bF$buf2 ;
wire SEL_B_8_bF$buf3 ;
wire SEL_B_8_bF$buf4 ;
wire _474_ ;
wire _283_ ;
wire _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire SEL_A_11_bF$buf0 ;
wire SEL_A_11_bF$buf1 ;
wire SEL_A_11_bF$buf2 ;
wire SEL_A_11_bF$buf3 ;
wire SEL_A_11_bF$buf4 ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire [3:0] NIBBLE_MAYOR ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire SEL_A_2_bF$buf0 ;
wire SEL_A_2_bF$buf1 ;
wire SEL_A_2_bF$buf2 ;
wire SEL_A_2_bF$buf3 ;
wire SEL_A_2_bF$buf4 ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire vdd = 1'b1 ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _66_ ;
wire [15:0] NIBBLES ;
wire _615_ ;
wire [11:0] SEL_A ;
wire [11:0] SEL_B ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire [3:0] \nibble_mayor.nibble_B  ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire SEL_A_5_bF$buf0 ;
wire SEL_A_5_bF$buf1 ;
wire SEL_A_5_bF$buf2 ;
wire SEL_A_5_bF$buf3 ;
wire SEL_A_5_bF$buf4 ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

NAND2X1 _1257_ (
    .A(SEL_A[7]),
    .B(_433_),
    .Y(_434_)
);

INVX1 _800_ (
    .A(DATA_A[22]),
    .Y(_152_)
);

OAI21X1 _1486_ (
    .A(_762_),
    .B(_763_),
    .C(_765_),
    .Y(_766_)
);

NAND2X1 _1066_ (
    .A(SEL_B_5_bF$buf3),
    .B(_250_),
    .Y(_251_)
);

NAND3X1 _1295_ (
    .A(SEL_A[10]),
    .B(_625_),
    .C(_624_),
    .Y(_626_)
);

NAND2X1 _1389_ (
    .A(SEL_B_11_bF$buf2),
    .B(_559_),
    .Y(_560_)
);

FILL FILL_7_1 (
);

DFFPOSX1 _1601_ (
    .Q(NIBBLE_MAYOR[0]),
    .CLK(CLK_bF$buf4),
    .D(_639_[0])
);

INVX1 _932_ (
    .A(DATA_B[29]),
    .Y(_123_)
);

NAND2X1 _1198_ (
    .A(SEL_B[7]),
    .B(_376_),
    .Y(_377_)
);

NAND3X1 _1410_ (
    .A(_618_),
    .B(_577_),
    .C(_579_),
    .Y(_580_)
);

BUFX2 BUFX2_insert30 (
    .A(SEL_A[2]),
    .Y(SEL_A_2_bF$buf4)
);

BUFX2 BUFX2_insert31 (
    .A(SEL_A[2]),
    .Y(SEL_A_2_bF$buf3)
);

BUFX2 BUFX2_insert32 (
    .A(SEL_A[2]),
    .Y(SEL_A_2_bF$buf2)
);

BUFX2 BUFX2_insert33 (
    .A(SEL_A[2]),
    .Y(SEL_A_2_bF$buf1)
);

BUFX2 BUFX2_insert34 (
    .A(SEL_A[2]),
    .Y(SEL_A_2_bF$buf0)
);

BUFX2 BUFX2_insert35 (
    .A(SEL_A[11]),
    .Y(SEL_A_11_bF$buf4)
);

BUFX2 BUFX2_insert36 (
    .A(SEL_A[11]),
    .Y(SEL_A_11_bF$buf3)
);

BUFX2 BUFX2_insert37 (
    .A(SEL_A[11]),
    .Y(SEL_A_11_bF$buf2)
);

BUFX2 BUFX2_insert38 (
    .A(SEL_A[11]),
    .Y(SEL_A_11_bF$buf1)
);

BUFX2 BUFX2_insert39 (
    .A(SEL_A[11]),
    .Y(SEL_A_11_bF$buf0)
);

NAND2X1 _970_ (
    .A(SEL_A_5_bF$buf0),
    .B(DATA_A[30]),
    .Y(_315_)
);

OAI22X1 _1504_ (
    .A(_651_),
    .B(\nibble_mayor.nibble_A [3]),
    .C(\nibble_mayor.nibble_A [1]),
    .D(_652_),
    .Y(_653_)
);

INVX1 _835_ (
    .A(DATA_A[27]),
    .Y(_28_)
);

INVX1 _1313_ (
    .A(DATA_B[26]),
    .Y(_486_)
);

NAND2X1 _1542_ (
    .A(_659_),
    .B(_677_),
    .Y(_691_)
);

OR2X2 _1122_ (
    .A(SEL_A_8_bF$buf1),
    .B(DATA_A[2]),
    .Y(_460_)
);

NAND3X1 _873_ (
    .A(_141_),
    .B(_62_),
    .C(_64_),
    .Y(_65_)
);

INVX1 _929_ (
    .A(DATA_B[21]),
    .Y(_120_)
);

NAND3X1 _1351_ (
    .A(_481_),
    .B(_520_),
    .C(_522_),
    .Y(_523_)
);

OR2X2 _1407_ (
    .A(SEL_A_11_bF$buf1),
    .B(DATA_A[1]),
    .Y(_577_)
);

OAI21X1 _1580_ (
    .A(_701_),
    .B(_702_),
    .C(_706_),
    .Y(_729_)
);

NAND3X1 _1160_ (
    .A(SEL_B[6]),
    .B(_335_),
    .C(_339_),
    .Y(_340_)
);

NAND2X1 _1216_ (
    .A(SEL_A_8_bF$buf3),
    .B(DATA_A[28]),
    .Y(_394_)
);

NAND2X1 _967_ (
    .A(SEL_A_5_bF$buf0),
    .B(_311_),
    .Y(_312_)
);

AOI21X1 _1445_ (
    .A(_595_),
    .B(_614_),
    .C(_615_),
    .Y(_479_[1])
);

OR2X2 _1025_ (
    .A(SEL_B_5_bF$buf1),
    .B(DATA_B[3]),
    .Y(_211_)
);

AND2X2 _776_ (
    .A(RESET_L_bF$buf2),
    .B(NIBBLE_MAYOR[2]),
    .Y(_0_[2])
);

INVX1 _1254_ (
    .A(DATA_A[13]),
    .Y(_431_)
);

AND2X2 _1483_ (
    .A(\nibble_mayor.nibble_C [3]),
    .B(\nibble_mayor.nibble_D [3]),
    .Y(_763_)
);

NAND3X1 _1063_ (
    .A(SEL_B[3]),
    .B(_243_),
    .C(_247_),
    .Y(_248_)
);

FILL FILL_13_1_0 (
);

FILL FILL_13_1_1 (
);

NAND2X1 _1539_ (
    .A(_680_),
    .B(_687_),
    .Y(_688_)
);

INVX2 _1119_ (
    .A(SEL_AB[2]),
    .Y(_457_)
);

INVX1 _1292_ (
    .A(DATA_A[26]),
    .Y(_623_)
);

OR2X2 _1348_ (
    .A(SEL_B_11_bF$buf0),
    .B(DATA_B[7]),
    .Y(_520_)
);

INVX1 _1577_ (
    .A(_646_),
    .Y(_726_)
);

NAND2X1 _1157_ (
    .A(SEL_B_8_bF$buf4),
    .B(DATA_B[30]),
    .Y(_337_)
);

NAND3X1 _1386_ (
    .A(_616_),
    .B(_547_),
    .C(_556_),
    .Y(_557_)
);

INVX1 _1195_ (
    .A(DATA_B[11]),
    .Y(_374_)
);

FILL FILL_5_1_0 (
);

FILL FILL_5_1_1 (
);

INVX1 _1289_ (
    .A(DATA_A[18]),
    .Y(_620_)
);

FILL FILL_0_1_0 (
);

FILL FILL_0_1_1 (
);

NOR2X1 _1501_ (
    .A(\nibble_mayor.nibble_A [2]),
    .B(_649_),
    .Y(_650_)
);

INVX1 _832_ (
    .A(DATA_A[19]),
    .Y(_25_)
);

INVX1 _1098_ (
    .A(DATA_B[29]),
    .Y(_282_)
);

INVX1 _1310_ (
    .A(DATA_B[18]),
    .Y(_483_)
);

FILL FILL_15_0_0 (
);

FILL FILL_15_0_1 (
);

OR2X2 _870_ (
    .A(SEL_A_2_bF$buf3),
    .B(DATA_A[0]),
    .Y(_62_)
);

NAND3X1 _926_ (
    .A(SEL_A[0]),
    .B(_112_),
    .C(_116_),
    .Y(_117_)
);

FILL FILL_10_0_0 (
);

FILL FILL_10_0_1 (
);

NAND3X1 _1404_ (
    .A(_480_),
    .B(_570_),
    .C(_574_),
    .Y(_575_)
);

NAND2X1 _1213_ (
    .A(SEL_A_8_bF$buf4),
    .B(_390_),
    .Y(_391_)
);

NAND3X1 _964_ (
    .A(_299_),
    .B(_304_),
    .C(_308_),
    .Y(_309_)
);

NAND2X1 _1442_ (
    .A(SEL_B[10]),
    .B(_611_),
    .Y(_612_)
);

OR2X2 _1022_ (
    .A(SEL_B_5_bF$buf0),
    .B(DATA_B[15]),
    .Y(_208_)
);

NAND3X1 _829_ (
    .A(SEL_AB[0]),
    .B(_13_),
    .C(_22_),
    .Y(_23_)
);

INVX1 _1251_ (
    .A(DATA_A[21]),
    .Y(_428_)
);

INVX2 _1307_ (
    .A(SEL_B[9]),
    .Y(_480_)
);

NAND2X1 _1480_ (
    .A(_759_),
    .B(_754_),
    .Y(_760_)
);

NAND2X1 _1060_ (
    .A(SEL_B_5_bF$buf2),
    .B(_244_),
    .Y(_245_)
);

FILL FILL_7_0_0 (
);

FILL FILL_7_0_1 (
);

OAI21X1 _1536_ (
    .A(\nibble_mayor.nibble_C [3]),
    .B(_748_),
    .C(_766_),
    .Y(_685_)
);

DFFPOSX1 _1116_ (
    .Q(NIBBLES[6]),
    .CLK(CLK_bF$buf1),
    .D(_161_[2])
);

NAND3X1 _867_ (
    .A(_3_),
    .B(_55_),
    .C(_59_),
    .Y(_60_)
);

NAND2X1 _1345_ (
    .A(SEL_A[10]),
    .B(_516_),
    .Y(_517_)
);

FILL FILL_2_0_0 (
);

FILL FILL_2_0_1 (
);

OAI21X1 _1574_ (
    .A(_694_),
    .B(_695_),
    .C(_679_),
    .Y(_723_)
);

NAND2X1 _1154_ (
    .A(SEL_B_8_bF$buf0),
    .B(_333_),
    .Y(_334_)
);

OAI21X1 _1383_ (
    .A(_552_),
    .B(SEL_A_11_bF$buf2),
    .C(_553_),
    .Y(_554_)
);

INVX1 _1439_ (
    .A(DATA_B[9]),
    .Y(_609_)
);

NAND3X1 _1019_ (
    .A(_163_),
    .B(_202_),
    .C(_204_),
    .Y(_205_)
);

INVX1 _1192_ (
    .A(DATA_B[19]),
    .Y(_371_)
);

NAND3X1 _1248_ (
    .A(SEL_A[7]),
    .B(_424_),
    .C(_423_),
    .Y(_425_)
);

NAND2X1 _999_ (
    .A(SEL_A_5_bF$buf4),
    .B(_184_),
    .Y(_185_)
);

INVX2 _1477_ (
    .A(\nibble_mayor.nibble_C [0]),
    .Y(_757_)
);

NAND2X1 _1057_ (
    .A(SEL_B_5_bF$buf2),
    .B(_241_),
    .Y(_242_)
);

INVX2 _1286_ (
    .A(SEL_A[9]),
    .Y(_617_)
);

INVX1 _1095_ (
    .A(DATA_B[21]),
    .Y(_279_)
);

NAND2X1 _923_ (
    .A(SEL_A_2_bF$buf1),
    .B(DATA_A[29]),
    .Y(_114_)
);

NAND3X1 _1189_ (
    .A(SEL_B[7]),
    .B(_367_),
    .C(_366_),
    .Y(_368_)
);

NAND2X1 _1401_ (
    .A(SEL_B_11_bF$buf1),
    .B(DATA_B[24]),
    .Y(_572_)
);

NAND3X1 _1210_ (
    .A(_458_),
    .B(_383_),
    .C(_387_),
    .Y(_388_)
);

NAND2X1 _961_ (
    .A(SEL_A_5_bF$buf3),
    .B(_305_),
    .Y(_306_)
);

OAI21X1 _826_ (
    .A(_18_),
    .B(SEL_B_2_bF$buf0),
    .C(_19_),
    .Y(_20_)
);

NAND2X1 _1304_ (
    .A(SEL_A[10]),
    .B(_634_),
    .Y(_635_)
);

OAI22X1 _1533_ (
    .A(_763_),
    .B(_762_),
    .C(_681_),
    .D(_752_),
    .Y(_682_)
);

AOI21X1 _1113_ (
    .A(_277_),
    .B(_296_),
    .C(_297_),
    .Y(_161_[1])
);

FILL FILL_12_1 (
);

NAND2X1 _864_ (
    .A(SEL_B_2_bF$buf2),
    .B(DATA_B[27]),
    .Y(_57_)
);

INVX1 _1342_ (
    .A(DATA_A[15]),
    .Y(_514_)
);

AOI22X1 _1571_ (
    .A(_709_),
    .B(_703_),
    .C(_715_),
    .D(_719_),
    .Y(_720_)
);

NAND3X1 _1151_ (
    .A(_321_),
    .B(_326_),
    .C(_330_),
    .Y(_331_)
);

NAND2X1 _1207_ (
    .A(SEL_A_8_bF$buf1),
    .B(_384_),
    .Y(_385_)
);

NAND2X1 _958_ (
    .A(SEL_A_5_bF$buf2),
    .B(_302_),
    .Y(_303_)
);

NAND3X1 _1380_ (
    .A(_618_),
    .B(_548_),
    .C(_550_),
    .Y(_551_)
);

INVX1 _1436_ (
    .A(DATA_B[17]),
    .Y(_606_)
);

OR2X2 _1016_ (
    .A(SEL_B_5_bF$buf3),
    .B(DATA_B[7]),
    .Y(_202_)
);

INVX1 _1245_ (
    .A(DATA_A[25]),
    .Y(_422_)
);

AOI21X1 _996_ (
    .A(_319_),
    .B(_182_),
    .C(_297_),
    .Y(_161_[2])
);

AOI22X1 _1474_ (
    .A(_749_),
    .B(_750_),
    .C(_753_),
    .D(_751_),
    .Y(_754_)
);

NAND3X1 _1054_ (
    .A(_298_),
    .B(_229_),
    .C(_238_),
    .Y(_239_)
);

DFFPOSX1 _1283_ (
    .Q(NIBBLES[11]),
    .CLK(CLK_bF$buf2),
    .D(_320_[3])
);

INVX1 _1339_ (
    .A(DATA_A[23]),
    .Y(_511_)
);

FILL FILL_2_1 (
);

FILL FILL_2_2 (
);

NAND3X1 _1092_ (
    .A(SEL_A[3]),
    .B(_271_),
    .C(_275_),
    .Y(_276_)
);

NAND2X1 _1568_ (
    .A(_757_),
    .B(_687_),
    .Y(_717_)
);

NAND2X1 _1148_ (
    .A(SEL_B_8_bF$buf3),
    .B(_327_),
    .Y(_328_)
);

INVX1 _899_ (
    .A(DATA_B[16]),
    .Y(_91_)
);

OR2X2 _1377_ (
    .A(SEL_A_11_bF$buf3),
    .B(DATA_A[4]),
    .Y(_548_)
);

NAND2X1 _920_ (
    .A(SEL_A_2_bF$buf2),
    .B(_110_),
    .Y(_111_)
);

INVX1 _1186_ (
    .A(DATA_B[31]),
    .Y(_365_)
);

NAND3X1 _823_ (
    .A(_4_),
    .B(_14_),
    .C(_16_),
    .Y(_17_)
);

NAND2X1 _1089_ (
    .A(SEL_A_5_bF$buf1),
    .B(DATA_A[29]),
    .Y(_273_)
);

INVX1 _1301_ (
    .A(DATA_A[14]),
    .Y(_632_)
);

AOI21X1 _1530_ (
    .A(_678_),
    .B(_667_),
    .C(_746_),
    .Y(_679_)
);

NAND2X1 _1110_ (
    .A(SEL_B[4]),
    .B(_293_),
    .Y(_294_)
);

NAND2X1 _861_ (
    .A(SEL_B_2_bF$buf2),
    .B(_53_),
    .Y(_54_)
);

NAND3X1 _917_ (
    .A(_140_),
    .B(_103_),
    .C(_107_),
    .Y(_108_)
);

NAND2X1 _1204_ (
    .A(SEL_A_8_bF$buf3),
    .B(_381_),
    .Y(_382_)
);

INVX4 _955_ (
    .A(SEL_A[4]),
    .Y(_300_)
);

NAND3X1 _1433_ (
    .A(SEL_B[10]),
    .B(_602_),
    .C(_601_),
    .Y(_603_)
);

NAND2X1 _1013_ (
    .A(SEL_A[4]),
    .B(_198_),
    .Y(_199_)
);

INVX1 _1242_ (
    .A(DATA_A[17]),
    .Y(_419_)
);

NAND2X1 _993_ (
    .A(SEL_B[4]),
    .B(_179_),
    .Y(_180_)
);

NAND2X1 _1471_ (
    .A(\nibble_mayor.nibble_C [2]),
    .B(\nibble_mayor.nibble_D [2]),
    .Y(_751_)
);

OAI21X1 _1051_ (
    .A(_234_),
    .B(SEL_A_5_bF$buf1),
    .C(_235_),
    .Y(_236_)
);

OAI21X1 _1527_ (
    .A(_672_),
    .B(_674_),
    .C(_675_),
    .Y(_676_)
);

INVX1 _1107_ (
    .A(DATA_B[9]),
    .Y(_291_)
);

NAND3X1 _858_ (
    .A(SEL_B[0]),
    .B(_46_),
    .C(_50_),
    .Y(_51_)
);

DFFPOSX1 _1280_ (
    .Q(NIBBLES[8]),
    .CLK(CLK_bF$buf2),
    .D(_320_[0])
);

NAND3X1 _1336_ (
    .A(SEL_A[10]),
    .B(_507_),
    .C(_506_),
    .Y(_508_)
);

OAI21X1 _1565_ (
    .A(_687_),
    .B(\nibble_mayor.nibble_D [0]),
    .C(RESET_L_bF$buf2),
    .Y(_714_)
);

NAND2X1 _1145_ (
    .A(SEL_B_8_bF$buf3),
    .B(_324_),
    .Y(_325_)
);

NAND3X1 _896_ (
    .A(SEL_B[1]),
    .B(_87_),
    .C(_86_),
    .Y(_88_)
);

OR2X2 _1374_ (
    .A(SEL_A_11_bF$buf1),
    .B(DATA_A[8]),
    .Y(_545_)
);

INVX1 _1183_ (
    .A(DATA_B[23]),
    .Y(_362_)
);

NAND3X1 _1239_ (
    .A(SEL_AB[2]),
    .B(_407_),
    .C(_416_),
    .Y(_417_)
);

INVX1 _1468_ (
    .A(\nibble_mayor.nibble_D [3]),
    .Y(_748_)
);

NAND3X1 _1048_ (
    .A(_300_),
    .B(_230_),
    .C(_232_),
    .Y(_233_)
);

OR2X2 _799_ (
    .A(SEL_A_2_bF$buf1),
    .B(DATA_A[6]),
    .Y(_151_)
);

NAND3X1 _1277_ (
    .A(_321_),
    .B(_449_),
    .C(_453_),
    .Y(_454_)
);

OR2X2 _820_ (
    .A(SEL_B_2_bF$buf4),
    .B(DATA_B[6]),
    .Y(_14_)
);

NAND2X1 _1086_ (
    .A(SEL_A_5_bF$buf0),
    .B(_269_),
    .Y(_270_)
);

NAND2X1 _914_ (
    .A(SEL_A_2_bF$buf0),
    .B(_104_),
    .Y(_105_)
);

AOI21X1 _1201_ (
    .A(_360_),
    .B(_379_),
    .C(_456_),
    .Y(_320_[3])
);

INVX2 _952_ (
    .A(RESET_L_bF$buf3),
    .Y(_297_)
);

INVX1 _1430_ (
    .A(DATA_B[29]),
    .Y(_600_)
);

INVX1 _1010_ (
    .A(DATA_A[15]),
    .Y(_196_)
);

OR2X2 _817_ (
    .A(SEL_B_2_bF$buf1),
    .B(DATA_B[10]),
    .Y(_11_)
);

INVX1 _990_ (
    .A(DATA_B[14]),
    .Y(_177_)
);

INVX1 _1524_ (
    .A(\nibble_mayor.nibble_A [0]),
    .Y(_673_)
);

INVX1 _1104_ (
    .A(DATA_B[17]),
    .Y(_288_)
);

NAND2X1 _855_ (
    .A(SEL_B_2_bF$buf1),
    .B(_47_),
    .Y(_48_)
);

INVX1 _1333_ (
    .A(DATA_A[27]),
    .Y(_505_)
);

NOR2X1 _1562_ (
    .A(\nibble_mayor.nibble_A [0]),
    .B(_710_),
    .Y(_711_)
);

INVX4 _1142_ (
    .A(SEL_B[7]),
    .Y(_322_)
);

INVX1 _893_ (
    .A(DATA_B[28]),
    .Y(_85_)
);

DFFPOSX1 _1618_ (
    .Q(\nibble_mayor.nibble_D [1]),
    .CLK(CLK_bF$buf5),
    .D(_643_[1])
);

DFFPOSX1 _949_ (
    .Q(NIBBLES[1]),
    .CLK(CLK_bF$buf3),
    .D(_2_[1])
);

NAND3X1 _1371_ (
    .A(_618_),
    .B(_539_),
    .C(_541_),
    .Y(_542_)
);

INVX1 _1427_ (
    .A(DATA_B[21]),
    .Y(_597_)
);

INVX1 _1007_ (
    .A(DATA_A[23]),
    .Y(_193_)
);

NAND3X1 _1180_ (
    .A(SEL_A[6]),
    .B(_354_),
    .C(_358_),
    .Y(_359_)
);

OAI21X1 _1236_ (
    .A(_412_),
    .B(SEL_B_8_bF$buf1),
    .C(_413_),
    .Y(_414_)
);

INVX1 _987_ (
    .A(DATA_B[22]),
    .Y(_174_)
);

AND2X2 _1465_ (
    .A(RESET_L_bF$buf3),
    .B(NIBBLES[3]),
    .Y(_640_[3])
);

OR2X2 _1045_ (
    .A(SEL_A_5_bF$buf1),
    .B(DATA_A[4]),
    .Y(_230_)
);

OR2X2 _796_ (
    .A(SEL_A_2_bF$buf4),
    .B(DATA_A[10]),
    .Y(_148_)
);

NAND2X1 _1274_ (
    .A(SEL_B_8_bF$buf4),
    .B(DATA_B[25]),
    .Y(_451_)
);

NAND3X1 _1083_ (
    .A(_299_),
    .B(_262_),
    .C(_266_),
    .Y(_267_)
);

AOI21X1 _1559_ (
    .A(_755_),
    .B(_644_),
    .C(_746_),
    .Y(_708_)
);

NAND3X1 _1139_ (
    .A(SEL_A[6]),
    .B(_472_),
    .C(_476_),
    .Y(_477_)
);

OR2X2 _1368_ (
    .A(SEL_A_11_bF$buf1),
    .B(DATA_A[0]),
    .Y(_539_)
);

NAND2X1 _911_ (
    .A(SEL_A_2_bF$buf0),
    .B(_101_),
    .Y(_102_)
);

OAI21X1 _1597_ (
    .A(_638_[1]),
    .B(_700_),
    .C(_743_),
    .Y(_639_[1])
);

NAND2X1 _1177_ (
    .A(SEL_A_8_bF$buf2),
    .B(DATA_A[31]),
    .Y(_356_)
);

NAND3X1 _814_ (
    .A(_4_),
    .B(_5_),
    .C(_7_),
    .Y(_8_)
);

NAND2X1 _1521_ (
    .A(\nibble_mayor.nibble_B [1]),
    .B(_669_),
    .Y(_670_)
);

NAND3X1 _1101_ (
    .A(SEL_B[4]),
    .B(_284_),
    .C(_283_),
    .Y(_285_)
);

NAND2X1 _852_ (
    .A(SEL_B_2_bF$buf1),
    .B(_44_),
    .Y(_45_)
);

AOI21X1 _908_ (
    .A(_80_),
    .B(_99_),
    .C(_138_),
    .Y(_2_[0])
);

INVX1 _1330_ (
    .A(DATA_A[19]),
    .Y(_502_)
);

INVX1 _890_ (
    .A(DATA_B[20]),
    .Y(_82_)
);

DFFPOSX1 _1615_ (
    .Q(\nibble_mayor.nibble_C [2]),
    .CLK(CLK_bF$buf5),
    .D(_642_[2])
);

NAND3X1 _946_ (
    .A(SEL_AB[0]),
    .B(_127_),
    .C(_136_),
    .Y(_137_)
);

CLKBUF1 CLKBUF1_insert50 (
    .A(CLK),
    .Y(CLK_bF$buf0)
);

NAND3X1 _1424_ (
    .A(SEL_A[9]),
    .B(_589_),
    .C(_593_),
    .Y(_594_)
);

NAND3X1 _1004_ (
    .A(SEL_A[4]),
    .B(_189_),
    .C(_188_),
    .Y(_190_)
);

NAND3X1 _1233_ (
    .A(_322_),
    .B(_408_),
    .C(_410_),
    .Y(_411_)
);

NAND3X1 _984_ (
    .A(SEL_B[4]),
    .B(_170_),
    .C(_169_),
    .Y(_171_)
);

AND2X2 _1462_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLES[0]),
    .Y(_640_[0])
);

OR2X2 _1042_ (
    .A(SEL_A_5_bF$buf2),
    .B(DATA_A[8]),
    .Y(_227_)
);

NAND3X1 _793_ (
    .A(_141_),
    .B(_142_),
    .C(_144_),
    .Y(_145_)
);

NAND3X1 _1518_ (
    .A(\nibble_mayor.nibble_B [2]),
    .B(_666_),
    .C(_662_),
    .Y(_667_)
);

NAND3X1 _849_ (
    .A(_139_),
    .B(_32_),
    .C(_41_),
    .Y(_42_)
);

NAND2X1 _1271_ (
    .A(SEL_B_8_bF$buf3),
    .B(_447_),
    .Y(_448_)
);

NAND3X1 _1327_ (
    .A(SEL_AB[3]),
    .B(_490_),
    .C(_499_),
    .Y(_500_)
);

NAND2X1 _1080_ (
    .A(SEL_A_5_bF$buf3),
    .B(_263_),
    .Y(_264_)
);

NAND2X1 _1556_ (
    .A(\nibble_mayor.nibble_A [1]),
    .B(_677_),
    .Y(_705_)
);

NAND2X1 _1136_ (
    .A(SEL_A_8_bF$buf3),
    .B(DATA_A[30]),
    .Y(_474_)
);

NAND3X1 _887_ (
    .A(SEL_A[0]),
    .B(_74_),
    .C(_78_),
    .Y(_79_)
);

NAND3X1 _1365_ (
    .A(_480_),
    .B(_532_),
    .C(_536_),
    .Y(_537_)
);

OAI21X1 _1594_ (
    .A(_740_),
    .B(_733_),
    .C(_741_),
    .Y(_639_[0])
);

NAND2X1 _1174_ (
    .A(SEL_A_8_bF$buf1),
    .B(_352_),
    .Y(_353_)
);

AND2X2 _1459_ (
    .A(RESET_L_bF$buf3),
    .B(NIBBLES[5]),
    .Y(_641_[1])
);

NAND3X1 _1039_ (
    .A(_300_),
    .B(_221_),
    .C(_223_),
    .Y(_224_)
);

NAND3X1 _1268_ (
    .A(SEL_B[6]),
    .B(_440_),
    .C(_444_),
    .Y(_445_)
);

FILL FILL_12_1_0 (
);

FILL FILL_12_1_1 (
);

OR2X2 _811_ (
    .A(DATA_B[2]),
    .B(SEL_B_2_bF$buf3),
    .Y(_5_)
);

OAI21X1 _1497_ (
    .A(_645_),
    .B(_746_),
    .C(_646_),
    .Y(_639_[3])
);

NAND2X1 _1077_ (
    .A(SEL_A_5_bF$buf3),
    .B(_260_),
    .Y(_261_)
);

NAND2X1 _905_ (
    .A(SEL_B[1]),
    .B(_96_),
    .Y(_97_)
);

FILL FILL_9_1_0 (
);

FILL FILL_9_1_1 (
);

DFFPOSX1 _1612_ (
    .Q(\nibble_mayor.nibble_B [3]),
    .CLK(CLK_bF$buf4),
    .D(_641_[3])
);

OAI21X1 _943_ (
    .A(_132_),
    .B(SEL_B_2_bF$buf2),
    .C(_133_),
    .Y(_134_)
);

FILL FILL_4_1_0 (
);

FILL FILL_4_1_1 (
);

NAND2X1 _1421_ (
    .A(SEL_A_11_bF$buf3),
    .B(DATA_A[29]),
    .Y(_591_)
);

INVX1 _1001_ (
    .A(DATA_A[27]),
    .Y(_187_)
);

NAND3X1 _808_ (
    .A(_139_),
    .B(_150_),
    .C(_159_),
    .Y(_160_)
);

OR2X2 _1230_ (
    .A(SEL_B_8_bF$buf1),
    .B(DATA_B[0]),
    .Y(_408_)
);

INVX1 _981_ (
    .A(DATA_B[26]),
    .Y(_168_)
);

OR2X2 _790_ (
    .A(SEL_A_2_bF$buf4),
    .B(DATA_A[2]),
    .Y(_142_)
);

NOR2X1 _1515_ (
    .A(\nibble_mayor.nibble_B [3]),
    .B(_658_),
    .Y(_664_)
);

OAI21X1 _846_ (
    .A(_37_),
    .B(SEL_A_2_bF$buf3),
    .C(_38_),
    .Y(_39_)
);

FILL FILL_14_0_0 (
);

FILL FILL_14_0_1 (
);

OAI21X1 _1324_ (
    .A(_495_),
    .B(SEL_B_11_bF$buf4),
    .C(_496_),
    .Y(_497_)
);

OAI21X1 _1553_ (
    .A(_687_),
    .B(\nibble_mayor.nibble_D [1]),
    .C(RESET_L_bF$buf2),
    .Y(_702_)
);

NAND2X1 _1133_ (
    .A(SEL_A_8_bF$buf4),
    .B(_470_),
    .Y(_471_)
);

NAND2X1 _884_ (
    .A(SEL_A_2_bF$buf2),
    .B(DATA_A[28]),
    .Y(_76_)
);

FILL FILL_14_1 (
);

DFFPOSX1 _1609_ (
    .Q(\nibble_mayor.nibble_B [0]),
    .CLK(CLK_bF$buf3),
    .D(_641_[0])
);

NAND2X1 _1362_ (
    .A(SEL_B_11_bF$buf2),
    .B(DATA_B[27]),
    .Y(_534_)
);

NAND2X1 _1418_ (
    .A(SEL_A_11_bF$buf3),
    .B(_587_),
    .Y(_588_)
);

NAND2X1 _1591_ (
    .A(_736_),
    .B(_739_),
    .Y(_638_[1])
);

NAND3X1 _1171_ (
    .A(_458_),
    .B(_345_),
    .C(_349_),
    .Y(_350_)
);

OR2X2 _1227_ (
    .A(SEL_B_8_bF$buf0),
    .B(DATA_B[12]),
    .Y(_405_)
);

INVX1 _978_ (
    .A(DATA_B[18]),
    .Y(_165_)
);

AND2X2 _1456_ (
    .A(RESET_L_bF$buf0),
    .B(NIBBLES[10]),
    .Y(_642_[2])
);

OR2X2 _1036_ (
    .A(SEL_A_5_bF$buf2),
    .B(DATA_A[0]),
    .Y(_221_)
);

INVX2 _787_ (
    .A(SEL_AB[0]),
    .Y(_139_)
);

FILL FILL_6_0_0 (
);

FILL FILL_6_0_1 (
);

NAND2X1 _1265_ (
    .A(SEL_B_8_bF$buf2),
    .B(_441_),
    .Y(_442_)
);

AOI22X1 _1494_ (
    .A(_754_),
    .B(_773_),
    .C(_760_),
    .D(_767_),
    .Y(_644_)
);

AOI21X1 _1074_ (
    .A(_239_),
    .B(_258_),
    .C(_297_),
    .Y(_161_[0])
);

FILL FILL_1_0_0 (
);

FILL FILL_1_0_1 (
);

BUFX2 BUFX2_insert0 (
    .A(SEL_B[11]),
    .Y(SEL_B_11_bF$buf4)
);

BUFX2 BUFX2_insert1 (
    .A(SEL_B[11]),
    .Y(SEL_B_11_bF$buf3)
);

BUFX2 BUFX2_insert2 (
    .A(SEL_B[11]),
    .Y(SEL_B_11_bF$buf2)
);

BUFX2 BUFX2_insert3 (
    .A(SEL_B[11]),
    .Y(SEL_B_11_bF$buf1)
);

BUFX2 BUFX2_insert4 (
    .A(SEL_B[11]),
    .Y(SEL_B_11_bF$buf0)
);

BUFX2 BUFX2_insert5 (
    .A(SEL_B[8]),
    .Y(SEL_B_8_bF$buf4)
);

BUFX2 BUFX2_insert6 (
    .A(SEL_B[8]),
    .Y(SEL_B_8_bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .A(SEL_B[8]),
    .Y(SEL_B_8_bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .A(SEL_B[8]),
    .Y(SEL_B_8_bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .A(SEL_B[8]),
    .Y(SEL_B_8_bF$buf0)
);

NAND2X1 _1359_ (
    .A(SEL_B_11_bF$buf3),
    .B(_530_),
    .Y(_531_)
);

FILL FILL_4_1 (
);

FILL FILL_4_2 (
);

INVX1 _902_ (
    .A(DATA_B[8]),
    .Y(_94_)
);

NAND2X1 _1588_ (
    .A(_645_),
    .B(_726_),
    .Y(_737_)
);

NAND2X1 _1168_ (
    .A(SEL_A_8_bF$buf0),
    .B(_346_),
    .Y(_347_)
);

INVX1 _1397_ (
    .A(DATA_B[16]),
    .Y(_568_)
);

NAND3X1 _940_ (
    .A(_4_),
    .B(_128_),
    .C(_130_),
    .Y(_131_)
);

OAI21X1 _805_ (
    .A(_155_),
    .B(SEL_A_2_bF$buf1),
    .C(_156_),
    .Y(_157_)
);

AOI21X1 _1512_ (
    .A(_655_),
    .B(_657_),
    .C(_660_),
    .Y(_661_)
);

NAND3X1 _843_ (
    .A(_141_),
    .B(_33_),
    .C(_35_),
    .Y(_36_)
);

NAND3X1 _1321_ (
    .A(_481_),
    .B(_491_),
    .C(_493_),
    .Y(_494_)
);

NAND3X1 _1550_ (
    .A(_652_),
    .B(_666_),
    .C(_662_),
    .Y(_699_)
);

NAND3X1 _1130_ (
    .A(_458_),
    .B(_463_),
    .C(_467_),
    .Y(_468_)
);

NAND2X1 _881_ (
    .A(SEL_A_2_bF$buf2),
    .B(_72_),
    .Y(_73_)
);

DFFPOSX1 _1606_ (
    .Q(\nibble_mayor.nibble_A [1]),
    .CLK(CLK_bF$buf3),
    .D(_640_[1])
);

OR2X2 _937_ (
    .A(SEL_B_2_bF$buf3),
    .B(DATA_B[1]),
    .Y(_128_)
);

NAND3X1 _1415_ (
    .A(_617_),
    .B(_580_),
    .C(_584_),
    .Y(_585_)
);

NAND3X1 _1224_ (
    .A(_322_),
    .B(_399_),
    .C(_401_),
    .Y(_402_)
);

INVX2 _975_ (
    .A(SEL_B[3]),
    .Y(_162_)
);

AND2X2 _1453_ (
    .A(RESET_L_bF$buf0),
    .B(NIBBLES[15]),
    .Y(_643_[3])
);

NAND3X1 _1033_ (
    .A(_162_),
    .B(_214_),
    .C(_218_),
    .Y(_219_)
);

DFFPOSX1 _784_ (
    .Q(_1_[2]),
    .CLK(CLK_bF$buf4),
    .D(_0_[2])
);

INVX2 _1509_ (
    .A(\nibble_mayor.nibble_A [3]),
    .Y(_658_)
);

NAND2X1 _1262_ (
    .A(SEL_B_8_bF$buf4),
    .B(_438_),
    .Y(_439_)
);

OR2X2 _1318_ (
    .A(SEL_B_11_bF$buf3),
    .B(DATA_B[6]),
    .Y(_491_)
);

INVX1 _1491_ (
    .A(\nibble_mayor.nibble_D [0]),
    .Y(_771_)
);

NAND2X1 _1071_ (
    .A(SEL_B[4]),
    .B(_255_),
    .Y(_256_)
);

OAI21X1 _1547_ (
    .A(_694_),
    .B(_695_),
    .C(_693_),
    .Y(_696_)
);

NAND2X1 _1127_ (
    .A(SEL_A_8_bF$buf2),
    .B(_464_),
    .Y(_465_)
);

NAND3X1 _878_ (
    .A(_140_),
    .B(_65_),
    .C(_69_),
    .Y(_70_)
);

NAND3X1 _1356_ (
    .A(SEL_B[9]),
    .B(_523_),
    .C(_527_),
    .Y(_528_)
);

AOI22X1 _1585_ (
    .A(_716_),
    .B(_733_),
    .C(_709_),
    .D(_703_),
    .Y(_734_)
);

NAND2X1 _1165_ (
    .A(SEL_A_8_bF$buf2),
    .B(_343_),
    .Y(_344_)
);

NAND3X1 _1394_ (
    .A(SEL_B[10]),
    .B(_564_),
    .C(_563_),
    .Y(_565_)
);

NAND3X1 _1259_ (
    .A(_457_),
    .B(_426_),
    .C(_435_),
    .Y(_436_)
);

NAND3X1 _802_ (
    .A(_141_),
    .B(_151_),
    .C(_153_),
    .Y(_154_)
);

NAND2X1 _1488_ (
    .A(\nibble_mayor.nibble_C [1]),
    .B(\nibble_mayor.nibble_D [1]),
    .Y(_768_)
);

INVX1 _1068_ (
    .A(DATA_B[8]),
    .Y(_253_)
);

OR2X2 _1297_ (
    .A(SEL_A_11_bF$buf3),
    .B(DATA_A[6]),
    .Y(_628_)
);

OR2X2 _840_ (
    .A(SEL_A_2_bF$buf3),
    .B(DATA_A[7]),
    .Y(_33_)
);

DFFPOSX1 _1603_ (
    .Q(NIBBLE_MAYOR[2]),
    .CLK(CLK_bF$buf4),
    .D(_639_[2])
);

OR2X2 _934_ (
    .A(SEL_B_2_bF$buf0),
    .B(DATA_B[13]),
    .Y(_125_)
);

NAND2X1 _1412_ (
    .A(SEL_A_11_bF$buf0),
    .B(_581_),
    .Y(_582_)
);

OR2X2 _1221_ (
    .A(SEL_B_8_bF$buf0),
    .B(DATA_B[4]),
    .Y(_399_)
);

NAND2X1 _972_ (
    .A(SEL_A[4]),
    .B(_316_),
    .Y(_317_)
);

AND2X2 _1450_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLES[12]),
    .Y(_643_[0])
);

NAND2X1 _1030_ (
    .A(SEL_B_5_bF$buf1),
    .B(DATA_B[27]),
    .Y(_216_)
);

BUFX2 _781_ (
    .A(_1_[3]),
    .Y(DATA_OUT[3])
);

NAND2X1 _1506_ (
    .A(\nibble_mayor.nibble_A [1]),
    .B(_652_),
    .Y(_655_)
);

OR2X2 _837_ (
    .A(SEL_A_2_bF$buf0),
    .B(DATA_A[11]),
    .Y(_30_)
);

OR2X2 _1315_ (
    .A(SEL_B_11_bF$buf1),
    .B(DATA_B[10]),
    .Y(_488_)
);

NAND3X1 _1544_ (
    .A(RESET_L_bF$buf1),
    .B(_691_),
    .C(_692_),
    .Y(_693_)
);

NAND2X1 _1124_ (
    .A(SEL_A_8_bF$buf1),
    .B(_461_),
    .Y(_462_)
);

NAND2X1 _875_ (
    .A(SEL_A_2_bF$buf4),
    .B(_66_),
    .Y(_67_)
);

NAND2X1 _1353_ (
    .A(SEL_B_11_bF$buf1),
    .B(_524_),
    .Y(_525_)
);

NAND2X1 _1409_ (
    .A(SEL_A_11_bF$buf1),
    .B(_578_),
    .Y(_579_)
);

AOI21X1 _1582_ (
    .A(_729_),
    .B(_730_),
    .C(_728_),
    .Y(_731_)
);

AOI21X1 _1162_ (
    .A(_478_),
    .B(_341_),
    .C(_456_),
    .Y(_320_[2])
);

NAND2X1 _1218_ (
    .A(SEL_A[7]),
    .B(_395_),
    .Y(_396_)
);

INVX1 _969_ (
    .A(DATA_A[14]),
    .Y(_314_)
);

INVX1 _1391_ (
    .A(DATA_B[28]),
    .Y(_562_)
);

DFFPOSX1 _1447_ (
    .Q(NIBBLES[13]),
    .CLK(CLK_bF$buf3),
    .D(_479_[1])
);

NAND2X1 _1027_ (
    .A(SEL_B_5_bF$buf2),
    .B(_212_),
    .Y(_213_)
);

BUFX2 _778_ (
    .A(_1_[0]),
    .Y(DATA_OUT[0])
);

OAI21X1 _1256_ (
    .A(_431_),
    .B(SEL_A_8_bF$buf3),
    .C(_432_),
    .Y(_433_)
);

NOR2X1 _1485_ (
    .A(\nibble_mayor.nibble_C [2]),
    .B(_764_),
    .Y(_765_)
);

INVX1 _1065_ (
    .A(DATA_B[16]),
    .Y(_250_)
);

OR2X2 _1294_ (
    .A(SEL_A_11_bF$buf3),
    .B(DATA_A[10]),
    .Y(_625_)
);

NOR3X1 _1579_ (
    .A(_701_),
    .B(_702_),
    .C(_706_),
    .Y(_728_)
);

NAND2X1 _1159_ (
    .A(SEL_B[7]),
    .B(_338_),
    .Y(_339_)
);

INVX1 _1388_ (
    .A(DATA_B[20]),
    .Y(_559_)
);

OAI21X1 _1600_ (
    .A(_638_[1]),
    .B(_693_),
    .C(_745_),
    .Y(_639_[2])
);

NAND3X1 _931_ (
    .A(_4_),
    .B(_119_),
    .C(_121_),
    .Y(_122_)
);

OAI21X1 _1197_ (
    .A(_374_),
    .B(SEL_B_8_bF$buf2),
    .C(_375_),
    .Y(_376_)
);

BUFX2 BUFX2_insert20 (
    .A(SEL_B[2]),
    .Y(SEL_B_2_bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(SEL_B[2]),
    .Y(SEL_B_2_bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(SEL_B[2]),
    .Y(SEL_B_2_bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(SEL_B[2]),
    .Y(SEL_B_2_bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(SEL_B[2]),
    .Y(SEL_B_2_bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(SEL_A[5]),
    .Y(SEL_A_5_bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .A(SEL_A[5]),
    .Y(SEL_A_5_bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(SEL_A[5]),
    .Y(SEL_A_5_bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(SEL_A[5]),
    .Y(SEL_A_5_bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(SEL_A[5]),
    .Y(SEL_A_5_bF$buf0)
);

INVX2 _1503_ (
    .A(\nibble_mayor.nibble_B [1]),
    .Y(_652_)
);

NAND3X1 _834_ (
    .A(_141_),
    .B(_24_),
    .C(_26_),
    .Y(_27_)
);

NAND3X1 _1312_ (
    .A(_481_),
    .B(_482_),
    .C(_484_),
    .Y(_485_)
);

NAND3X1 _1541_ (
    .A(_688_),
    .B(_679_),
    .C(_689_),
    .Y(_690_)
);

INVX4 _1121_ (
    .A(SEL_A[7]),
    .Y(_459_)
);

NAND2X1 _872_ (
    .A(SEL_A_2_bF$buf4),
    .B(_63_),
    .Y(_64_)
);

OR2X2 _928_ (
    .A(SEL_B_2_bF$buf2),
    .B(DATA_B[5]),
    .Y(_119_)
);

NAND2X1 _1350_ (
    .A(SEL_B_11_bF$buf0),
    .B(_521_),
    .Y(_522_)
);

AOI21X1 _1406_ (
    .A(_557_),
    .B(_576_),
    .C(_615_),
    .Y(_479_[0])
);

INVX1 _1215_ (
    .A(DATA_A[12]),
    .Y(_393_)
);

INVX1 _966_ (
    .A(DATA_A[22]),
    .Y(_311_)
);

NAND3X1 _1444_ (
    .A(SEL_AB[3]),
    .B(_604_),
    .C(_613_),
    .Y(_614_)
);

NAND3X1 _1024_ (
    .A(SEL_B[3]),
    .B(_205_),
    .C(_209_),
    .Y(_210_)
);

AND2X2 _775_ (
    .A(RESET_L_bF$buf2),
    .B(NIBBLE_MAYOR[1]),
    .Y(_0_[1])
);

NAND3X1 _1253_ (
    .A(_459_),
    .B(_427_),
    .C(_429_),
    .Y(_430_)
);

OR2X2 _1309_ (
    .A(DATA_B[2]),
    .B(SEL_B_11_bF$buf0),
    .Y(_482_)
);

NOR2X1 _1482_ (
    .A(\nibble_mayor.nibble_C [3]),
    .B(\nibble_mayor.nibble_D [3]),
    .Y(_762_)
);

NAND3X1 _1062_ (
    .A(SEL_B[4]),
    .B(_246_),
    .C(_245_),
    .Y(_247_)
);

OAI21X1 _1538_ (
    .A(_685_),
    .B(_684_),
    .C(_686_),
    .Y(_687_)
);

INVX2 _1118_ (
    .A(RESET_L_bF$buf0),
    .Y(_456_)
);

AOI21X1 _869_ (
    .A(_42_),
    .B(_61_),
    .C(_138_),
    .Y(_2_[3])
);

NAND3X1 _1291_ (
    .A(_618_),
    .B(_619_),
    .C(_621_),
    .Y(_622_)
);

NAND3X1 _1347_ (
    .A(_616_),
    .B(_509_),
    .C(_518_),
    .Y(_519_)
);

NOR3X1 _1576_ (
    .A(_694_),
    .B(_695_),
    .C(_679_),
    .Y(_725_)
);

INVX1 _1156_ (
    .A(DATA_B[14]),
    .Y(_336_)
);

NAND3X1 _1385_ (
    .A(SEL_A[9]),
    .B(_551_),
    .C(_555_),
    .Y(_556_)
);

NAND3X1 _1194_ (
    .A(_322_),
    .B(_370_),
    .C(_372_),
    .Y(_373_)
);

OAI21X1 _1479_ (
    .A(\nibble_mayor.nibble_C [1]),
    .B(_755_),
    .C(_758_),
    .Y(_759_)
);

INVX1 _1059_ (
    .A(DATA_B[28]),
    .Y(_244_)
);

OR2X2 _1288_ (
    .A(SEL_A_11_bF$buf4),
    .B(DATA_A[2]),
    .Y(_619_)
);

INVX2 _1500_ (
    .A(\nibble_mayor.nibble_B [2]),
    .Y(_649_)
);

OR2X2 _831_ (
    .A(DATA_A[3]),
    .B(SEL_A_2_bF$buf3),
    .Y(_24_)
);

NAND3X1 _1097_ (
    .A(_163_),
    .B(_278_),
    .C(_280_),
    .Y(_281_)
);

NAND2X1 _925_ (
    .A(SEL_A[1]),
    .B(_115_),
    .Y(_116_)
);

NAND2X1 _1403_ (
    .A(SEL_B[10]),
    .B(_573_),
    .Y(_574_)
);

INVX1 _1212_ (
    .A(DATA_A[20]),
    .Y(_390_)
);

NAND3X1 _963_ (
    .A(SEL_A[4]),
    .B(_307_),
    .C(_306_),
    .Y(_308_)
);

OAI21X1 _1441_ (
    .A(_609_),
    .B(SEL_B_11_bF$buf4),
    .C(_610_),
    .Y(_611_)
);

NAND2X1 _1021_ (
    .A(SEL_B_5_bF$buf0),
    .B(_206_),
    .Y(_207_)
);

NAND3X1 _828_ (
    .A(SEL_B[0]),
    .B(_17_),
    .C(_21_),
    .Y(_22_)
);

OR2X2 _1250_ (
    .A(SEL_A_8_bF$buf4),
    .B(DATA_A[5]),
    .Y(_427_)
);

NAND3X1 _1306_ (
    .A(_616_),
    .B(_627_),
    .C(_636_),
    .Y(_637_)
);

AOI21X1 _1535_ (
    .A(_683_),
    .B(_758_),
    .C(_682_),
    .Y(_684_)
);

DFFPOSX1 _1115_ (
    .Q(NIBBLES[5]),
    .CLK(CLK_bF$buf1),
    .D(_161_[1])
);

NAND2X1 _866_ (
    .A(SEL_B[1]),
    .B(_58_),
    .Y(_59_)
);

OAI21X1 _1344_ (
    .A(_514_),
    .B(SEL_A_11_bF$buf0),
    .C(_515_),
    .Y(_516_)
);

NAND3X1 _1573_ (
    .A(_693_),
    .B(_688_),
    .C(_689_),
    .Y(_722_)
);

INVX1 _1153_ (
    .A(DATA_B[22]),
    .Y(_333_)
);

FILL FILL_16_1 (
);

FILL FILL_16_2 (
);

NAND3X1 _1209_ (
    .A(SEL_A[7]),
    .B(_386_),
    .C(_385_),
    .Y(_387_)
);

NAND2X1 _1382_ (
    .A(SEL_A_11_bF$buf2),
    .B(DATA_A[28]),
    .Y(_553_)
);

NAND3X1 _1438_ (
    .A(_481_),
    .B(_605_),
    .C(_607_),
    .Y(_608_)
);

NAND2X1 _1018_ (
    .A(SEL_B_5_bF$buf0),
    .B(_203_),
    .Y(_204_)
);

OR2X2 _1191_ (
    .A(SEL_B_8_bF$buf0),
    .B(DATA_B[3]),
    .Y(_370_)
);

OR2X2 _1247_ (
    .A(SEL_A_8_bF$buf0),
    .B(DATA_A[9]),
    .Y(_424_)
);

INVX1 _998_ (
    .A(DATA_A[19]),
    .Y(_184_)
);

INVX2 _1476_ (
    .A(\nibble_mayor.nibble_C [1]),
    .Y(_756_)
);

INVX1 _1056_ (
    .A(DATA_B[20]),
    .Y(_241_)
);

INVX2 _1285_ (
    .A(SEL_AB[3]),
    .Y(_616_)
);

OR2X2 _1094_ (
    .A(SEL_B_5_bF$buf1),
    .B(DATA_B[5]),
    .Y(_278_)
);

NAND2X1 _1379_ (
    .A(SEL_A_11_bF$buf2),
    .B(_549_),
    .Y(_550_)
);

FILL FILL_6_1 (
);

INVX1 _922_ (
    .A(DATA_A[13]),
    .Y(_113_)
);

OR2X2 _1188_ (
    .A(SEL_B_8_bF$buf1),
    .B(DATA_B[15]),
    .Y(_367_)
);

INVX1 _1400_ (
    .A(DATA_B[8]),
    .Y(_571_)
);

FILL FILL_11_1_0 (
);

FILL FILL_11_1_1 (
);

INVX1 _960_ (
    .A(DATA_A[26]),
    .Y(_305_)
);

NAND2X1 _825_ (
    .A(SEL_B_2_bF$buf4),
    .B(DATA_B[30]),
    .Y(_19_)
);

OAI21X1 _1303_ (
    .A(_632_),
    .B(SEL_A_11_bF$buf2),
    .C(_633_),
    .Y(_634_)
);

AND2X2 _1532_ (
    .A(\nibble_mayor.nibble_C [2]),
    .B(\nibble_mayor.nibble_D [2]),
    .Y(_681_)
);

NAND3X1 _1112_ (
    .A(SEL_AB[1]),
    .B(_286_),
    .C(_295_),
    .Y(_296_)
);

INVX1 _863_ (
    .A(DATA_B[11]),
    .Y(_56_)
);

FILL FILL_8_1_0 (
);

FILL FILL_8_1_1 (
);

INVX1 _919_ (
    .A(DATA_A[21]),
    .Y(_110_)
);

NAND3X1 _1341_ (
    .A(_618_),
    .B(_510_),
    .C(_512_),
    .Y(_513_)
);

NAND3X1 _1570_ (
    .A(_717_),
    .B(_718_),
    .C(_716_),
    .Y(_719_)
);

NAND3X1 _1150_ (
    .A(SEL_B[7]),
    .B(_329_),
    .C(_328_),
    .Y(_330_)
);

FILL FILL_3_1_0 (
);

FILL FILL_3_1_1 (
);

INVX1 _1206_ (
    .A(DATA_A[24]),
    .Y(_384_)
);

INVX1 _957_ (
    .A(DATA_A[18]),
    .Y(_302_)
);

OR2X2 _1435_ (
    .A(SEL_B_11_bF$buf2),
    .B(DATA_B[1]),
    .Y(_605_)
);

NAND3X1 _1015_ (
    .A(_298_),
    .B(_191_),
    .C(_200_),
    .Y(_201_)
);

NAND3X1 _1244_ (
    .A(_459_),
    .B(_418_),
    .C(_420_),
    .Y(_421_)
);

NAND3X1 _995_ (
    .A(SEL_AB[1]),
    .B(_172_),
    .C(_181_),
    .Y(_182_)
);

INVX1 _1473_ (
    .A(_752_),
    .Y(_753_)
);

NAND3X1 _1053_ (
    .A(SEL_A[3]),
    .B(_233_),
    .C(_237_),
    .Y(_238_)
);

FILL FILL_13_0_0 (
);

FILL FILL_13_0_1 (
);

NAND2X1 _1529_ (
    .A(\nibble_mayor.nibble_A [2]),
    .B(_677_),
    .Y(_678_)
);

OAI21X1 _1109_ (
    .A(_291_),
    .B(SEL_B_5_bF$buf1),
    .C(_292_),
    .Y(_293_)
);

DFFPOSX1 _1282_ (
    .Q(NIBBLES[10]),
    .CLK(CLK_bF$buf0),
    .D(_320_[2])
);

OR2X2 _1338_ (
    .A(SEL_A_11_bF$buf0),
    .B(DATA_A[7]),
    .Y(_510_)
);

NAND2X1 _1091_ (
    .A(SEL_A[4]),
    .B(_274_),
    .Y(_275_)
);

AOI21X1 _1567_ (
    .A(_673_),
    .B(_677_),
    .C(_712_),
    .Y(_716_)
);

INVX1 _1147_ (
    .A(DATA_B[26]),
    .Y(_327_)
);

OR2X2 _898_ (
    .A(SEL_B_2_bF$buf3),
    .B(DATA_B[0]),
    .Y(_90_)
);

NAND3X1 _1376_ (
    .A(_617_),
    .B(_542_),
    .C(_546_),
    .Y(_547_)
);

NAND3X1 _1185_ (
    .A(_322_),
    .B(_361_),
    .C(_363_),
    .Y(_364_)
);

FILL FILL_5_0_0 (
);

FILL FILL_5_0_1 (
);

AOI21X1 _1279_ (
    .A(_436_),
    .B(_455_),
    .C(_456_),
    .Y(_320_[1])
);

FILL FILL_0_0_0 (
);

FILL FILL_0_0_1 (
);

NAND2X1 _822_ (
    .A(SEL_B_2_bF$buf4),
    .B(_15_),
    .Y(_16_)
);

INVX1 _1088_ (
    .A(DATA_A[13]),
    .Y(_272_)
);

NAND3X1 _1300_ (
    .A(_618_),
    .B(_628_),
    .C(_630_),
    .Y(_631_)
);

INVX1 _860_ (
    .A(DATA_B[19]),
    .Y(_53_)
);

NAND3X1 _916_ (
    .A(SEL_A[1]),
    .B(_106_),
    .C(_105_),
    .Y(_107_)
);

INVX1 _1203_ (
    .A(DATA_A[16]),
    .Y(_381_)
);

INVX2 _954_ (
    .A(SEL_A[3]),
    .Y(_299_)
);

OR2X2 _1432_ (
    .A(SEL_B_11_bF$buf3),
    .B(DATA_B[13]),
    .Y(_602_)
);

OAI21X1 _1012_ (
    .A(_196_),
    .B(SEL_A_5_bF$buf3),
    .C(_197_),
    .Y(_198_)
);

NAND3X1 _819_ (
    .A(_3_),
    .B(_8_),
    .C(_12_),
    .Y(_13_)
);

OR2X2 _1241_ (
    .A(SEL_A_8_bF$buf0),
    .B(DATA_A[1]),
    .Y(_418_)
);

OAI21X1 _992_ (
    .A(_177_),
    .B(SEL_B_5_bF$buf4),
    .C(_178_),
    .Y(_179_)
);

NAND2X1 _1470_ (
    .A(\nibble_mayor.nibble_C [3]),
    .B(\nibble_mayor.nibble_D [3]),
    .Y(_750_)
);

NAND2X1 _1050_ (
    .A(SEL_A_5_bF$buf1),
    .B(DATA_A[28]),
    .Y(_235_)
);

AOI22X1 _1526_ (
    .A(_651_),
    .B(\nibble_mayor.nibble_A [3]),
    .C(\nibble_mayor.nibble_A [2]),
    .D(_649_),
    .Y(_675_)
);

NAND3X1 _1106_ (
    .A(_163_),
    .B(_287_),
    .C(_289_),
    .Y(_290_)
);

NAND3X1 _857_ (
    .A(SEL_B[1]),
    .B(_49_),
    .C(_48_),
    .Y(_50_)
);

OR2X2 _1335_ (
    .A(SEL_A_11_bF$buf4),
    .B(DATA_A[11]),
    .Y(_507_)
);

NOR2X1 _1564_ (
    .A(\nibble_mayor.nibble_C [0]),
    .B(_644_),
    .Y(_713_)
);

INVX1 _1144_ (
    .A(DATA_B[18]),
    .Y(_324_)
);

OR2X2 _895_ (
    .A(SEL_B_2_bF$buf0),
    .B(DATA_B[12]),
    .Y(_87_)
);

NAND2X1 _1373_ (
    .A(SEL_A_11_bF$buf4),
    .B(_543_),
    .Y(_544_)
);

NAND3X1 _1429_ (
    .A(_481_),
    .B(_596_),
    .C(_598_),
    .Y(_599_)
);

NAND3X1 _1009_ (
    .A(_300_),
    .B(_192_),
    .C(_194_),
    .Y(_195_)
);

OR2X2 _1182_ (
    .A(SEL_B_8_bF$buf3),
    .B(DATA_B[7]),
    .Y(_361_)
);

NAND3X1 _1238_ (
    .A(_321_),
    .B(_411_),
    .C(_415_),
    .Y(_416_)
);

NAND3X1 _989_ (
    .A(_163_),
    .B(_173_),
    .C(_175_),
    .Y(_176_)
);

INVX1 _1467_ (
    .A(\nibble_mayor.nibble_C [3]),
    .Y(_747_)
);

NAND2X1 _1047_ (
    .A(SEL_A_5_bF$buf1),
    .B(_231_),
    .Y(_232_)
);

NAND3X1 _798_ (
    .A(_140_),
    .B(_145_),
    .C(_149_),
    .Y(_150_)
);

NAND2X1 _1276_ (
    .A(SEL_B[7]),
    .B(_452_),
    .Y(_453_)
);

INVX1 _1085_ (
    .A(DATA_A[21]),
    .Y(_269_)
);

INVX1 _913_ (
    .A(DATA_A[25]),
    .Y(_104_)
);

NAND3X1 _1599_ (
    .A(_744_),
    .B(_721_),
    .C(_732_),
    .Y(_745_)
);

NAND2X1 _1179_ (
    .A(SEL_A[7]),
    .B(_357_),
    .Y(_358_)
);

DFFPOSX1 _1620_ (
    .Q(\nibble_mayor.nibble_D [3]),
    .CLK(CLK_bF$buf0),
    .D(_643_[3])
);

NAND3X1 _1200_ (
    .A(SEL_AB[2]),
    .B(_369_),
    .C(_378_),
    .Y(_379_)
);

DFFPOSX1 _951_ (
    .Q(NIBBLES[3]),
    .CLK(CLK_bF$buf1),
    .D(_2_[3])
);

NAND2X1 _816_ (
    .A(SEL_B_2_bF$buf1),
    .B(_9_),
    .Y(_10_)
);

NOR2X1 _1523_ (
    .A(\nibble_mayor.nibble_B [1]),
    .B(_669_),
    .Y(_672_)
);

OR2X2 _1103_ (
    .A(SEL_B_5_bF$buf4),
    .B(DATA_B[1]),
    .Y(_287_)
);

FILL FILL_11_1 (
);

INVX1 _854_ (
    .A(DATA_B[31]),
    .Y(_47_)
);

FILL FILL_11_2 (
);

NAND3X1 _1332_ (
    .A(_618_),
    .B(_501_),
    .C(_503_),
    .Y(_504_)
);

INVX1 _1561_ (
    .A(_677_),
    .Y(_710_)
);

INVX2 _1141_ (
    .A(SEL_B[6]),
    .Y(_321_)
);

NAND3X1 _892_ (
    .A(_4_),
    .B(_81_),
    .C(_83_),
    .Y(_84_)
);

DFFPOSX1 _1617_ (
    .Q(\nibble_mayor.nibble_D [0]),
    .CLK(CLK_bF$buf5),
    .D(_643_[0])
);

DFFPOSX1 _948_ (
    .Q(NIBBLES[0]),
    .CLK(CLK_bF$buf0),
    .D(_2_[0])
);

NAND2X1 _1370_ (
    .A(SEL_A_11_bF$buf1),
    .B(_540_),
    .Y(_541_)
);

OR2X2 _1426_ (
    .A(SEL_B_11_bF$buf4),
    .B(DATA_B[5]),
    .Y(_596_)
);

OR2X2 _1006_ (
    .A(SEL_A_5_bF$buf4),
    .B(DATA_A[7]),
    .Y(_192_)
);

NAND2X1 _1235_ (
    .A(SEL_B_8_bF$buf1),
    .B(DATA_B[24]),
    .Y(_413_)
);

OR2X2 _986_ (
    .A(SEL_B_5_bF$buf3),
    .B(DATA_B[6]),
    .Y(_173_)
);

AND2X2 _1464_ (
    .A(RESET_L_bF$buf1),
    .B(NIBBLES[2]),
    .Y(_640_[2])
);

NAND3X1 _1044_ (
    .A(_299_),
    .B(_224_),
    .C(_228_),
    .Y(_229_)
);

NAND2X1 _795_ (
    .A(SEL_A_2_bF$buf4),
    .B(_146_),
    .Y(_147_)
);

INVX1 _1273_ (
    .A(DATA_B[9]),
    .Y(_450_)
);

OR2X2 _1329_ (
    .A(DATA_A[3]),
    .B(SEL_A_11_bF$buf4),
    .Y(_501_)
);

FILL FILL_1_1 (
);

NAND3X1 _1082_ (
    .A(SEL_A[4]),
    .B(_265_),
    .C(_264_),
    .Y(_266_)
);

NAND2X1 _1558_ (
    .A(_756_),
    .B(_687_),
    .Y(_707_)
);

NAND2X1 _1138_ (
    .A(SEL_A[7]),
    .B(_475_),
    .Y(_476_)
);

OR2X2 _889_ (
    .A(SEL_B_2_bF$buf0),
    .B(DATA_B[4]),
    .Y(_81_)
);

AOI21X1 _1367_ (
    .A(_519_),
    .B(_538_),
    .C(_615_),
    .Y(_479_[3])
);

INVX1 _910_ (
    .A(DATA_A[17]),
    .Y(_101_)
);

NAND3X1 _1596_ (
    .A(_742_),
    .B(_721_),
    .C(_732_),
    .Y(_743_)
);

INVX1 _1176_ (
    .A(DATA_A[15]),
    .Y(_355_)
);

NAND2X1 _813_ (
    .A(SEL_B_2_bF$buf3),
    .B(_6_),
    .Y(_7_)
);

INVX1 _1499_ (
    .A(_647_),
    .Y(_648_)
);

INVX1 _1079_ (
    .A(DATA_A[25]),
    .Y(_263_)
);

INVX1 _1520_ (
    .A(\nibble_mayor.nibble_A [1]),
    .Y(_669_)
);

OR2X2 _1100_ (
    .A(SEL_B_5_bF$buf1),
    .B(DATA_B[13]),
    .Y(_284_)
);

INVX1 _851_ (
    .A(DATA_B[23]),
    .Y(_44_)
);

NAND3X1 _907_ (
    .A(SEL_AB[0]),
    .B(_89_),
    .C(_98_),
    .Y(_99_)
);

DFFPOSX1 _1614_ (
    .Q(\nibble_mayor.nibble_C [1]),
    .CLK(CLK_bF$buf5),
    .D(_642_[1])
);

NAND3X1 _945_ (
    .A(_3_),
    .B(_131_),
    .C(_135_),
    .Y(_136_)
);

CLKBUF1 CLKBUF1_insert45 (
    .A(CLK),
    .Y(CLK_bF$buf5)
);

CLKBUF1 CLKBUF1_insert46 (
    .A(CLK),
    .Y(CLK_bF$buf4)
);

CLKBUF1 CLKBUF1_insert47 (
    .A(CLK),
    .Y(CLK_bF$buf3)
);

CLKBUF1 CLKBUF1_insert48 (
    .A(CLK),
    .Y(CLK_bF$buf2)
);

CLKBUF1 CLKBUF1_insert49 (
    .A(CLK),
    .Y(CLK_bF$buf1)
);

NAND2X1 _1423_ (
    .A(SEL_A[10]),
    .B(_592_),
    .Y(_593_)
);

OR2X2 _1003_ (
    .A(SEL_A_5_bF$buf4),
    .B(DATA_A[11]),
    .Y(_189_)
);

NAND2X1 _1232_ (
    .A(SEL_B_8_bF$buf1),
    .B(_409_),
    .Y(_410_)
);

OR2X2 _983_ (
    .A(SEL_B_5_bF$buf0),
    .B(DATA_B[10]),
    .Y(_170_)
);

AND2X2 _1461_ (
    .A(RESET_L_bF$buf3),
    .B(NIBBLES[7]),
    .Y(_641_[3])
);

NAND2X1 _1041_ (
    .A(SEL_A_5_bF$buf2),
    .B(_225_),
    .Y(_226_)
);

NAND2X1 _792_ (
    .A(SEL_A_2_bF$buf4),
    .B(_143_),
    .Y(_144_)
);

AOI21X1 _1517_ (
    .A(_663_),
    .B(_665_),
    .C(_664_),
    .Y(_666_)
);

NAND3X1 _848_ (
    .A(SEL_A[0]),
    .B(_36_),
    .C(_40_),
    .Y(_41_)
);

INVX1 _1270_ (
    .A(DATA_B[17]),
    .Y(_447_)
);

NAND3X1 _1326_ (
    .A(SEL_B[9]),
    .B(_494_),
    .C(_498_),
    .Y(_499_)
);

NAND3X1 _1555_ (
    .A(\nibble_mayor.nibble_B [1]),
    .B(_666_),
    .C(_662_),
    .Y(_704_)
);

INVX1 _1135_ (
    .A(DATA_A[14]),
    .Y(_473_)
);

NAND2X1 _886_ (
    .A(SEL_A[1]),
    .B(_77_),
    .Y(_78_)
);

NAND2X1 _1364_ (
    .A(SEL_B[10]),
    .B(_535_),
    .Y(_536_)
);

NAND2X1 _1593_ (
    .A(_716_),
    .B(_739_),
    .Y(_741_)
);

INVX1 _1173_ (
    .A(DATA_A[23]),
    .Y(_352_)
);

NAND3X1 _1229_ (
    .A(SEL_B[6]),
    .B(_402_),
    .C(_406_),
    .Y(_407_)
);

AND2X2 _1458_ (
    .A(RESET_L_bF$buf3),
    .B(NIBBLES[4]),
    .Y(_641_[0])
);

NAND2X1 _1038_ (
    .A(SEL_A_5_bF$buf2),
    .B(_222_),
    .Y(_223_)
);

INVX4 _789_ (
    .A(SEL_A[1]),
    .Y(_141_)
);

NAND3X1 _1267_ (
    .A(SEL_B[7]),
    .B(_443_),
    .C(_442_),
    .Y(_444_)
);

INVX4 _810_ (
    .A(SEL_B[1]),
    .Y(_4_)
);

OAI21X1 _1496_ (
    .A(\nibble_mayor.nibble_C [3]),
    .B(\nibble_mayor.nibble_D [3]),
    .C(RESET_L_bF$buf1),
    .Y(_646_)
);

INVX1 _1076_ (
    .A(DATA_A[17]),
    .Y(_260_)
);

OAI21X1 _904_ (
    .A(_94_),
    .B(SEL_B_2_bF$buf3),
    .C(_95_),
    .Y(_96_)
);

NAND3X1 _1399_ (
    .A(_481_),
    .B(_567_),
    .C(_569_),
    .Y(_570_)
);

FILL FILL_8_1 (
);

DFFPOSX1 _1611_ (
    .Q(\nibble_mayor.nibble_B [2]),
    .CLK(CLK_bF$buf3),
    .D(_641_[2])
);

NAND2X1 _942_ (
    .A(SEL_B_2_bF$buf4),
    .B(DATA_B[25]),
    .Y(_133_)
);

INVX1 _1420_ (
    .A(DATA_A[13]),
    .Y(_590_)
);

NAND3X1 _1000_ (
    .A(_300_),
    .B(_183_),
    .C(_185_),
    .Y(_186_)
);

NAND3X1 _807_ (
    .A(SEL_A[0]),
    .B(_154_),
    .C(_158_),
    .Y(_159_)
);

NAND3X1 _980_ (
    .A(_163_),
    .B(_164_),
    .C(_166_),
    .Y(_167_)
);

NAND2X1 _1514_ (
    .A(\nibble_mayor.nibble_B [3]),
    .B(_658_),
    .Y(_663_)
);

NAND2X1 _845_ (
    .A(SEL_A_2_bF$buf3),
    .B(DATA_A[31]),
    .Y(_38_)
);

NAND2X1 _1323_ (
    .A(SEL_B_11_bF$buf3),
    .B(DATA_B[30]),
    .Y(_496_)
);

AND2X2 _1552_ (
    .A(_687_),
    .B(_756_),
    .Y(_701_)
);

INVX1 _1132_ (
    .A(DATA_A[22]),
    .Y(_470_)
);

INVX1 _883_ (
    .A(DATA_A[12]),
    .Y(_75_)
);

DFFPOSX1 _1608_ (
    .Q(\nibble_mayor.nibble_A [3]),
    .CLK(CLK_bF$buf1),
    .D(_640_[3])
);

NAND2X1 _939_ (
    .A(SEL_B_2_bF$buf4),
    .B(_129_),
    .Y(_130_)
);

INVX1 _1361_ (
    .A(DATA_B[11]),
    .Y(_533_)
);

INVX1 _1417_ (
    .A(DATA_A[21]),
    .Y(_587_)
);

AOI21X1 _1590_ (
    .A(_728_),
    .B(_697_),
    .C(_738_),
    .Y(_739_)
);

NAND3X1 _1170_ (
    .A(SEL_A[7]),
    .B(_348_),
    .C(_347_),
    .Y(_349_)
);

NAND2X1 _1226_ (
    .A(SEL_B_8_bF$buf0),
    .B(_403_),
    .Y(_404_)
);

OR2X2 _977_ (
    .A(DATA_B[2]),
    .B(SEL_B_5_bF$buf4),
    .Y(_164_)
);

AND2X2 _1455_ (
    .A(RESET_L_bF$buf0),
    .B(NIBBLES[9]),
    .Y(_642_[1])
);

AOI21X1 _1035_ (
    .A(_201_),
    .B(_220_),
    .C(_297_),
    .Y(_161_[3])
);

INVX2 _786_ (
    .A(RESET_L_bF$buf4),
    .Y(_138_)
);

INVX1 _1264_ (
    .A(DATA_B[29]),
    .Y(_441_)
);

AOI22X1 _1493_ (
    .A(_769_),
    .B(_768_),
    .C(_770_),
    .D(_772_),
    .Y(_773_)
);

NAND3X1 _1073_ (
    .A(SEL_AB[1]),
    .B(_248_),
    .C(_257_),
    .Y(_258_)
);

NAND2X1 _1549_ (
    .A(_669_),
    .B(_677_),
    .Y(_698_)
);

NAND3X1 _1129_ (
    .A(SEL_A[7]),
    .B(_466_),
    .C(_465_),
    .Y(_467_)
);

INVX1 _1358_ (
    .A(DATA_B[19]),
    .Y(_530_)
);

NAND3X1 _901_ (
    .A(_4_),
    .B(_90_),
    .C(_92_),
    .Y(_93_)
);

NAND3X1 _1587_ (
    .A(_735_),
    .B(_697_),
    .C(_734_),
    .Y(_736_)
);

INVX1 _1167_ (
    .A(DATA_A[27]),
    .Y(_346_)
);

OR2X2 _1396_ (
    .A(SEL_B_11_bF$buf0),
    .B(DATA_B[0]),
    .Y(_567_)
);

NAND2X1 _804_ (
    .A(SEL_A_2_bF$buf1),
    .B(DATA_A[30]),
    .Y(_156_)
);

NAND2X1 _1299_ (
    .A(SEL_A_11_bF$buf2),
    .B(_629_),
    .Y(_630_)
);

OAI22X1 _1511_ (
    .A(_658_),
    .B(\nibble_mayor.nibble_B [3]),
    .C(_659_),
    .D(\nibble_mayor.nibble_B [2]),
    .Y(_660_)
);

NAND2X1 _842_ (
    .A(SEL_A_2_bF$buf3),
    .B(_34_),
    .Y(_35_)
);

NAND2X1 _1320_ (
    .A(SEL_B_11_bF$buf3),
    .B(_492_),
    .Y(_493_)
);

FILL FILL_15_1_0 (
);

FILL FILL_15_1_1 (
);

INVX1 _880_ (
    .A(DATA_A[20]),
    .Y(_72_)
);

DFFPOSX1 _1605_ (
    .Q(\nibble_mayor.nibble_A [0]),
    .CLK(CLK_bF$buf5),
    .D(_640_[0])
);

NAND3X1 _936_ (
    .A(SEL_B[0]),
    .B(_122_),
    .C(_126_),
    .Y(_127_)
);

FILL FILL_10_1_0 (
);

FILL FILL_10_1_1 (
);

NAND3X1 _1414_ (
    .A(SEL_A[10]),
    .B(_583_),
    .C(_582_),
    .Y(_584_)
);

NAND2X1 _1223_ (
    .A(SEL_B_8_bF$buf4),
    .B(_400_),
    .Y(_401_)
);

NAND3X1 _974_ (
    .A(_298_),
    .B(_309_),
    .C(_318_),
    .Y(_319_)
);

AND2X2 _1452_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLES[14]),
    .Y(_643_[2])
);

NAND2X1 _1032_ (
    .A(SEL_B[4]),
    .B(_217_),
    .Y(_218_)
);

DFFPOSX1 _783_ (
    .Q(_1_[1]),
    .CLK(CLK_bF$buf2),
    .D(_0_[1])
);

NOR2X1 _1508_ (
    .A(\nibble_mayor.nibble_A [0]),
    .B(_656_),
    .Y(_657_)
);

NAND3X1 _839_ (
    .A(_140_),
    .B(_27_),
    .C(_31_),
    .Y(_32_)
);

INVX1 _1261_ (
    .A(DATA_B[21]),
    .Y(_438_)
);

NAND3X1 _1317_ (
    .A(_480_),
    .B(_485_),
    .C(_489_),
    .Y(_490_)
);

NAND2X1 _1490_ (
    .A(\nibble_mayor.nibble_C [0]),
    .B(\nibble_mayor.nibble_D [0]),
    .Y(_770_)
);

OAI21X1 _1070_ (
    .A(_253_),
    .B(SEL_B_5_bF$buf3),
    .C(_254_),
    .Y(_255_)
);

FILL FILL_7_1_0 (
);

FILL FILL_7_1_1 (
);

OAI21X1 _1546_ (
    .A(_687_),
    .B(\nibble_mayor.nibble_D [2]),
    .C(RESET_L_bF$buf2),
    .Y(_695_)
);

INVX1 _1126_ (
    .A(DATA_A[26]),
    .Y(_464_)
);

NAND3X1 _877_ (
    .A(SEL_A[1]),
    .B(_68_),
    .C(_67_),
    .Y(_69_)
);

NAND3X1 _1355_ (
    .A(SEL_B[10]),
    .B(_526_),
    .C(_525_),
    .Y(_527_)
);

FILL FILL_2_1_0 (
);

FILL FILL_2_1_1 (
);

OAI21X1 _1584_ (
    .A(\nibble_mayor.nibble_C [0]),
    .B(_644_),
    .C(_718_),
    .Y(_733_)
);

INVX1 _1164_ (
    .A(DATA_A[19]),
    .Y(_343_)
);

OR2X2 _1393_ (
    .A(SEL_B_11_bF$buf4),
    .B(DATA_B[12]),
    .Y(_564_)
);

DFFPOSX1 _1449_ (
    .Q(NIBBLES[15]),
    .CLK(CLK_bF$buf0),
    .D(_479_[3])
);

INVX1 _1029_ (
    .A(DATA_B[11]),
    .Y(_215_)
);

NAND3X1 _1258_ (
    .A(SEL_A[6]),
    .B(_430_),
    .C(_434_),
    .Y(_435_)
);

FILL FILL_12_0_0 (
);

FILL FILL_12_0_1 (
);

NAND2X1 _801_ (
    .A(SEL_A_2_bF$buf1),
    .B(_152_),
    .Y(_153_)
);

AND2X2 _1487_ (
    .A(_766_),
    .B(_761_),
    .Y(_767_)
);

NAND3X1 _1067_ (
    .A(_163_),
    .B(_249_),
    .C(_251_),
    .Y(_252_)
);

NAND3X1 _1296_ (
    .A(_617_),
    .B(_622_),
    .C(_626_),
    .Y(_627_)
);

FILL FILL_9_0_0 (
);

FILL FILL_9_0_1 (
);

DFFPOSX1 _1602_ (
    .Q(NIBBLE_MAYOR[1]),
    .CLK(CLK_bF$buf4),
    .D(_639_[1])
);

NAND2X1 _933_ (
    .A(SEL_B_2_bF$buf0),
    .B(_123_),
    .Y(_124_)
);

NAND3X1 _1199_ (
    .A(_321_),
    .B(_373_),
    .C(_377_),
    .Y(_378_)
);

FILL FILL_4_0_0 (
);

FILL FILL_4_0_1 (
);

INVX1 _1411_ (
    .A(DATA_A[25]),
    .Y(_581_)
);

BUFX2 BUFX2_insert40 (
    .A(RESET_L),
    .Y(RESET_L_bF$buf4)
);

BUFX2 BUFX2_insert41 (
    .A(RESET_L),
    .Y(RESET_L_bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(RESET_L),
    .Y(RESET_L_bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(RESET_L),
    .Y(RESET_L_bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(RESET_L),
    .Y(RESET_L_bF$buf0)
);

NAND3X1 _1220_ (
    .A(_457_),
    .B(_388_),
    .C(_397_),
    .Y(_398_)
);

OAI21X1 _971_ (
    .A(_314_),
    .B(SEL_A_5_bF$buf0),
    .C(_315_),
    .Y(_316_)
);

BUFX2 _780_ (
    .A(_1_[2]),
    .Y(DATA_OUT[2])
);

NOR2X1 _1505_ (
    .A(_650_),
    .B(_653_),
    .Y(_654_)
);

NAND2X1 _836_ (
    .A(SEL_A_2_bF$buf0),
    .B(_28_),
    .Y(_29_)
);

NAND2X1 _1314_ (
    .A(SEL_B_11_bF$buf1),
    .B(_486_),
    .Y(_487_)
);

NAND3X1 _1543_ (
    .A(_649_),
    .B(_666_),
    .C(_662_),
    .Y(_692_)
);

INVX1 _1123_ (
    .A(DATA_A[18]),
    .Y(_461_)
);

INVX1 _874_ (
    .A(DATA_A[24]),
    .Y(_66_)
);

INVX1 _1352_ (
    .A(DATA_B[31]),
    .Y(_524_)
);

INVX1 _1408_ (
    .A(DATA_A[17]),
    .Y(_578_)
);

OAI21X1 _1581_ (
    .A(_713_),
    .B(_714_),
    .C(_716_),
    .Y(_730_)
);

NAND3X1 _1161_ (
    .A(SEL_AB[2]),
    .B(_331_),
    .C(_340_),
    .Y(_341_)
);

OAI21X1 _1217_ (
    .A(_393_),
    .B(SEL_A_8_bF$buf4),
    .C(_394_),
    .Y(_395_)
);

NAND3X1 _968_ (
    .A(_300_),
    .B(_310_),
    .C(_312_),
    .Y(_313_)
);

NAND3X1 _1390_ (
    .A(_481_),
    .B(_558_),
    .C(_560_),
    .Y(_561_)
);

DFFPOSX1 _1446_ (
    .Q(NIBBLES[12]),
    .CLK(CLK_bF$buf3),
    .D(_479_[0])
);

INVX1 _1026_ (
    .A(DATA_B[19]),
    .Y(_212_)
);

AND2X2 _777_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLE_MAYOR[3]),
    .Y(_0_[3])
);

NAND2X1 _1255_ (
    .A(SEL_A_8_bF$buf4),
    .B(DATA_A[29]),
    .Y(_432_)
);

INVX1 _1484_ (
    .A(\nibble_mayor.nibble_D [2]),
    .Y(_764_)
);

OR2X2 _1064_ (
    .A(SEL_B_5_bF$buf3),
    .B(DATA_B[0]),
    .Y(_249_)
);

NAND2X1 _1293_ (
    .A(SEL_A_11_bF$buf1),
    .B(_623_),
    .Y(_624_)
);

INVX1 _1349_ (
    .A(DATA_B[23]),
    .Y(_521_)
);

FILL FILL_3_1 (
);

FILL FILL_3_2 (
);

AOI22X1 _1578_ (
    .A(_645_),
    .B(_726_),
    .C(_725_),
    .D(_647_),
    .Y(_727_)
);

OAI21X1 _1158_ (
    .A(_336_),
    .B(SEL_B_8_bF$buf4),
    .C(_337_),
    .Y(_338_)
);

OR2X2 _1387_ (
    .A(SEL_B_11_bF$buf2),
    .B(DATA_B[4]),
    .Y(_558_)
);

NAND2X1 _930_ (
    .A(SEL_B_2_bF$buf0),
    .B(_120_),
    .Y(_121_)
);

NAND2X1 _1196_ (
    .A(SEL_B_8_bF$buf2),
    .B(DATA_B[27]),
    .Y(_375_)
);

BUFX2 BUFX2_insert10 (
    .A(SEL_B[5]),
    .Y(SEL_B_5_bF$buf4)
);

BUFX2 BUFX2_insert11 (
    .A(SEL_B[5]),
    .Y(SEL_B_5_bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .A(SEL_B[5]),
    .Y(SEL_B_5_bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .A(SEL_B[5]),
    .Y(SEL_B_5_bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .A(SEL_B[5]),
    .Y(SEL_B_5_bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .A(SEL_A[8]),
    .Y(SEL_A_8_bF$buf4)
);

BUFX2 BUFX2_insert16 (
    .A(SEL_A[8]),
    .Y(SEL_A_8_bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .A(SEL_A[8]),
    .Y(SEL_A_8_bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .A(SEL_A[8]),
    .Y(SEL_A_8_bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .A(SEL_A[8]),
    .Y(SEL_A_8_bF$buf0)
);

INVX1 _1502_ (
    .A(\nibble_mayor.nibble_B [3]),
    .Y(_651_)
);

NAND2X1 _833_ (
    .A(SEL_A_2_bF$buf3),
    .B(_25_),
    .Y(_26_)
);

NAND2X1 _1099_ (
    .A(SEL_B_5_bF$buf2),
    .B(_282_),
    .Y(_283_)
);

NAND2X1 _1311_ (
    .A(SEL_B_11_bF$buf0),
    .B(_483_),
    .Y(_484_)
);

AOI21X1 _1540_ (
    .A(_764_),
    .B(_644_),
    .C(_746_),
    .Y(_689_)
);

INVX2 _1120_ (
    .A(SEL_A[6]),
    .Y(_458_)
);

INVX1 _871_ (
    .A(DATA_A[16]),
    .Y(_63_)
);

NAND3X1 _927_ (
    .A(_139_),
    .B(_108_),
    .C(_117_),
    .Y(_118_)
);

NAND3X1 _1405_ (
    .A(SEL_AB[3]),
    .B(_566_),
    .C(_575_),
    .Y(_576_)
);

NAND3X1 _1214_ (
    .A(_459_),
    .B(_389_),
    .C(_391_),
    .Y(_392_)
);

OR2X2 _965_ (
    .A(SEL_A_5_bF$buf0),
    .B(DATA_A[6]),
    .Y(_310_)
);

NAND3X1 _1443_ (
    .A(_480_),
    .B(_608_),
    .C(_612_),
    .Y(_613_)
);

NAND3X1 _1023_ (
    .A(SEL_B[4]),
    .B(_208_),
    .C(_207_),
    .Y(_209_)
);

AND2X2 _774_ (
    .A(RESET_L_bF$buf2),
    .B(NIBBLE_MAYOR[0]),
    .Y(_0_[0])
);

NAND2X1 _1252_ (
    .A(SEL_A_8_bF$buf4),
    .B(_428_),
    .Y(_429_)
);

INVX4 _1308_ (
    .A(SEL_B[10]),
    .Y(_481_)
);

NAND2X1 _1481_ (
    .A(\nibble_mayor.nibble_D [3]),
    .B(_747_),
    .Y(_761_)
);

OR2X2 _1061_ (
    .A(SEL_B_5_bF$buf4),
    .B(DATA_B[12]),
    .Y(_246_)
);

NAND2X1 _1537_ (
    .A(_773_),
    .B(_754_),
    .Y(_686_)
);

DFFPOSX1 _1117_ (
    .Q(NIBBLES[7]),
    .CLK(CLK_bF$buf1),
    .D(_161_[3])
);

NAND3X1 _868_ (
    .A(SEL_AB[0]),
    .B(_51_),
    .C(_60_),
    .Y(_61_)
);

NAND2X1 _1290_ (
    .A(SEL_A_11_bF$buf4),
    .B(_620_),
    .Y(_621_)
);

NAND3X1 _1346_ (
    .A(SEL_A[9]),
    .B(_513_),
    .C(_517_),
    .Y(_518_)
);

NAND3X1 _1575_ (
    .A(_647_),
    .B(_723_),
    .C(_722_),
    .Y(_724_)
);

NAND3X1 _1155_ (
    .A(_322_),
    .B(_332_),
    .C(_334_),
    .Y(_335_)
);

NAND2X1 _1384_ (
    .A(SEL_A[10]),
    .B(_554_),
    .Y(_555_)
);

NAND2X1 _1193_ (
    .A(SEL_B_8_bF$buf2),
    .B(_371_),
    .Y(_372_)
);

NAND3X1 _1249_ (
    .A(_458_),
    .B(_421_),
    .C(_425_),
    .Y(_426_)
);

OAI22X1 _1478_ (
    .A(_756_),
    .B(\nibble_mayor.nibble_D [1]),
    .C(_757_),
    .D(\nibble_mayor.nibble_D [0]),
    .Y(_758_)
);

NAND3X1 _1058_ (
    .A(_163_),
    .B(_240_),
    .C(_242_),
    .Y(_243_)
);

INVX4 _1287_ (
    .A(SEL_A[10]),
    .Y(_618_)
);

AOI21X1 _830_ (
    .A(_160_),
    .B(_23_),
    .C(_138_),
    .Y(_2_[2])
);

NAND2X1 _1096_ (
    .A(SEL_B_5_bF$buf2),
    .B(_279_),
    .Y(_280_)
);

OAI21X1 _924_ (
    .A(_113_),
    .B(SEL_A_2_bF$buf1),
    .C(_114_),
    .Y(_115_)
);

OAI21X1 _1402_ (
    .A(_571_),
    .B(SEL_B_11_bF$buf1),
    .C(_572_),
    .Y(_573_)
);

OR2X2 _1211_ (
    .A(SEL_A_8_bF$buf4),
    .B(DATA_A[4]),
    .Y(_389_)
);

OR2X2 _962_ (
    .A(SEL_A_5_bF$buf3),
    .B(DATA_A[10]),
    .Y(_307_)
);

NAND2X1 _1440_ (
    .A(SEL_B_11_bF$buf2),
    .B(DATA_B[25]),
    .Y(_610_)
);

INVX1 _1020_ (
    .A(DATA_B[31]),
    .Y(_206_)
);

NAND2X1 _827_ (
    .A(SEL_B[1]),
    .B(_20_),
    .Y(_21_)
);

NAND3X1 _1305_ (
    .A(SEL_A[9]),
    .B(_631_),
    .C(_635_),
    .Y(_636_)
);

NAND2X1 _1534_ (
    .A(\nibble_mayor.nibble_D [1]),
    .B(_756_),
    .Y(_683_)
);

DFFPOSX1 _1114_ (
    .Q(NIBBLES[4]),
    .CLK(CLK_bF$buf1),
    .D(_161_[0])
);

OAI21X1 _865_ (
    .A(_56_),
    .B(SEL_B_2_bF$buf2),
    .C(_57_),
    .Y(_58_)
);

NAND2X1 _1343_ (
    .A(SEL_A_11_bF$buf0),
    .B(DATA_A[31]),
    .Y(_515_)
);

NAND2X1 _1572_ (
    .A(_697_),
    .B(_720_),
    .Y(_721_)
);

OR2X2 _1152_ (
    .A(SEL_B_8_bF$buf4),
    .B(DATA_B[6]),
    .Y(_332_)
);

OR2X2 _1208_ (
    .A(SEL_A_8_bF$buf1),
    .B(DATA_A[8]),
    .Y(_386_)
);

NAND3X1 _959_ (
    .A(_300_),
    .B(_301_),
    .C(_303_),
    .Y(_304_)
);

INVX1 _1381_ (
    .A(DATA_A[12]),
    .Y(_552_)
);

NAND2X1 _1437_ (
    .A(SEL_B_11_bF$buf2),
    .B(_606_),
    .Y(_607_)
);

INVX1 _1017_ (
    .A(DATA_B[23]),
    .Y(_203_)
);

NAND3X1 _1190_ (
    .A(SEL_B[6]),
    .B(_364_),
    .C(_368_),
    .Y(_369_)
);

NAND2X1 _1246_ (
    .A(SEL_A_8_bF$buf0),
    .B(_422_),
    .Y(_423_)
);

OR2X2 _997_ (
    .A(DATA_A[3]),
    .B(SEL_A_5_bF$buf3),
    .Y(_183_)
);

INVX2 _1475_ (
    .A(\nibble_mayor.nibble_D [1]),
    .Y(_755_)
);

OR2X2 _1055_ (
    .A(SEL_B_5_bF$buf3),
    .B(DATA_B[4]),
    .Y(_240_)
);

INVX2 _1284_ (
    .A(RESET_L_bF$buf3),
    .Y(_615_)
);

NAND3X1 _1093_ (
    .A(_298_),
    .B(_267_),
    .C(_276_),
    .Y(_277_)
);

AOI21X1 _1569_ (
    .A(_771_),
    .B(_644_),
    .C(_746_),
    .Y(_718_)
);

OR2X2 _1149_ (
    .A(SEL_B_8_bF$buf3),
    .B(DATA_B[10]),
    .Y(_329_)
);

INVX1 _1378_ (
    .A(DATA_A[20]),
    .Y(_549_)
);

NAND3X1 _921_ (
    .A(_141_),
    .B(_109_),
    .C(_111_),
    .Y(_112_)
);

NAND2X1 _1187_ (
    .A(SEL_B_8_bF$buf1),
    .B(_365_),
    .Y(_366_)
);

INVX1 _824_ (
    .A(DATA_B[14]),
    .Y(_18_)
);

NAND2X1 _1302_ (
    .A(SEL_A_11_bF$buf2),
    .B(DATA_A[30]),
    .Y(_633_)
);

INVX1 _1531_ (
    .A(\nibble_mayor.nibble_C [2]),
    .Y(_680_)
);

NAND3X1 _1111_ (
    .A(_162_),
    .B(_290_),
    .C(_294_),
    .Y(_295_)
);

NAND3X1 _862_ (
    .A(_4_),
    .B(_52_),
    .C(_54_),
    .Y(_55_)
);

OR2X2 _918_ (
    .A(SEL_A_2_bF$buf2),
    .B(DATA_A[5]),
    .Y(_109_)
);

NAND2X1 _1340_ (
    .A(SEL_A_11_bF$buf4),
    .B(_511_),
    .Y(_512_)
);

NAND3X1 _1205_ (
    .A(_459_),
    .B(_380_),
    .C(_382_),
    .Y(_383_)
);

OR2X2 _956_ (
    .A(SEL_A_5_bF$buf2),
    .B(DATA_A[2]),
    .Y(_301_)
);

NAND3X1 _1434_ (
    .A(SEL_B[9]),
    .B(_599_),
    .C(_603_),
    .Y(_604_)
);

NAND3X1 _1014_ (
    .A(SEL_A[3]),
    .B(_195_),
    .C(_199_),
    .Y(_200_)
);

NAND2X1 _1243_ (
    .A(SEL_A_8_bF$buf0),
    .B(_419_),
    .Y(_420_)
);

NAND3X1 _994_ (
    .A(SEL_B[3]),
    .B(_176_),
    .C(_180_),
    .Y(_181_)
);

NOR2X1 _1472_ (
    .A(\nibble_mayor.nibble_C [2]),
    .B(\nibble_mayor.nibble_D [2]),
    .Y(_752_)
);

NAND2X1 _1052_ (
    .A(SEL_A[4]),
    .B(_236_),
    .Y(_237_)
);

OAI21X1 _1528_ (
    .A(_676_),
    .B(_671_),
    .C(_666_),
    .Y(_677_)
);

NAND2X1 _1108_ (
    .A(SEL_B_5_bF$buf2),
    .B(DATA_B[25]),
    .Y(_292_)
);

OR2X2 _859_ (
    .A(SEL_B_2_bF$buf2),
    .B(DATA_B[3]),
    .Y(_52_)
);

DFFPOSX1 _1281_ (
    .Q(NIBBLES[9]),
    .CLK(CLK_bF$buf2),
    .D(_320_[1])
);

NAND3X1 _1337_ (
    .A(_617_),
    .B(_504_),
    .C(_508_),
    .Y(_509_)
);

OAI21X1 _1090_ (
    .A(_272_),
    .B(SEL_A_5_bF$buf1),
    .C(_273_),
    .Y(_274_)
);

OAI22X1 _1566_ (
    .A(_711_),
    .B(_712_),
    .C(_713_),
    .D(_714_),
    .Y(_715_)
);

NAND3X1 _1146_ (
    .A(_322_),
    .B(_323_),
    .C(_325_),
    .Y(_326_)
);

NAND3X1 _897_ (
    .A(SEL_B[0]),
    .B(_84_),
    .C(_88_),
    .Y(_89_)
);

NAND3X1 _1375_ (
    .A(SEL_A[10]),
    .B(_545_),
    .C(_544_),
    .Y(_546_)
);

NAND2X1 _1184_ (
    .A(SEL_B_8_bF$buf3),
    .B(_362_),
    .Y(_363_)
);

NAND2X1 _1469_ (
    .A(_747_),
    .B(_748_),
    .Y(_749_)
);

INVX1 _1049_ (
    .A(DATA_A[12]),
    .Y(_234_)
);

NAND3X1 _1278_ (
    .A(SEL_AB[2]),
    .B(_445_),
    .C(_454_),
    .Y(_455_)
);

INVX1 _821_ (
    .A(DATA_B[22]),
    .Y(_15_)
);

NAND3X1 _1087_ (
    .A(_300_),
    .B(_268_),
    .C(_270_),
    .Y(_271_)
);

OR2X2 _915_ (
    .A(SEL_A_2_bF$buf0),
    .B(DATA_A[9]),
    .Y(_106_)
);

OR2X2 _1202_ (
    .A(SEL_A_8_bF$buf3),
    .B(DATA_A[0]),
    .Y(_380_)
);

INVX2 _953_ (
    .A(SEL_AB[1]),
    .Y(_298_)
);

NAND2X1 _1431_ (
    .A(SEL_B_11_bF$buf3),
    .B(_600_),
    .Y(_601_)
);

NAND2X1 _1011_ (
    .A(SEL_A_5_bF$buf4),
    .B(DATA_A[31]),
    .Y(_197_)
);

NAND3X1 _818_ (
    .A(SEL_B[1]),
    .B(_11_),
    .C(_10_),
    .Y(_12_)
);

AOI21X1 _1240_ (
    .A(_398_),
    .B(_417_),
    .C(_456_),
    .Y(_320_[0])
);

NAND2X1 _991_ (
    .A(SEL_B_5_bF$buf4),
    .B(DATA_B[30]),
    .Y(_178_)
);

NAND2X1 _1525_ (
    .A(\nibble_mayor.nibble_B [0]),
    .B(_673_),
    .Y(_674_)
);

NAND2X1 _1105_ (
    .A(SEL_B_5_bF$buf4),
    .B(_288_),
    .Y(_289_)
);

OR2X2 _856_ (
    .A(SEL_B_2_bF$buf1),
    .B(DATA_B[15]),
    .Y(_49_)
);

FILL FILL_14_1_0 (
);

FILL FILL_14_1_1 (
);

NAND2X1 _1334_ (
    .A(SEL_A_11_bF$buf0),
    .B(_505_),
    .Y(_506_)
);

OAI21X1 _1563_ (
    .A(_677_),
    .B(\nibble_mayor.nibble_B [0]),
    .C(RESET_L_bF$buf1),
    .Y(_712_)
);

OR2X2 _1143_ (
    .A(DATA_B[2]),
    .B(SEL_B_8_bF$buf3),
    .Y(_323_)
);

FILL FILL_15_1 (
);

NAND2X1 _894_ (
    .A(SEL_B_2_bF$buf4),
    .B(_85_),
    .Y(_86_)
);

FILL FILL_15_2 (
);

DFFPOSX1 _1619_ (
    .Q(\nibble_mayor.nibble_D [2]),
    .CLK(CLK_bF$buf0),
    .D(_643_[2])
);

INVX1 _1372_ (
    .A(DATA_A[24]),
    .Y(_543_)
);

NAND2X1 _1428_ (
    .A(SEL_B_11_bF$buf3),
    .B(_597_),
    .Y(_598_)
);

NAND2X1 _1008_ (
    .A(SEL_A_5_bF$buf4),
    .B(_193_),
    .Y(_194_)
);

NAND3X1 _1181_ (
    .A(_457_),
    .B(_350_),
    .C(_359_),
    .Y(_360_)
);

NAND2X1 _1237_ (
    .A(SEL_B[7]),
    .B(_414_),
    .Y(_415_)
);

NAND2X1 _988_ (
    .A(SEL_B_5_bF$buf3),
    .B(_174_),
    .Y(_175_)
);

INVX4 _1466_ (
    .A(RESET_L_bF$buf1),
    .Y(_746_)
);

INVX1 _1046_ (
    .A(DATA_A[20]),
    .Y(_231_)
);

NAND3X1 _797_ (
    .A(SEL_A[1]),
    .B(_148_),
    .C(_147_),
    .Y(_149_)
);

FILL FILL_6_1_0 (
);

FILL FILL_6_1_1 (
);

OAI21X1 _1275_ (
    .A(_450_),
    .B(SEL_B_8_bF$buf4),
    .C(_451_),
    .Y(_452_)
);

OR2X2 _1084_ (
    .A(SEL_A_5_bF$buf0),
    .B(DATA_A[5]),
    .Y(_268_)
);

FILL FILL_1_1_0 (
);

FILL FILL_1_1_1 (
);

INVX1 _1369_ (
    .A(DATA_A[16]),
    .Y(_540_)
);

FILL FILL_5_1 (
);

FILL FILL_5_2 (
);

NAND3X1 _912_ (
    .A(_141_),
    .B(_100_),
    .C(_102_),
    .Y(_103_)
);

NOR2X1 _1598_ (
    .A(_695_),
    .B(_694_),
    .Y(_744_)
);

OAI21X1 _1178_ (
    .A(_355_),
    .B(SEL_A_8_bF$buf2),
    .C(_356_),
    .Y(_357_)
);

FILL FILL_11_0_0 (
);

FILL FILL_11_0_1 (
);

DFFPOSX1 _950_ (
    .Q(NIBBLES[2]),
    .CLK(CLK_bF$buf5),
    .D(_2_[2])
);

INVX1 _815_ (
    .A(DATA_B[26]),
    .Y(_9_)
);

NAND3X1 _1522_ (
    .A(_668_),
    .B(_670_),
    .C(_663_),
    .Y(_671_)
);

NAND3X1 _1102_ (
    .A(SEL_B[3]),
    .B(_281_),
    .C(_285_),
    .Y(_286_)
);

NAND3X1 _853_ (
    .A(_4_),
    .B(_43_),
    .C(_45_),
    .Y(_46_)
);

FILL FILL_8_0_0 (
);

FILL FILL_8_0_1 (
);

OR2X2 _909_ (
    .A(SEL_A_2_bF$buf0),
    .B(DATA_A[1]),
    .Y(_100_)
);

NAND2X1 _1331_ (
    .A(SEL_A_11_bF$buf4),
    .B(_502_),
    .Y(_503_)
);

NAND3X1 _1560_ (
    .A(_707_),
    .B(_706_),
    .C(_708_),
    .Y(_709_)
);

NAND3X1 _1140_ (
    .A(_457_),
    .B(_468_),
    .C(_477_),
    .Y(_478_)
);

NAND2X1 _891_ (
    .A(SEL_B_2_bF$buf4),
    .B(_82_),
    .Y(_83_)
);

FILL FILL_3_0_0 (
);

FILL FILL_3_0_1 (
);

DFFPOSX1 _1616_ (
    .Q(\nibble_mayor.nibble_C [3]),
    .CLK(CLK_bF$buf2),
    .D(_642_[3])
);

AOI21X1 _947_ (
    .A(_118_),
    .B(_137_),
    .C(_138_),
    .Y(_2_[1])
);

NAND3X1 _1425_ (
    .A(_616_),
    .B(_585_),
    .C(_594_),
    .Y(_595_)
);

NAND3X1 _1005_ (
    .A(_299_),
    .B(_186_),
    .C(_190_),
    .Y(_191_)
);

INVX1 _1234_ (
    .A(DATA_B[8]),
    .Y(_412_)
);

NAND3X1 _985_ (
    .A(_162_),
    .B(_167_),
    .C(_171_),
    .Y(_172_)
);

AND2X2 _1463_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLES[1]),
    .Y(_640_[1])
);

NAND3X1 _1043_ (
    .A(SEL_A[4]),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

INVX1 _794_ (
    .A(DATA_A[26]),
    .Y(_146_)
);

NAND2X1 _1519_ (
    .A(\nibble_mayor.nibble_B [2]),
    .B(_659_),
    .Y(_668_)
);

NAND3X1 _1272_ (
    .A(_322_),
    .B(_446_),
    .C(_448_),
    .Y(_449_)
);

AOI21X1 _1328_ (
    .A(_637_),
    .B(_500_),
    .C(_615_),
    .Y(_479_[2])
);

OR2X2 _1081_ (
    .A(SEL_A_5_bF$buf3),
    .B(DATA_A[9]),
    .Y(_265_)
);

AOI21X1 _1557_ (
    .A(_705_),
    .B(_704_),
    .C(_746_),
    .Y(_706_)
);

OAI21X1 _1137_ (
    .A(_473_),
    .B(SEL_A_8_bF$buf3),
    .C(_474_),
    .Y(_475_)
);

NAND3X1 _888_ (
    .A(_139_),
    .B(_70_),
    .C(_79_),
    .Y(_80_)
);

NAND3X1 _1366_ (
    .A(SEL_AB[3]),
    .B(_528_),
    .C(_537_),
    .Y(_538_)
);

NOR2X1 _1595_ (
    .A(_702_),
    .B(_701_),
    .Y(_742_)
);

NAND3X1 _1175_ (
    .A(_459_),
    .B(_351_),
    .C(_353_),
    .Y(_354_)
);

OR2X2 _1269_ (
    .A(SEL_B_8_bF$buf0),
    .B(DATA_B[1]),
    .Y(_446_)
);

INVX1 _812_ (
    .A(DATA_B[18]),
    .Y(_6_)
);

OAI21X1 _1498_ (
    .A(_645_),
    .B(_646_),
    .C(_639_[3]),
    .Y(_647_)
);

NAND3X1 _1078_ (
    .A(_300_),
    .B(_259_),
    .C(_261_),
    .Y(_262_)
);

OR2X2 _850_ (
    .A(SEL_B_2_bF$buf1),
    .B(DATA_B[7]),
    .Y(_43_)
);

NAND3X1 _906_ (
    .A(_3_),
    .B(_93_),
    .C(_97_),
    .Y(_98_)
);

DFFPOSX1 _1613_ (
    .Q(\nibble_mayor.nibble_C [0]),
    .CLK(CLK_bF$buf2),
    .D(_642_[0])
);

NAND2X1 _944_ (
    .A(SEL_B[1]),
    .B(_134_),
    .Y(_135_)
);

OAI21X1 _1422_ (
    .A(_590_),
    .B(SEL_A_11_bF$buf3),
    .C(_591_),
    .Y(_592_)
);

NAND2X1 _1002_ (
    .A(SEL_A_5_bF$buf4),
    .B(_187_),
    .Y(_188_)
);

INVX2 _809_ (
    .A(SEL_B[0]),
    .Y(_3_)
);

INVX1 _1231_ (
    .A(DATA_B[16]),
    .Y(_409_)
);

NAND2X1 _982_ (
    .A(SEL_B_5_bF$buf0),
    .B(_168_),
    .Y(_169_)
);

AND2X2 _1460_ (
    .A(RESET_L_bF$buf3),
    .B(NIBBLES[6]),
    .Y(_641_[2])
);

INVX1 _1040_ (
    .A(DATA_A[24]),
    .Y(_225_)
);

INVX1 _791_ (
    .A(DATA_A[18]),
    .Y(_143_)
);

NOR2X1 _1516_ (
    .A(\nibble_mayor.nibble_B [2]),
    .B(_659_),
    .Y(_665_)
);

NAND2X1 _847_ (
    .A(SEL_A[1]),
    .B(_39_),
    .Y(_40_)
);

NAND2X1 _1325_ (
    .A(SEL_B[10]),
    .B(_497_),
    .Y(_498_)
);

OAI21X1 _1554_ (
    .A(_701_),
    .B(_702_),
    .C(_700_),
    .Y(_703_)
);

NAND3X1 _1134_ (
    .A(_459_),
    .B(_469_),
    .C(_471_),
    .Y(_472_)
);

OAI21X1 _885_ (
    .A(_75_),
    .B(SEL_A_2_bF$buf2),
    .C(_76_),
    .Y(_77_)
);

OAI21X1 _1363_ (
    .A(_533_),
    .B(SEL_B_11_bF$buf4),
    .C(_534_),
    .Y(_535_)
);

NAND3X1 _1419_ (
    .A(_618_),
    .B(_586_),
    .C(_588_),
    .Y(_589_)
);

NAND2X1 _1592_ (
    .A(_721_),
    .B(_732_),
    .Y(_740_)
);

OR2X2 _1172_ (
    .A(SEL_A_8_bF$buf1),
    .B(DATA_A[7]),
    .Y(_351_)
);

NAND3X1 _1228_ (
    .A(SEL_B[7]),
    .B(_405_),
    .C(_404_),
    .Y(_406_)
);

NAND2X1 _979_ (
    .A(SEL_B_5_bF$buf4),
    .B(_165_),
    .Y(_166_)
);

AND2X2 _1457_ (
    .A(RESET_L_bF$buf0),
    .B(NIBBLES[11]),
    .Y(_642_[3])
);

INVX1 _1037_ (
    .A(DATA_A[16]),
    .Y(_222_)
);

INVX2 _788_ (
    .A(SEL_A[0]),
    .Y(_140_)
);

OR2X2 _1266_ (
    .A(SEL_B_8_bF$buf2),
    .B(DATA_B[13]),
    .Y(_443_)
);

NOR2X1 _1495_ (
    .A(\nibble_mayor.nibble_A [3]),
    .B(\nibble_mayor.nibble_B [3]),
    .Y(_645_)
);

OR2X2 _1075_ (
    .A(SEL_A_5_bF$buf4),
    .B(DATA_A[1]),
    .Y(_259_)
);

NAND2X1 _903_ (
    .A(SEL_B_2_bF$buf3),
    .B(DATA_B[24]),
    .Y(_95_)
);

OAI21X1 _1589_ (
    .A(_722_),
    .B(_648_),
    .C(_737_),
    .Y(_738_)
);

OR2X2 _1169_ (
    .A(SEL_A_8_bF$buf0),
    .B(DATA_A[11]),
    .Y(_348_)
);

NAND2X1 _1398_ (
    .A(SEL_B_11_bF$buf4),
    .B(_568_),
    .Y(_569_)
);

DFFPOSX1 _1610_ (
    .Q(\nibble_mayor.nibble_B [1]),
    .CLK(CLK_bF$buf3),
    .D(_641_[1])
);

INVX1 _941_ (
    .A(DATA_B[9]),
    .Y(_132_)
);

NAND2X1 _806_ (
    .A(SEL_A[1]),
    .B(_157_),
    .Y(_158_)
);

NAND2X1 _1513_ (
    .A(_654_),
    .B(_661_),
    .Y(_662_)
);

FILL FILL_10_1 (
);

INVX1 _844_ (
    .A(DATA_A[15]),
    .Y(_37_)
);

INVX1 _1322_ (
    .A(DATA_B[14]),
    .Y(_495_)
);

NAND3X1 _1551_ (
    .A(RESET_L_bF$buf1),
    .B(_698_),
    .C(_699_),
    .Y(_700_)
);

OR2X2 _1131_ (
    .A(SEL_A_8_bF$buf3),
    .B(DATA_A[6]),
    .Y(_469_)
);

NAND3X1 _882_ (
    .A(_141_),
    .B(_71_),
    .C(_73_),
    .Y(_74_)
);

DFFPOSX1 _1607_ (
    .Q(\nibble_mayor.nibble_A [2]),
    .CLK(CLK_bF$buf4),
    .D(_640_[2])
);

INVX1 _938_ (
    .A(DATA_B[17]),
    .Y(_129_)
);

NAND3X1 _1360_ (
    .A(_481_),
    .B(_529_),
    .C(_531_),
    .Y(_532_)
);

OR2X2 _1416_ (
    .A(SEL_A_11_bF$buf3),
    .B(DATA_A[5]),
    .Y(_586_)
);

INVX1 _1225_ (
    .A(DATA_B[28]),
    .Y(_403_)
);

INVX4 _976_ (
    .A(SEL_B[4]),
    .Y(_163_)
);

AND2X2 _1454_ (
    .A(RESET_L_bF$buf0),
    .B(NIBBLES[8]),
    .Y(_642_[0])
);

NAND3X1 _1034_ (
    .A(SEL_AB[1]),
    .B(_210_),
    .C(_219_),
    .Y(_220_)
);

DFFPOSX1 _785_ (
    .Q(_1_[3]),
    .CLK(CLK_bF$buf4),
    .D(_0_[3])
);

NAND3X1 _1263_ (
    .A(_322_),
    .B(_437_),
    .C(_439_),
    .Y(_440_)
);

INVX1 _1319_ (
    .A(DATA_B[22]),
    .Y(_492_)
);

NAND2X1 _1492_ (
    .A(_757_),
    .B(_771_),
    .Y(_772_)
);

NAND3X1 _1072_ (
    .A(_162_),
    .B(_252_),
    .C(_256_),
    .Y(_257_)
);

AOI21X1 _1548_ (
    .A(_696_),
    .B(_690_),
    .C(_648_),
    .Y(_697_)
);

OR2X2 _1128_ (
    .A(SEL_A_8_bF$buf2),
    .B(DATA_A[10]),
    .Y(_466_)
);

OR2X2 _879_ (
    .A(SEL_A_2_bF$buf2),
    .B(DATA_A[4]),
    .Y(_71_)
);

OR2X2 _1357_ (
    .A(SEL_B_11_bF$buf4),
    .B(DATA_B[3]),
    .Y(_529_)
);

NAND2X1 _900_ (
    .A(SEL_B_2_bF$buf3),
    .B(_91_),
    .Y(_92_)
);

NOR2X1 _1586_ (
    .A(_716_),
    .B(_733_),
    .Y(_735_)
);

NAND3X1 _1166_ (
    .A(_459_),
    .B(_342_),
    .C(_344_),
    .Y(_345_)
);

NAND3X1 _1395_ (
    .A(SEL_B[9]),
    .B(_561_),
    .C(_565_),
    .Y(_566_)
);

INVX1 _803_ (
    .A(DATA_A[14]),
    .Y(_155_)
);

NAND2X1 _1489_ (
    .A(_756_),
    .B(_755_),
    .Y(_769_)
);

NAND2X1 _1069_ (
    .A(SEL_B_5_bF$buf0),
    .B(DATA_B[24]),
    .Y(_254_)
);

INVX1 _1298_ (
    .A(DATA_A[22]),
    .Y(_629_)
);

INVX2 _1510_ (
    .A(\nibble_mayor.nibble_A [2]),
    .Y(_659_)
);

INVX1 _841_ (
    .A(DATA_A[23]),
    .Y(_34_)
);

DFFPOSX1 _1604_ (
    .Q(NIBBLE_MAYOR[3]),
    .CLK(CLK_bF$buf5),
    .D(_639_[3])
);

NAND3X1 _935_ (
    .A(SEL_B[1]),
    .B(_125_),
    .C(_124_),
    .Y(_126_)
);

OR2X2 _1413_ (
    .A(SEL_A_11_bF$buf0),
    .B(DATA_A[9]),
    .Y(_583_)
);

INVX1 _1222_ (
    .A(DATA_B[20]),
    .Y(_400_)
);

NAND3X1 _973_ (
    .A(SEL_A[3]),
    .B(_313_),
    .C(_317_),
    .Y(_318_)
);

AND2X2 _1451_ (
    .A(RESET_L_bF$buf4),
    .B(NIBBLES[13]),
    .Y(_643_[1])
);

OAI21X1 _1031_ (
    .A(_215_),
    .B(SEL_B_5_bF$buf1),
    .C(_216_),
    .Y(_217_)
);

DFFPOSX1 _782_ (
    .Q(_1_[0]),
    .CLK(CLK_bF$buf2),
    .D(_0_[0])
);

INVX1 _1507_ (
    .A(\nibble_mayor.nibble_B [0]),
    .Y(_656_)
);

NAND3X1 _838_ (
    .A(SEL_A[1]),
    .B(_30_),
    .C(_29_),
    .Y(_31_)
);

OR2X2 _1260_ (
    .A(SEL_B_8_bF$buf2),
    .B(DATA_B[5]),
    .Y(_437_)
);

NAND3X1 _1316_ (
    .A(SEL_B[10]),
    .B(_488_),
    .C(_487_),
    .Y(_489_)
);

NOR2X1 _1545_ (
    .A(\nibble_mayor.nibble_C [2]),
    .B(_644_),
    .Y(_694_)
);

NAND3X1 _1125_ (
    .A(_459_),
    .B(_460_),
    .C(_462_),
    .Y(_463_)
);

OR2X2 _876_ (
    .A(SEL_A_2_bF$buf4),
    .B(DATA_A[8]),
    .Y(_68_)
);

OR2X2 _1354_ (
    .A(SEL_B_11_bF$buf1),
    .B(DATA_B[15]),
    .Y(_526_)
);

OAI21X1 _1583_ (
    .A(_731_),
    .B(_724_),
    .C(_727_),
    .Y(_732_)
);

OR2X2 _1163_ (
    .A(DATA_A[3]),
    .B(SEL_A_8_bF$buf2),
    .Y(_342_)
);

NAND3X1 _1219_ (
    .A(SEL_A[6]),
    .B(_392_),
    .C(_396_),
    .Y(_397_)
);

NAND2X1 _1392_ (
    .A(SEL_B_11_bF$buf0),
    .B(_562_),
    .Y(_563_)
);

DFFPOSX1 _1448_ (
    .Q(NIBBLES[14]),
    .CLK(CLK_bF$buf0),
    .D(_479_[2])
);

NAND3X1 _1028_ (
    .A(_163_),
    .B(_211_),
    .C(_213_),
    .Y(_214_)
);

BUFX2 _779_ (
    .A(_1_[1]),
    .Y(DATA_OUT[1])
);

endmodule
