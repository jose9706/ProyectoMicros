VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO nibble_top
   CLASS BLOCK ;
   FOREIGN nibble_top ;
   ORIGIN 2.6000 3.0000 ;
   SIZE 178.8000 BY 167.2000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.2000 160.2000 173.4000 160.8000 ;
	    RECT 0.6000 157.9000 1.0000 160.2000 ;
	    RECT 2.2000 157.9000 2.6000 160.2000 ;
	    RECT 3.8000 157.9000 4.2000 160.2000 ;
	    RECT 4.6000 157.9000 5.0000 160.2000 ;
	    RECT 6.2000 157.9000 6.6000 160.2000 ;
	    RECT 7.8000 157.9000 8.2000 160.2000 ;
	    RECT 8.6000 155.9000 9.0000 160.2000 ;
	    RECT 10.7000 157.9000 11.1000 160.2000 ;
	    RECT 11.8000 157.9000 12.2000 160.2000 ;
	    RECT 13.4000 157.9000 13.8000 160.2000 ;
	    RECT 14.2000 157.9000 14.6000 160.2000 ;
	    RECT 15.8000 157.9000 16.2000 160.2000 ;
	    RECT 17.4000 156.5000 17.8000 160.2000 ;
	    RECT 19.0000 157.9000 19.4000 160.2000 ;
	    RECT 20.6000 157.9000 21.0000 160.2000 ;
	    RECT 21.4000 157.9000 21.8000 160.2000 ;
	    RECT 23.0000 157.9000 23.4000 160.2000 ;
	    RECT 24.6000 157.9000 25.0000 160.2000 ;
	    RECT 25.4000 157.9000 25.8000 160.2000 ;
	    RECT 27.0000 157.9000 27.4000 160.2000 ;
	    RECT 27.8000 157.9000 28.2000 160.2000 ;
	    RECT 30.2000 157.9000 30.6000 160.2000 ;
	    RECT 31.0000 157.9000 31.4000 160.2000 ;
	    RECT 32.6000 155.9000 33.0000 160.2000 ;
	    RECT 34.7000 157.9000 35.1000 160.2000 ;
	    RECT 35.8000 157.9000 36.2000 160.2000 ;
	    RECT 37.4000 157.9000 37.8000 160.2000 ;
	    RECT 38.2000 157.9000 38.6000 160.2000 ;
	    RECT 39.8000 157.9000 40.2000 160.2000 ;
	    RECT 41.4000 156.5000 41.8000 160.2000 ;
	    RECT 43.0000 157.9000 43.4000 160.2000 ;
	    RECT 44.6000 157.9000 45.0000 160.2000 ;
	    RECT 45.4000 157.9000 45.8000 160.2000 ;
	    RECT 47.0000 157.9000 47.4000 160.2000 ;
	    RECT 48.6000 157.9000 49.0000 160.2000 ;
	    RECT 49.4000 157.9000 49.8000 160.2000 ;
	    RECT 51.0000 157.9000 51.4000 160.2000 ;
	    RECT 51.8000 157.9000 52.2000 160.2000 ;
	    RECT 53.4000 157.9000 53.8000 160.2000 ;
	    RECT 55.0000 156.5000 55.4000 160.2000 ;
	    RECT 56.6000 157.9000 57.0000 160.2000 ;
	    RECT 58.2000 155.9000 58.6000 160.2000 ;
	    RECT 60.3000 157.9000 60.7000 160.2000 ;
	    RECT 63.0000 157.9000 63.4000 160.2000 ;
	    RECT 64.6000 157.9000 65.0000 160.2000 ;
	    RECT 65.4000 157.9000 65.8000 160.2000 ;
	    RECT 67.0000 157.9000 67.4000 160.2000 ;
	    RECT 68.6000 157.9000 69.0000 160.2000 ;
	    RECT 69.4000 157.9000 69.8000 160.2000 ;
	    RECT 71.0000 157.9000 71.4000 160.2000 ;
	    RECT 71.8000 157.9000 72.2000 160.2000 ;
	    RECT 73.4000 157.9000 73.8000 160.2000 ;
	    RECT 75.0000 157.9000 75.4000 160.2000 ;
	    RECT 77.4000 155.9000 77.8000 160.2000 ;
	    RECT 78.2000 157.9000 78.6000 160.2000 ;
	    RECT 79.8000 157.9000 80.2000 160.2000 ;
	    RECT 81.4000 155.9000 81.8000 160.2000 ;
	    RECT 84.2000 157.9000 84.6000 160.2000 ;
	    RECT 85.8000 157.9000 86.2000 160.2000 ;
	    RECT 88.6000 156.0000 89.0000 160.2000 ;
	    RECT 91.0000 155.9000 91.4000 160.2000 ;
	    RECT 91.8000 155.9000 92.2000 160.2000 ;
	    RECT 95.0000 155.9000 95.4000 160.2000 ;
	    RECT 95.8000 155.9000 96.2000 160.2000 ;
	    RECT 99.0000 155.9000 99.4000 160.2000 ;
	    RECT 101.4000 155.9000 101.8000 160.2000 ;
	    RECT 102.2000 157.9000 102.6000 160.2000 ;
	    RECT 103.8000 157.9000 104.2000 160.2000 ;
	    RECT 106.2000 156.5000 106.6000 160.2000 ;
	    RECT 107.8000 157.9000 108.2000 160.2000 ;
	    RECT 109.4000 157.9000 109.8000 160.2000 ;
	    RECT 111.8000 155.9000 112.2000 160.2000 ;
	    RECT 114.2000 157.9000 114.6000 160.2000 ;
	    RECT 115.8000 157.9000 116.2000 160.2000 ;
	    RECT 117.4000 157.9000 117.8000 160.2000 ;
	    RECT 119.0000 156.5000 119.4000 160.2000 ;
	    RECT 123.0000 156.9000 123.4000 160.2000 ;
	    RECT 128.6000 157.9000 129.0000 160.2000 ;
	    RECT 130.5000 157.9000 130.9000 160.2000 ;
	    RECT 132.6000 155.9000 133.0000 160.2000 ;
	    RECT 135.0000 156.5000 135.4000 160.2000 ;
	    RECT 136.9000 157.9000 137.3000 160.2000 ;
	    RECT 139.0000 155.9000 139.4000 160.2000 ;
	    RECT 141.4000 155.9000 141.8000 160.2000 ;
	    RECT 143.8000 156.5000 144.2000 160.2000 ;
	    RECT 145.4000 157.9000 145.8000 160.2000 ;
	    RECT 147.0000 157.9000 147.4000 160.2000 ;
	    RECT 147.8000 157.9000 148.2000 160.2000 ;
	    RECT 149.4000 158.1000 149.8000 160.2000 ;
	    RECT 151.8000 158.1000 152.2000 160.2000 ;
	    RECT 153.4000 157.9000 153.8000 160.2000 ;
	    RECT 154.2000 157.9000 154.6000 160.2000 ;
	    RECT 155.8000 157.9000 156.2000 160.2000 ;
	    RECT 156.6000 155.9000 157.0000 160.2000 ;
	    RECT 158.7000 157.9000 159.1000 160.2000 ;
	    RECT 159.8000 157.9000 160.2000 160.2000 ;
	    RECT 161.4000 157.9000 161.8000 160.2000 ;
	    RECT 163.0000 156.0000 163.4000 160.2000 ;
	    RECT 165.8000 157.9000 166.2000 160.2000 ;
	    RECT 167.4000 157.9000 167.8000 160.2000 ;
	    RECT 170.2000 155.9000 170.6000 160.2000 ;
	    RECT 1.4000 140.8000 1.8000 142.9000 ;
	    RECT 3.0000 140.8000 3.4000 143.1000 ;
	    RECT 4.9000 140.8000 5.3000 145.1000 ;
	    RECT 7.3000 140.8000 7.7000 143.1000 ;
	    RECT 9.4000 140.8000 9.8000 145.1000 ;
	    RECT 11.0000 140.8000 11.4000 143.1000 ;
	    RECT 12.6000 140.8000 13.0000 144.5000 ;
	    RECT 14.5000 140.8000 14.9000 143.1000 ;
	    RECT 16.6000 140.8000 17.0000 145.1000 ;
	    RECT 18.2000 140.8000 18.6000 143.1000 ;
	    RECT 19.8000 140.8000 20.2000 143.1000 ;
	    RECT 20.6000 140.8000 21.0000 143.1000 ;
	    RECT 22.2000 140.8000 22.6000 142.9000 ;
	    RECT 24.9000 140.8000 25.3000 145.1000 ;
	    RECT 27.3000 140.8000 27.7000 143.1000 ;
	    RECT 29.4000 140.8000 29.8000 145.1000 ;
	    RECT 31.0000 140.8000 31.4000 143.1000 ;
	    RECT 32.1000 140.8000 32.5000 143.1000 ;
	    RECT 34.2000 140.8000 34.6000 145.1000 ;
	    RECT 35.8000 140.8000 36.2000 143.1000 ;
	    RECT 36.6000 140.8000 37.0000 145.1000 ;
	    RECT 38.7000 140.8000 39.1000 143.1000 ;
	    RECT 40.6000 140.8000 41.0000 144.5000 ;
	    RECT 42.2000 140.8000 42.6000 143.1000 ;
	    RECT 43.8000 140.8000 44.2000 145.1000 ;
	    RECT 45.9000 140.8000 46.3000 143.1000 ;
	    RECT 48.3000 140.8000 48.7000 145.1000 ;
	    RECT 50.2000 140.8000 50.6000 143.1000 ;
	    RECT 52.6000 140.8000 53.0000 142.9000 ;
	    RECT 54.2000 140.8000 54.6000 143.1000 ;
	    RECT 55.0000 140.8000 55.4000 143.1000 ;
	    RECT 57.4000 140.8000 57.8000 142.9000 ;
	    RECT 59.0000 140.8000 59.4000 143.1000 ;
	    RECT 62.7000 140.8000 63.1000 145.1000 ;
	    RECT 64.6000 140.8000 65.0000 143.1000 ;
	    RECT 66.2000 140.8000 66.6000 142.9000 ;
	    RECT 67.8000 140.8000 68.2000 143.1000 ;
	    RECT 69.4000 140.8000 69.8000 142.9000 ;
	    RECT 71.0000 140.8000 71.4000 143.1000 ;
	    RECT 73.4000 140.8000 73.8000 144.5000 ;
	    RECT 75.8000 140.8000 76.2000 145.1000 ;
	    RECT 78.2000 140.8000 78.6000 143.1000 ;
	    RECT 79.8000 140.8000 80.2000 143.1000 ;
	    RECT 80.6000 140.8000 81.0000 143.1000 ;
	    RECT 82.2000 140.8000 82.6000 142.9000 ;
	    RECT 83.8000 140.8000 84.2000 143.1000 ;
	    RECT 85.4000 140.8000 85.8000 145.1000 ;
	    RECT 87.8000 140.8000 88.2000 144.5000 ;
	    RECT 91.8000 140.8000 92.2000 145.1000 ;
	    RECT 93.4000 140.8000 93.8000 142.9000 ;
	    RECT 95.0000 140.8000 95.4000 143.1000 ;
	    RECT 95.8000 140.8000 96.2000 143.1000 ;
	    RECT 97.4000 140.8000 97.8000 143.1000 ;
	    RECT 99.8000 140.8000 100.2000 145.1000 ;
	    RECT 101.4000 140.8000 101.8000 142.9000 ;
	    RECT 103.0000 140.8000 103.4000 143.1000 ;
	    RECT 103.8000 140.8000 104.2000 145.1000 ;
	    RECT 105.4000 140.8000 105.8000 145.1000 ;
	    RECT 106.5000 140.8000 106.9000 143.1000 ;
	    RECT 108.6000 140.8000 109.0000 145.1000 ;
	    RECT 109.7000 140.8000 110.1000 143.1000 ;
	    RECT 111.8000 140.8000 112.2000 145.1000 ;
	    RECT 115.0000 140.8000 115.4000 142.9000 ;
	    RECT 116.6000 140.8000 117.0000 143.1000 ;
	    RECT 117.4000 140.8000 117.8000 145.1000 ;
	    RECT 119.5000 140.8000 119.9000 143.1000 ;
	    RECT 120.9000 140.8000 121.3000 143.1000 ;
	    RECT 123.0000 140.8000 123.4000 145.1000 ;
	    RECT 123.8000 140.8000 124.2000 143.1000 ;
	    RECT 125.4000 140.8000 125.8000 142.9000 ;
	    RECT 128.6000 140.8000 129.0000 144.5000 ;
	    RECT 130.5000 140.8000 130.9000 143.1000 ;
	    RECT 132.6000 140.8000 133.0000 145.1000 ;
	    RECT 138.2000 140.8000 138.6000 144.1000 ;
	    RECT 139.8000 140.8000 140.2000 145.1000 ;
	    RECT 141.9000 140.8000 142.3000 143.1000 ;
	    RECT 145.4000 140.8000 145.8000 144.5000 ;
	    RECT 149.4000 140.8000 149.8000 144.5000 ;
	    RECT 151.0000 140.8000 151.4000 145.1000 ;
	    RECT 153.4000 140.8000 153.8000 143.1000 ;
	    RECT 155.0000 140.8000 155.4000 142.9000 ;
	    RECT 156.6000 140.8000 157.0000 145.1000 ;
	    RECT 158.7000 140.8000 159.1000 143.1000 ;
	    RECT 159.8000 140.8000 160.2000 145.1000 ;
	    RECT 163.0000 140.8000 163.4000 145.0000 ;
	    RECT 165.8000 140.8000 166.2000 143.1000 ;
	    RECT 167.4000 140.8000 167.8000 143.1000 ;
	    RECT 170.2000 140.8000 170.6000 145.1000 ;
	    RECT 0.2000 140.2000 173.4000 140.8000 ;
	    RECT 1.4000 136.5000 1.8000 140.2000 ;
	    RECT 3.0000 137.9000 3.4000 140.2000 ;
	    RECT 4.6000 137.9000 5.0000 140.2000 ;
	    RECT 6.7000 135.9000 7.1000 140.2000 ;
	    RECT 8.6000 137.9000 9.0000 140.2000 ;
	    RECT 10.2000 138.1000 10.6000 140.2000 ;
	    RECT 11.8000 137.9000 12.2000 140.2000 ;
	    RECT 13.4000 137.9000 13.8000 140.2000 ;
	    RECT 14.2000 137.9000 14.6000 140.2000 ;
	    RECT 15.8000 137.9000 16.2000 140.2000 ;
	    RECT 16.6000 137.9000 17.0000 140.2000 ;
	    RECT 18.2000 137.9000 18.6000 140.2000 ;
	    RECT 19.0000 137.9000 19.4000 140.2000 ;
	    RECT 20.6000 137.9000 21.0000 140.2000 ;
	    RECT 21.4000 137.9000 21.8000 140.2000 ;
	    RECT 23.0000 137.9000 23.4000 140.2000 ;
	    RECT 24.6000 136.5000 25.0000 140.2000 ;
	    RECT 27.0000 137.9000 27.4000 140.2000 ;
	    RECT 27.8000 137.9000 28.2000 140.2000 ;
	    RECT 29.4000 137.9000 29.8000 140.2000 ;
	    RECT 30.2000 137.9000 30.6000 140.2000 ;
	    RECT 31.8000 137.9000 32.2000 140.2000 ;
	    RECT 33.9000 135.9000 34.3000 140.2000 ;
	    RECT 35.8000 137.9000 36.2000 140.2000 ;
	    RECT 37.4000 137.9000 37.8000 140.2000 ;
	    RECT 38.2000 137.9000 38.6000 140.2000 ;
	    RECT 39.8000 135.9000 40.2000 140.2000 ;
	    RECT 41.9000 137.9000 42.3000 140.2000 ;
	    RECT 43.0000 137.9000 43.4000 140.2000 ;
	    RECT 44.6000 137.9000 45.0000 140.2000 ;
	    RECT 45.4000 137.9000 45.8000 140.2000 ;
	    RECT 47.0000 135.9000 47.4000 140.2000 ;
	    RECT 49.1000 137.9000 49.5000 140.2000 ;
	    RECT 50.2000 137.9000 50.6000 140.2000 ;
	    RECT 51.8000 137.9000 52.2000 140.2000 ;
	    RECT 52.6000 137.9000 53.0000 140.2000 ;
	    RECT 54.2000 137.9000 54.6000 140.2000 ;
	    RECT 55.3000 137.9000 55.7000 140.2000 ;
	    RECT 57.4000 135.9000 57.8000 140.2000 ;
	    RECT 58.2000 137.9000 58.6000 140.2000 ;
	    RECT 59.8000 137.9000 60.2000 140.2000 ;
	    RECT 62.2000 137.9000 62.6000 140.2000 ;
	    RECT 63.8000 137.9000 64.2000 140.2000 ;
	    RECT 65.9000 135.9000 66.3000 140.2000 ;
	    RECT 67.8000 137.9000 68.2000 140.2000 ;
	    RECT 69.4000 137.9000 69.8000 140.2000 ;
	    RECT 70.2000 137.9000 70.6000 140.2000 ;
	    RECT 71.8000 137.9000 72.2000 140.2000 ;
	    RECT 73.9000 135.9000 74.3000 140.2000 ;
	    RECT 76.6000 138.1000 77.0000 140.2000 ;
	    RECT 78.2000 137.9000 78.6000 140.2000 ;
	    RECT 79.0000 137.9000 79.4000 140.2000 ;
	    RECT 80.6000 137.9000 81.0000 140.2000 ;
	    RECT 81.7000 137.9000 82.1000 140.2000 ;
	    RECT 83.8000 135.9000 84.2000 140.2000 ;
	    RECT 84.6000 135.9000 85.0000 140.2000 ;
	    RECT 87.0000 135.9000 87.4000 140.2000 ;
	    RECT 89.1000 137.9000 89.5000 140.2000 ;
	    RECT 90.2000 135.9000 90.6000 140.2000 ;
	    RECT 91.8000 137.9000 92.2000 140.2000 ;
	    RECT 93.4000 138.1000 93.8000 140.2000 ;
	    RECT 95.0000 137.9000 95.4000 140.2000 ;
	    RECT 96.6000 138.1000 97.0000 140.2000 ;
	    RECT 99.0000 138.1000 99.4000 140.2000 ;
	    RECT 100.6000 137.9000 101.0000 140.2000 ;
	    RECT 102.2000 138.1000 102.6000 140.2000 ;
	    RECT 103.8000 137.9000 104.2000 140.2000 ;
	    RECT 104.6000 137.9000 105.0000 140.2000 ;
	    RECT 107.8000 135.9000 108.2000 140.2000 ;
	    RECT 109.4000 136.5000 109.8000 140.2000 ;
	    RECT 115.0000 136.5000 115.4000 140.2000 ;
	    RECT 116.6000 135.9000 117.0000 140.2000 ;
	    RECT 119.8000 137.9000 120.2000 140.2000 ;
	    RECT 121.4000 137.9000 121.8000 140.2000 ;
	    RECT 122.2000 137.9000 122.6000 140.2000 ;
	    RECT 123.8000 137.9000 124.2000 140.2000 ;
	    RECT 124.6000 137.9000 125.0000 140.2000 ;
	    RECT 126.2000 138.1000 126.6000 140.2000 ;
	    RECT 127.8000 135.9000 128.2000 140.2000 ;
	    RECT 129.9000 137.9000 130.3000 140.2000 ;
	    RECT 131.0000 135.9000 131.4000 140.2000 ;
	    RECT 133.4000 135.9000 133.8000 140.2000 ;
	    RECT 136.6000 135.9000 137.0000 140.2000 ;
	    RECT 137.7000 137.9000 138.1000 140.2000 ;
	    RECT 139.8000 135.9000 140.2000 140.2000 ;
	    RECT 140.9000 137.9000 141.3000 140.2000 ;
	    RECT 143.0000 135.9000 143.4000 140.2000 ;
	    RECT 145.4000 135.9000 145.8000 140.2000 ;
	    RECT 147.0000 138.1000 147.4000 140.2000 ;
	    RECT 148.6000 137.9000 149.0000 140.2000 ;
	    RECT 149.4000 137.9000 149.8000 140.2000 ;
	    RECT 151.0000 137.9000 151.4000 140.2000 ;
	    RECT 152.1000 137.9000 152.5000 140.2000 ;
	    RECT 154.2000 135.9000 154.6000 140.2000 ;
	    RECT 155.8000 136.1000 156.2000 140.2000 ;
	    RECT 157.4000 137.9000 157.8000 140.2000 ;
	    RECT 158.2000 137.9000 158.6000 140.2000 ;
	    RECT 159.8000 138.1000 160.2000 140.2000 ;
	    RECT 161.4000 137.9000 161.8000 140.2000 ;
	    RECT 164.6000 136.5000 165.0000 140.2000 ;
	    RECT 166.2000 135.9000 166.6000 140.2000 ;
	    RECT 168.3000 137.9000 168.7000 140.2000 ;
	    RECT 169.4000 135.9000 169.8000 140.2000 ;
	    RECT 171.5000 137.9000 171.9000 140.2000 ;
	    RECT 0.6000 120.8000 1.0000 125.1000 ;
	    RECT 2.2000 120.8000 2.6000 125.1000 ;
	    RECT 3.8000 120.8000 4.2000 122.9000 ;
	    RECT 5.4000 120.8000 5.8000 123.1000 ;
	    RECT 6.2000 120.8000 6.6000 125.1000 ;
	    RECT 7.8000 120.8000 8.2000 125.1000 ;
	    RECT 8.6000 120.8000 9.0000 123.1000 ;
	    RECT 10.2000 120.8000 10.6000 122.9000 ;
	    RECT 11.8000 120.8000 12.2000 123.1000 ;
	    RECT 13.4000 120.8000 13.8000 122.9000 ;
	    RECT 15.8000 120.8000 16.2000 122.9000 ;
	    RECT 17.4000 120.8000 17.8000 123.1000 ;
	    RECT 19.0000 120.8000 19.4000 122.9000 ;
	    RECT 20.6000 120.8000 21.0000 123.1000 ;
	    RECT 22.5000 120.8000 22.9000 125.1000 ;
	    RECT 25.9000 120.8000 26.3000 125.1000 ;
	    RECT 28.6000 120.8000 29.0000 122.9000 ;
	    RECT 30.2000 120.8000 30.6000 123.1000 ;
	    RECT 31.8000 120.8000 32.2000 122.9000 ;
	    RECT 33.4000 120.8000 33.8000 123.1000 ;
	    RECT 34.2000 120.8000 34.6000 123.1000 ;
	    RECT 35.8000 120.8000 36.2000 122.9000 ;
	    RECT 37.4000 120.8000 37.8000 123.1000 ;
	    RECT 39.0000 120.8000 39.4000 123.1000 ;
	    RECT 40.6000 120.8000 41.0000 123.1000 ;
	    RECT 41.4000 120.8000 41.8000 123.1000 ;
	    RECT 43.0000 120.8000 43.4000 123.1000 ;
	    RECT 45.1000 120.8000 45.5000 125.1000 ;
	    RECT 47.8000 120.8000 48.2000 122.9000 ;
	    RECT 49.4000 120.8000 49.8000 123.1000 ;
	    RECT 51.5000 120.8000 51.9000 125.1000 ;
	    RECT 54.2000 120.8000 54.6000 122.9000 ;
	    RECT 55.8000 120.8000 56.2000 123.1000 ;
	    RECT 57.4000 120.8000 57.8000 124.5000 ;
	    RECT 61.4000 120.8000 61.8000 122.9000 ;
	    RECT 63.0000 120.8000 63.4000 123.1000 ;
	    RECT 65.1000 120.8000 65.5000 125.1000 ;
	    RECT 67.0000 120.8000 67.4000 123.1000 ;
	    RECT 68.6000 120.8000 69.0000 122.9000 ;
	    RECT 70.2000 120.8000 70.6000 123.1000 ;
	    RECT 71.8000 120.8000 72.2000 122.9000 ;
	    RECT 73.4000 120.8000 73.8000 123.1000 ;
	    RECT 75.0000 120.8000 75.4000 123.1000 ;
	    RECT 76.6000 120.8000 77.0000 123.1000 ;
	    RECT 77.4000 120.8000 77.8000 123.1000 ;
	    RECT 79.0000 120.8000 79.4000 122.9000 ;
	    RECT 80.6000 120.8000 81.0000 125.1000 ;
	    RECT 82.2000 120.8000 82.6000 125.1000 ;
	    RECT 83.0000 120.8000 83.4000 123.1000 ;
	    RECT 84.6000 120.8000 85.0000 123.1000 ;
	    RECT 86.2000 120.8000 86.6000 125.1000 ;
	    RECT 89.0000 120.8000 89.4000 123.1000 ;
	    RECT 90.6000 120.8000 91.0000 123.1000 ;
	    RECT 93.4000 120.8000 93.8000 125.0000 ;
	    RECT 95.0000 120.8000 95.4000 123.1000 ;
	    RECT 96.6000 120.8000 97.0000 123.1000 ;
	    RECT 98.2000 120.8000 98.6000 123.1000 ;
	    RECT 99.0000 120.8000 99.4000 123.1000 ;
	    RECT 100.6000 120.8000 101.0000 123.1000 ;
	    RECT 101.4000 120.8000 101.8000 123.1000 ;
	    RECT 103.0000 120.8000 103.4000 123.1000 ;
	    RECT 104.6000 120.8000 105.0000 125.1000 ;
	    RECT 107.4000 120.8000 107.8000 123.1000 ;
	    RECT 109.0000 120.8000 109.4000 123.1000 ;
	    RECT 111.8000 120.8000 112.2000 125.0000 ;
	    RECT 115.0000 120.8000 115.4000 123.1000 ;
	    RECT 116.6000 120.8000 117.0000 123.1000 ;
	    RECT 117.4000 120.8000 117.8000 123.1000 ;
	    RECT 119.8000 120.8000 120.2000 124.9000 ;
	    RECT 121.4000 120.8000 121.8000 123.1000 ;
	    RECT 123.0000 120.8000 123.4000 124.5000 ;
	    RECT 124.9000 120.8000 125.3000 123.1000 ;
	    RECT 127.0000 120.8000 127.4000 125.1000 ;
	    RECT 128.6000 120.8000 129.0000 124.5000 ;
	    RECT 132.6000 120.8000 133.0000 124.5000 ;
	    RECT 135.8000 120.8000 136.2000 125.1000 ;
	    RECT 137.4000 120.8000 137.8000 123.1000 ;
	    RECT 138.2000 120.8000 138.6000 123.1000 ;
	    RECT 139.8000 120.8000 140.2000 123.1000 ;
	    RECT 141.4000 120.8000 141.8000 124.5000 ;
	    RECT 144.6000 120.8000 145.0000 123.1000 ;
	    RECT 146.2000 120.8000 146.6000 123.1000 ;
	    RECT 148.6000 120.8000 149.0000 124.5000 ;
	    RECT 150.2000 120.8000 150.6000 123.1000 ;
	    RECT 151.8000 120.8000 152.2000 123.1000 ;
	    RECT 153.4000 120.8000 153.8000 124.5000 ;
	    RECT 156.6000 120.8000 157.0000 123.1000 ;
	    RECT 158.2000 120.8000 158.6000 123.1000 ;
	    RECT 159.0000 120.8000 159.4000 123.1000 ;
	    RECT 160.6000 120.8000 161.0000 123.1000 ;
	    RECT 161.4000 120.8000 161.8000 123.1000 ;
	    RECT 163.0000 120.8000 163.4000 123.1000 ;
	    RECT 164.6000 120.8000 165.0000 125.0000 ;
	    RECT 167.4000 120.8000 167.8000 123.1000 ;
	    RECT 169.0000 120.8000 169.4000 123.1000 ;
	    RECT 171.8000 120.8000 172.2000 125.1000 ;
	    RECT 0.2000 120.2000 173.4000 120.8000 ;
	    RECT 1.9000 115.9000 2.3000 120.2000 ;
	    RECT 3.8000 117.9000 4.2000 120.2000 ;
	    RECT 5.4000 117.9000 5.8000 120.2000 ;
	    RECT 7.0000 117.9000 7.4000 120.2000 ;
	    RECT 7.8000 117.9000 8.2000 120.2000 ;
	    RECT 9.4000 117.9000 9.8000 120.2000 ;
	    RECT 11.0000 117.9000 11.4000 120.2000 ;
	    RECT 12.6000 118.1000 13.0000 120.2000 ;
	    RECT 14.2000 117.9000 14.6000 120.2000 ;
	    RECT 16.1000 115.9000 16.5000 120.2000 ;
	    RECT 19.0000 116.5000 19.4000 120.2000 ;
	    RECT 20.6000 117.9000 21.0000 120.2000 ;
	    RECT 22.2000 117.9000 22.6000 120.2000 ;
	    RECT 23.8000 117.9000 24.2000 120.2000 ;
	    RECT 25.9000 115.9000 26.3000 120.2000 ;
	    RECT 27.8000 117.9000 28.2000 120.2000 ;
	    RECT 29.4000 118.1000 29.8000 120.2000 ;
	    RECT 31.0000 117.9000 31.4000 120.2000 ;
	    RECT 32.6000 117.9000 33.0000 120.2000 ;
	    RECT 34.2000 117.9000 34.6000 120.2000 ;
	    RECT 35.8000 118.1000 36.2000 120.2000 ;
	    RECT 37.4000 117.9000 37.8000 120.2000 ;
	    RECT 39.0000 117.9000 39.4000 120.2000 ;
	    RECT 40.6000 116.5000 41.0000 120.2000 ;
	    RECT 43.5000 115.9000 43.9000 120.2000 ;
	    RECT 46.2000 118.1000 46.6000 120.2000 ;
	    RECT 47.8000 117.9000 48.2000 120.2000 ;
	    RECT 49.9000 115.9000 50.3000 120.2000 ;
	    RECT 51.8000 117.9000 52.2000 120.2000 ;
	    RECT 53.4000 117.9000 53.8000 120.2000 ;
	    RECT 55.0000 117.9000 55.4000 120.2000 ;
	    RECT 55.8000 117.9000 56.2000 120.2000 ;
	    RECT 57.4000 118.1000 57.8000 120.2000 ;
	    RECT 59.8000 116.5000 60.2000 120.2000 ;
	    RECT 63.8000 116.5000 64.2000 120.2000 ;
	    RECT 66.2000 118.1000 66.6000 120.2000 ;
	    RECT 67.8000 117.9000 68.2000 120.2000 ;
	    RECT 69.4000 118.1000 69.8000 120.2000 ;
	    RECT 71.0000 117.9000 71.4000 120.2000 ;
	    RECT 72.6000 115.9000 73.0000 120.2000 ;
	    RECT 75.4000 117.9000 75.8000 120.2000 ;
	    RECT 77.0000 117.9000 77.4000 120.2000 ;
	    RECT 79.8000 116.0000 80.2000 120.2000 ;
	    RECT 82.2000 116.0000 82.6000 120.2000 ;
	    RECT 85.0000 117.9000 85.4000 120.2000 ;
	    RECT 86.6000 117.9000 87.0000 120.2000 ;
	    RECT 89.4000 115.9000 89.8000 120.2000 ;
	    RECT 91.8000 115.9000 92.2000 120.2000 ;
	    RECT 94.6000 117.9000 95.0000 120.2000 ;
	    RECT 96.2000 117.9000 96.6000 120.2000 ;
	    RECT 99.0000 116.0000 99.4000 120.2000 ;
	    RECT 101.4000 115.9000 101.8000 120.2000 ;
	    RECT 104.2000 117.9000 104.6000 120.2000 ;
	    RECT 105.8000 117.9000 106.2000 120.2000 ;
	    RECT 108.6000 116.0000 109.0000 120.2000 ;
	    RECT 112.6000 116.0000 113.0000 120.2000 ;
	    RECT 115.4000 117.9000 115.8000 120.2000 ;
	    RECT 117.0000 117.9000 117.4000 120.2000 ;
	    RECT 119.8000 115.9000 120.2000 120.2000 ;
	    RECT 121.7000 117.9000 122.1000 120.2000 ;
	    RECT 123.8000 115.9000 124.2000 120.2000 ;
	    RECT 126.2000 115.9000 126.6000 120.2000 ;
	    RECT 127.0000 117.9000 127.4000 120.2000 ;
	    RECT 128.6000 116.1000 129.0000 120.2000 ;
	    RECT 131.8000 115.9000 132.2000 120.2000 ;
	    RECT 132.6000 115.9000 133.0000 120.2000 ;
	    RECT 134.7000 117.9000 135.1000 120.2000 ;
	    RECT 135.8000 117.9000 136.2000 120.2000 ;
	    RECT 137.4000 117.9000 137.8000 120.2000 ;
	    RECT 138.2000 115.9000 138.6000 120.2000 ;
	    RECT 140.3000 117.9000 140.7000 120.2000 ;
	    RECT 141.4000 117.9000 141.8000 120.2000 ;
	    RECT 143.0000 116.1000 143.4000 120.2000 ;
	    RECT 144.6000 115.9000 145.0000 120.2000 ;
	    RECT 146.7000 117.9000 147.1000 120.2000 ;
	    RECT 148.1000 117.9000 148.5000 120.2000 ;
	    RECT 150.2000 115.9000 150.6000 120.2000 ;
	    RECT 151.0000 117.9000 151.4000 120.2000 ;
	    RECT 152.6000 117.9000 153.0000 120.2000 ;
	    RECT 154.2000 115.9000 154.6000 120.2000 ;
	    RECT 155.0000 117.9000 155.4000 120.2000 ;
	    RECT 156.6000 117.9000 157.0000 120.2000 ;
	    RECT 157.4000 115.9000 157.8000 120.2000 ;
	    RECT 159.0000 115.9000 159.4000 120.2000 ;
	    RECT 162.2000 115.9000 162.6000 120.2000 ;
	    RECT 163.8000 116.0000 164.2000 120.2000 ;
	    RECT 166.6000 117.9000 167.0000 120.2000 ;
	    RECT 168.2000 117.9000 168.6000 120.2000 ;
	    RECT 171.0000 115.9000 171.4000 120.2000 ;
	    RECT 0.6000 100.8000 1.0000 103.1000 ;
	    RECT 2.2000 100.8000 2.6000 103.1000 ;
	    RECT 3.8000 100.8000 4.2000 102.9000 ;
	    RECT 5.4000 100.8000 5.8000 103.1000 ;
	    RECT 7.0000 100.8000 7.4000 103.1000 ;
	    RECT 8.6000 100.8000 9.0000 102.9000 ;
	    RECT 10.2000 100.8000 10.6000 103.1000 ;
	    RECT 12.1000 100.8000 12.5000 105.1000 ;
	    RECT 15.0000 100.8000 15.4000 102.9000 ;
	    RECT 16.6000 100.8000 17.0000 103.1000 ;
	    RECT 18.2000 100.8000 18.6000 104.5000 ;
	    RECT 21.1000 100.8000 21.5000 105.1000 ;
	    RECT 23.8000 100.8000 24.2000 102.9000 ;
	    RECT 25.4000 100.8000 25.8000 103.1000 ;
	    RECT 27.0000 100.8000 27.4000 105.1000 ;
	    RECT 27.8000 100.8000 28.2000 103.1000 ;
	    RECT 29.4000 100.8000 29.8000 102.9000 ;
	    RECT 31.0000 100.8000 31.4000 103.1000 ;
	    RECT 32.6000 100.8000 33.0000 103.1000 ;
	    RECT 34.2000 100.8000 34.6000 103.1000 ;
	    RECT 35.8000 100.8000 36.2000 102.9000 ;
	    RECT 37.4000 100.8000 37.8000 103.1000 ;
	    RECT 39.0000 100.8000 39.4000 102.9000 ;
	    RECT 40.6000 100.8000 41.0000 103.1000 ;
	    RECT 42.7000 100.8000 43.1000 105.1000 ;
	    RECT 45.4000 100.8000 45.8000 103.1000 ;
	    RECT 46.2000 100.8000 46.6000 103.1000 ;
	    RECT 47.8000 100.8000 48.2000 103.1000 ;
	    RECT 49.4000 100.8000 49.8000 102.9000 ;
	    RECT 51.0000 100.8000 51.4000 103.1000 ;
	    RECT 53.1000 100.8000 53.5000 105.1000 ;
	    RECT 55.0000 100.8000 55.4000 103.1000 ;
	    RECT 56.6000 100.8000 57.0000 102.9000 ;
	    RECT 58.2000 100.8000 58.6000 103.1000 ;
	    RECT 59.8000 100.8000 60.2000 103.1000 ;
	    RECT 63.0000 100.8000 63.4000 102.9000 ;
	    RECT 64.6000 100.8000 65.0000 103.1000 ;
	    RECT 66.2000 100.8000 66.6000 102.9000 ;
	    RECT 67.8000 100.8000 68.2000 103.1000 ;
	    RECT 69.4000 100.8000 69.8000 102.9000 ;
	    RECT 71.0000 100.8000 71.4000 103.1000 ;
	    RECT 71.8000 100.8000 72.2000 105.1000 ;
	    RECT 73.4000 100.8000 73.8000 105.1000 ;
	    RECT 74.2000 100.8000 74.6000 105.1000 ;
	    RECT 76.6000 100.8000 77.0000 105.1000 ;
	    RECT 78.2000 100.8000 78.6000 102.9000 ;
	    RECT 79.8000 100.8000 80.2000 103.1000 ;
	    RECT 81.4000 100.8000 81.8000 102.9000 ;
	    RECT 83.0000 100.8000 83.4000 103.1000 ;
	    RECT 83.8000 100.8000 84.2000 103.1000 ;
	    RECT 85.4000 100.8000 85.8000 102.9000 ;
	    RECT 87.0000 100.8000 87.4000 103.1000 ;
	    RECT 88.6000 100.8000 89.0000 102.9000 ;
	    RECT 91.0000 100.8000 91.4000 102.9000 ;
	    RECT 92.6000 100.8000 93.0000 103.1000 ;
	    RECT 94.2000 100.8000 94.6000 105.0000 ;
	    RECT 97.0000 100.8000 97.4000 103.1000 ;
	    RECT 98.6000 100.8000 99.0000 103.1000 ;
	    RECT 101.4000 100.8000 101.8000 105.1000 ;
	    RECT 103.8000 100.8000 104.2000 104.9000 ;
	    RECT 105.4000 100.8000 105.8000 103.1000 ;
	    RECT 106.2000 100.8000 106.6000 103.1000 ;
	    RECT 107.8000 100.8000 108.2000 104.9000 ;
	    RECT 111.8000 100.8000 112.2000 105.1000 ;
	    RECT 114.6000 100.8000 115.0000 103.1000 ;
	    RECT 116.2000 100.8000 116.6000 103.1000 ;
	    RECT 119.0000 100.8000 119.4000 105.0000 ;
	    RECT 121.4000 100.8000 121.8000 104.9000 ;
	    RECT 123.0000 100.8000 123.4000 103.1000 ;
	    RECT 123.8000 100.8000 124.2000 103.1000 ;
	    RECT 125.4000 100.8000 125.8000 104.9000 ;
	    RECT 127.0000 100.8000 127.4000 105.1000 ;
	    RECT 130.2000 100.8000 130.6000 105.1000 ;
	    RECT 131.0000 100.8000 131.4000 103.1000 ;
	    RECT 135.0000 100.8000 135.4000 104.5000 ;
	    RECT 136.6000 100.8000 137.0000 103.1000 ;
	    RECT 138.2000 100.8000 138.6000 103.1000 ;
	    RECT 139.0000 100.8000 139.4000 103.1000 ;
	    RECT 140.6000 100.8000 141.0000 103.1000 ;
	    RECT 142.2000 100.8000 142.6000 103.1000 ;
	    RECT 143.8000 100.8000 144.2000 105.0000 ;
	    RECT 146.6000 100.8000 147.0000 103.1000 ;
	    RECT 148.2000 100.8000 148.6000 103.1000 ;
	    RECT 151.0000 100.8000 151.4000 105.1000 ;
	    RECT 153.4000 100.8000 153.8000 105.1000 ;
	    RECT 156.2000 100.8000 156.6000 103.1000 ;
	    RECT 157.8000 100.8000 158.2000 103.1000 ;
	    RECT 160.6000 100.8000 161.0000 105.0000 ;
	    RECT 163.0000 100.8000 163.4000 105.0000 ;
	    RECT 165.8000 100.8000 166.2000 103.1000 ;
	    RECT 167.4000 100.8000 167.8000 103.1000 ;
	    RECT 170.2000 100.8000 170.6000 105.1000 ;
	    RECT 0.2000 100.2000 173.4000 100.8000 ;
	    RECT 1.4000 96.5000 1.8000 100.2000 ;
	    RECT 3.0000 97.9000 3.4000 100.2000 ;
	    RECT 4.6000 97.9000 5.0000 100.2000 ;
	    RECT 6.2000 97.9000 6.6000 100.2000 ;
	    RECT 8.3000 95.9000 8.7000 100.2000 ;
	    RECT 11.0000 98.1000 11.4000 100.2000 ;
	    RECT 12.6000 97.9000 13.0000 100.2000 ;
	    RECT 14.7000 95.9000 15.1000 100.2000 ;
	    RECT 16.6000 97.9000 17.0000 100.2000 ;
	    RECT 18.2000 97.9000 18.6000 100.2000 ;
	    RECT 19.0000 97.9000 19.4000 100.2000 ;
	    RECT 21.4000 98.1000 21.8000 100.2000 ;
	    RECT 23.0000 97.9000 23.4000 100.2000 ;
	    RECT 24.6000 96.5000 25.0000 100.2000 ;
	    RECT 26.2000 97.9000 26.6000 100.2000 ;
	    RECT 27.8000 98.1000 28.2000 100.2000 ;
	    RECT 29.4000 97.9000 29.8000 100.2000 ;
	    RECT 31.0000 98.1000 31.4000 100.2000 ;
	    RECT 33.7000 95.9000 34.1000 100.2000 ;
	    RECT 36.6000 98.1000 37.0000 100.2000 ;
	    RECT 38.2000 97.9000 38.6000 100.2000 ;
	    RECT 39.0000 97.9000 39.4000 100.2000 ;
	    RECT 40.6000 97.9000 41.0000 100.2000 ;
	    RECT 42.2000 97.9000 42.6000 100.2000 ;
	    RECT 44.3000 95.9000 44.7000 100.2000 ;
	    RECT 47.0000 98.1000 47.4000 100.2000 ;
	    RECT 48.6000 97.9000 49.0000 100.2000 ;
	    RECT 49.4000 97.9000 49.8000 100.2000 ;
	    RECT 51.0000 97.9000 51.4000 100.2000 ;
	    RECT 52.6000 97.9000 53.0000 100.2000 ;
	    RECT 54.7000 95.9000 55.1000 100.2000 ;
	    RECT 56.6000 97.9000 57.0000 100.2000 ;
	    RECT 58.2000 98.1000 58.6000 100.2000 ;
	    RECT 62.2000 97.9000 62.6000 100.2000 ;
	    RECT 63.0000 97.9000 63.4000 100.2000 ;
	    RECT 64.6000 97.9000 65.0000 100.2000 ;
	    RECT 66.2000 97.9000 66.6000 100.2000 ;
	    RECT 68.3000 95.9000 68.7000 100.2000 ;
	    RECT 71.0000 98.1000 71.4000 100.2000 ;
	    RECT 72.6000 97.9000 73.0000 100.2000 ;
	    RECT 74.2000 98.1000 74.6000 100.2000 ;
	    RECT 75.8000 97.9000 76.2000 100.2000 ;
	    RECT 77.9000 95.9000 78.3000 100.2000 ;
	    RECT 79.8000 97.9000 80.2000 100.2000 ;
	    RECT 81.4000 97.9000 81.8000 100.2000 ;
	    RECT 83.0000 98.1000 83.4000 100.2000 ;
	    RECT 84.6000 97.9000 85.0000 100.2000 ;
	    RECT 86.2000 97.9000 86.6000 100.2000 ;
	    RECT 87.0000 97.9000 87.4000 100.2000 ;
	    RECT 88.6000 98.1000 89.0000 100.2000 ;
	    RECT 90.2000 97.9000 90.6000 100.2000 ;
	    RECT 91.8000 98.1000 92.2000 100.2000 ;
	    RECT 94.7000 95.9000 95.1000 100.2000 ;
	    RECT 97.4000 98.1000 97.8000 100.2000 ;
	    RECT 99.0000 97.9000 99.4000 100.2000 ;
	    RECT 100.6000 96.5000 101.0000 100.2000 ;
	    RECT 104.6000 96.5000 105.0000 100.2000 ;
	    RECT 107.0000 96.5000 107.4000 100.2000 ;
	    RECT 110.2000 96.5000 110.6000 100.2000 ;
	    RECT 115.0000 96.5000 115.4000 100.2000 ;
	    RECT 118.2000 96.0000 118.6000 100.2000 ;
	    RECT 121.0000 97.9000 121.4000 100.2000 ;
	    RECT 122.6000 97.9000 123.0000 100.2000 ;
	    RECT 125.4000 95.9000 125.8000 100.2000 ;
	    RECT 127.8000 95.9000 128.2000 100.2000 ;
	    RECT 130.6000 97.9000 131.0000 100.2000 ;
	    RECT 132.2000 97.9000 132.6000 100.2000 ;
	    RECT 135.0000 96.0000 135.4000 100.2000 ;
	    RECT 136.6000 97.9000 137.0000 100.2000 ;
	    RECT 138.2000 97.9000 138.6000 100.2000 ;
	    RECT 139.8000 97.9000 140.2000 100.2000 ;
	    RECT 141.4000 96.5000 141.8000 100.2000 ;
	    RECT 143.8000 95.9000 144.2000 100.2000 ;
	    RECT 146.6000 97.9000 147.0000 100.2000 ;
	    RECT 148.2000 97.9000 148.6000 100.2000 ;
	    RECT 151.0000 96.0000 151.4000 100.2000 ;
	    RECT 152.6000 95.9000 153.0000 100.2000 ;
	    RECT 154.2000 95.9000 154.6000 100.2000 ;
	    RECT 155.8000 95.9000 156.2000 100.2000 ;
	    RECT 157.4000 95.9000 157.8000 100.2000 ;
	    RECT 159.0000 95.9000 159.4000 100.2000 ;
	    RECT 160.6000 96.0000 161.0000 100.2000 ;
	    RECT 163.4000 97.9000 163.8000 100.2000 ;
	    RECT 165.0000 97.9000 165.4000 100.2000 ;
	    RECT 167.8000 95.9000 168.2000 100.2000 ;
	    RECT 170.2000 96.1000 170.6000 100.2000 ;
	    RECT 171.8000 97.9000 172.2000 100.2000 ;
	    RECT 0.6000 80.8000 1.0000 83.1000 ;
	    RECT 2.2000 80.8000 2.6000 83.1000 ;
	    RECT 3.8000 80.8000 4.2000 83.1000 ;
	    RECT 5.4000 80.8000 5.8000 83.1000 ;
	    RECT 7.5000 80.8000 7.9000 85.1000 ;
	    RECT 10.2000 80.8000 10.6000 82.9000 ;
	    RECT 11.8000 80.8000 12.2000 83.1000 ;
	    RECT 13.4000 80.8000 13.8000 82.9000 ;
	    RECT 15.0000 80.8000 15.4000 83.1000 ;
	    RECT 15.8000 80.8000 16.2000 83.1000 ;
	    RECT 17.4000 80.8000 17.8000 83.1000 ;
	    RECT 19.0000 80.8000 19.4000 83.1000 ;
	    RECT 21.1000 80.8000 21.5000 85.1000 ;
	    RECT 23.0000 80.8000 23.4000 83.1000 ;
	    RECT 24.6000 80.8000 25.0000 82.9000 ;
	    RECT 26.2000 80.8000 26.6000 83.1000 ;
	    RECT 27.8000 80.8000 28.2000 82.9000 ;
	    RECT 30.2000 80.8000 30.6000 82.9000 ;
	    RECT 31.8000 80.8000 32.2000 83.1000 ;
	    RECT 32.6000 80.8000 33.0000 83.1000 ;
	    RECT 34.2000 80.8000 34.6000 83.1000 ;
	    RECT 36.1000 80.8000 36.5000 85.1000 ;
	    RECT 38.2000 80.8000 38.6000 83.1000 ;
	    RECT 39.8000 80.8000 40.2000 83.1000 ;
	    RECT 40.6000 80.8000 41.0000 83.1000 ;
	    RECT 42.2000 80.8000 42.6000 82.9000 ;
	    RECT 43.8000 80.8000 44.2000 83.1000 ;
	    RECT 45.4000 80.8000 45.8000 82.9000 ;
	    RECT 47.0000 80.8000 47.4000 83.1000 ;
	    RECT 48.6000 80.8000 49.0000 83.1000 ;
	    RECT 50.2000 80.8000 50.6000 83.1000 ;
	    RECT 52.3000 80.8000 52.7000 85.1000 ;
	    RECT 55.0000 80.8000 55.4000 82.9000 ;
	    RECT 56.6000 80.8000 57.0000 83.1000 ;
	    RECT 58.7000 80.8000 59.1000 85.1000 ;
	    RECT 62.2000 80.8000 62.6000 83.1000 ;
	    RECT 64.6000 80.8000 65.0000 84.5000 ;
	    RECT 66.2000 80.8000 66.6000 83.1000 ;
	    RECT 67.8000 80.8000 68.2000 83.1000 ;
	    RECT 68.6000 80.8000 69.0000 83.1000 ;
	    RECT 70.2000 80.8000 70.6000 83.1000 ;
	    RECT 71.8000 80.8000 72.2000 82.9000 ;
	    RECT 73.4000 80.8000 73.8000 83.1000 ;
	    RECT 75.0000 80.8000 75.4000 82.9000 ;
	    RECT 76.6000 80.8000 77.0000 83.1000 ;
	    RECT 78.2000 80.8000 78.6000 82.9000 ;
	    RECT 79.8000 80.8000 80.2000 83.1000 ;
	    RECT 80.6000 80.8000 81.0000 83.1000 ;
	    RECT 82.2000 80.8000 82.6000 82.9000 ;
	    RECT 85.1000 80.8000 85.5000 85.1000 ;
	    RECT 87.0000 80.8000 87.4000 83.1000 ;
	    RECT 88.6000 80.8000 89.0000 83.1000 ;
	    RECT 89.4000 80.8000 89.8000 83.1000 ;
	    RECT 91.0000 80.8000 91.4000 83.1000 ;
	    RECT 92.6000 80.8000 93.0000 82.9000 ;
	    RECT 94.2000 80.8000 94.6000 83.1000 ;
	    RECT 95.8000 80.8000 96.2000 82.9000 ;
	    RECT 97.4000 80.8000 97.8000 83.1000 ;
	    RECT 99.0000 80.8000 99.4000 82.9000 ;
	    RECT 100.6000 80.8000 101.0000 83.1000 ;
	    RECT 102.2000 80.8000 102.6000 85.0000 ;
	    RECT 105.0000 80.8000 105.4000 83.1000 ;
	    RECT 106.6000 80.8000 107.0000 83.1000 ;
	    RECT 109.4000 80.8000 109.8000 85.1000 ;
	    RECT 113.4000 80.8000 113.8000 85.1000 ;
	    RECT 115.0000 80.8000 115.4000 84.5000 ;
	    RECT 117.4000 80.8000 117.8000 84.9000 ;
	    RECT 119.0000 80.8000 119.4000 83.1000 ;
	    RECT 120.6000 80.8000 121.0000 85.1000 ;
	    RECT 123.4000 80.8000 123.8000 83.1000 ;
	    RECT 125.0000 80.8000 125.4000 83.1000 ;
	    RECT 127.8000 80.8000 128.2000 85.0000 ;
	    RECT 129.4000 80.8000 129.8000 83.1000 ;
	    RECT 131.0000 80.8000 131.4000 84.9000 ;
	    RECT 133.4000 80.8000 133.8000 85.0000 ;
	    RECT 136.2000 80.8000 136.6000 83.1000 ;
	    RECT 137.8000 80.8000 138.2000 83.1000 ;
	    RECT 140.6000 80.8000 141.0000 85.1000 ;
	    RECT 143.8000 80.8000 144.2000 84.5000 ;
	    RECT 145.4000 80.8000 145.8000 85.1000 ;
	    RECT 147.0000 80.8000 147.4000 85.1000 ;
	    RECT 148.6000 80.8000 149.0000 85.1000 ;
	    RECT 150.2000 80.8000 150.6000 85.1000 ;
	    RECT 151.8000 80.8000 152.2000 85.1000 ;
	    RECT 153.4000 80.8000 153.8000 85.1000 ;
	    RECT 156.2000 80.8000 156.6000 83.1000 ;
	    RECT 157.8000 80.8000 158.2000 83.1000 ;
	    RECT 160.6000 80.8000 161.0000 85.0000 ;
	    RECT 162.2000 80.8000 162.6000 83.1000 ;
	    RECT 163.8000 80.8000 164.2000 84.9000 ;
	    RECT 166.2000 80.8000 166.6000 84.9000 ;
	    RECT 167.8000 80.8000 168.2000 83.1000 ;
	    RECT 169.4000 80.8000 169.8000 84.5000 ;
	    RECT 171.0000 80.8000 171.4000 83.1000 ;
	    RECT 172.6000 80.8000 173.0000 83.1000 ;
	    RECT 0.2000 80.2000 173.4000 80.8000 ;
	    RECT 0.6000 77.9000 1.0000 80.2000 ;
	    RECT 2.2000 77.9000 2.6000 80.2000 ;
	    RECT 4.1000 75.9000 4.5000 80.2000 ;
	    RECT 7.0000 76.5000 7.4000 80.2000 ;
	    RECT 9.4000 76.5000 9.8000 80.2000 ;
	    RECT 11.8000 77.9000 12.2000 80.2000 ;
	    RECT 12.6000 77.9000 13.0000 80.2000 ;
	    RECT 14.2000 77.9000 14.6000 80.2000 ;
	    RECT 16.3000 75.9000 16.7000 80.2000 ;
	    RECT 18.2000 77.9000 18.6000 80.2000 ;
	    RECT 19.8000 77.9000 20.2000 80.2000 ;
	    RECT 21.4000 77.9000 21.8000 80.2000 ;
	    RECT 22.2000 77.9000 22.6000 80.2000 ;
	    RECT 23.8000 77.9000 24.2000 80.2000 ;
	    RECT 25.4000 77.9000 25.8000 80.2000 ;
	    RECT 26.2000 77.9000 26.6000 80.2000 ;
	    RECT 27.8000 77.9000 28.2000 80.2000 ;
	    RECT 29.4000 77.9000 29.8000 80.2000 ;
	    RECT 31.3000 75.9000 31.7000 80.2000 ;
	    RECT 34.2000 77.9000 34.6000 80.2000 ;
	    RECT 35.8000 77.9000 36.2000 80.2000 ;
	    RECT 36.6000 75.9000 37.0000 80.2000 ;
	    RECT 38.7000 77.9000 39.1000 80.2000 ;
	    RECT 40.6000 75.9000 41.0000 80.2000 ;
	    RECT 41.4000 77.9000 41.8000 80.2000 ;
	    RECT 43.0000 77.9000 43.4000 80.2000 ;
	    RECT 44.6000 77.9000 45.0000 80.2000 ;
	    RECT 46.7000 75.9000 47.1000 80.2000 ;
	    RECT 49.4000 78.1000 49.8000 80.2000 ;
	    RECT 51.0000 77.9000 51.4000 80.2000 ;
	    RECT 53.1000 75.9000 53.5000 80.2000 ;
	    RECT 55.8000 76.5000 56.2000 80.2000 ;
	    RECT 58.2000 78.1000 58.6000 80.2000 ;
	    RECT 59.8000 77.9000 60.2000 80.2000 ;
	    RECT 63.0000 78.1000 63.4000 80.2000 ;
	    RECT 64.6000 77.9000 65.0000 80.2000 ;
	    RECT 66.2000 76.5000 66.6000 80.2000 ;
	    RECT 68.6000 78.1000 69.0000 80.2000 ;
	    RECT 70.2000 77.9000 70.6000 80.2000 ;
	    RECT 71.8000 78.1000 72.2000 80.2000 ;
	    RECT 73.4000 77.9000 73.8000 80.2000 ;
	    RECT 75.3000 75.9000 75.7000 80.2000 ;
	    RECT 78.7000 75.9000 79.1000 80.2000 ;
	    RECT 80.6000 77.9000 81.0000 80.2000 ;
	    RECT 82.2000 78.1000 82.6000 80.2000 ;
	    RECT 83.8000 77.9000 84.2000 80.2000 ;
	    RECT 85.4000 77.9000 85.8000 80.2000 ;
	    RECT 87.8000 76.1000 88.2000 80.2000 ;
	    RECT 89.4000 77.9000 89.8000 80.2000 ;
	    RECT 90.2000 77.9000 90.6000 80.2000 ;
	    RECT 91.8000 76.1000 92.2000 80.2000 ;
	    RECT 94.2000 78.1000 94.6000 80.2000 ;
	    RECT 95.8000 77.9000 96.2000 80.2000 ;
	    RECT 97.4000 76.5000 97.8000 80.2000 ;
	    RECT 100.6000 76.5000 101.0000 80.2000 ;
	    RECT 103.0000 75.9000 103.4000 80.2000 ;
	    RECT 104.6000 75.9000 105.0000 80.2000 ;
	    RECT 106.2000 75.9000 106.6000 80.2000 ;
	    RECT 107.8000 75.9000 108.2000 80.2000 ;
	    RECT 109.4000 75.9000 109.8000 80.2000 ;
	    RECT 111.0000 76.5000 111.4000 80.2000 ;
	    RECT 115.0000 76.0000 115.4000 80.2000 ;
	    RECT 117.8000 77.9000 118.2000 80.2000 ;
	    RECT 119.4000 77.9000 119.8000 80.2000 ;
	    RECT 122.2000 75.9000 122.6000 80.2000 ;
	    RECT 123.8000 77.9000 124.2000 80.2000 ;
	    RECT 125.4000 76.1000 125.8000 80.2000 ;
	    RECT 127.8000 76.0000 128.2000 80.2000 ;
	    RECT 130.6000 77.9000 131.0000 80.2000 ;
	    RECT 132.2000 77.9000 132.6000 80.2000 ;
	    RECT 135.0000 75.9000 135.4000 80.2000 ;
	    RECT 137.4000 76.5000 137.8000 80.2000 ;
	    RECT 140.6000 76.5000 141.0000 80.2000 ;
	    RECT 142.2000 75.9000 142.6000 80.2000 ;
	    RECT 144.6000 76.5000 145.0000 80.2000 ;
	    RECT 147.8000 76.5000 148.2000 80.2000 ;
	    RECT 151.8000 76.5000 152.2000 80.2000 ;
	    RECT 154.2000 76.0000 154.6000 80.2000 ;
	    RECT 157.0000 77.9000 157.4000 80.2000 ;
	    RECT 158.6000 77.9000 159.0000 80.2000 ;
	    RECT 161.4000 75.9000 161.8000 80.2000 ;
	    RECT 163.8000 76.0000 164.2000 80.2000 ;
	    RECT 166.6000 77.9000 167.0000 80.2000 ;
	    RECT 168.2000 77.9000 168.6000 80.2000 ;
	    RECT 171.0000 75.9000 171.4000 80.2000 ;
	    RECT 1.4000 60.8000 1.8000 62.9000 ;
	    RECT 3.0000 60.8000 3.4000 63.1000 ;
	    RECT 3.8000 60.8000 4.2000 65.1000 ;
	    RECT 6.7000 60.8000 7.1000 65.1000 ;
	    RECT 8.6000 60.8000 9.0000 63.1000 ;
	    RECT 10.2000 60.8000 10.6000 62.9000 ;
	    RECT 11.8000 60.8000 12.2000 63.1000 ;
	    RECT 13.4000 60.8000 13.8000 62.9000 ;
	    RECT 15.8000 60.8000 16.2000 62.9000 ;
	    RECT 17.4000 60.8000 17.8000 63.1000 ;
	    RECT 18.2000 60.8000 18.6000 63.1000 ;
	    RECT 19.8000 60.8000 20.2000 62.9000 ;
	    RECT 21.4000 60.8000 21.8000 63.1000 ;
	    RECT 23.0000 60.8000 23.4000 63.1000 ;
	    RECT 24.6000 60.8000 25.0000 62.9000 ;
	    RECT 26.2000 60.8000 26.6000 63.1000 ;
	    RECT 28.3000 60.8000 28.7000 65.1000 ;
	    RECT 30.2000 60.8000 30.6000 63.1000 ;
	    RECT 31.8000 60.8000 32.2000 62.9000 ;
	    RECT 33.4000 60.8000 33.8000 63.1000 ;
	    RECT 35.0000 60.8000 35.4000 63.1000 ;
	    RECT 36.6000 60.8000 37.0000 63.1000 ;
	    RECT 37.4000 60.8000 37.8000 63.1000 ;
	    RECT 39.0000 60.8000 39.4000 63.1000 ;
	    RECT 39.8000 60.8000 40.2000 63.1000 ;
	    RECT 41.4000 60.8000 41.8000 63.1000 ;
	    RECT 42.2000 60.8000 42.6000 63.1000 ;
	    RECT 43.8000 60.8000 44.2000 65.1000 ;
	    RECT 45.9000 60.8000 46.3000 63.1000 ;
	    RECT 47.0000 60.8000 47.4000 63.1000 ;
	    RECT 48.6000 60.8000 49.0000 63.1000 ;
	    RECT 49.4000 60.8000 49.8000 63.1000 ;
	    RECT 51.3000 60.8000 51.7000 63.1000 ;
	    RECT 53.4000 60.8000 53.8000 65.1000 ;
	    RECT 54.2000 60.8000 54.6000 63.1000 ;
	    RECT 55.8000 60.8000 56.2000 63.1000 ;
	    RECT 57.4000 60.8000 57.8000 63.1000 ;
	    RECT 58.2000 60.8000 58.6000 63.1000 ;
	    RECT 59.8000 60.8000 60.2000 63.1000 ;
	    RECT 62.2000 60.8000 62.6000 63.1000 ;
	    RECT 63.8000 60.8000 64.2000 63.1000 ;
	    RECT 65.4000 60.8000 65.8000 63.1000 ;
	    RECT 66.2000 60.8000 66.6000 63.1000 ;
	    RECT 67.8000 60.8000 68.2000 63.1000 ;
	    RECT 69.4000 60.8000 69.8000 63.1000 ;
	    RECT 71.3000 60.8000 71.7000 65.1000 ;
	    RECT 73.4000 60.8000 73.8000 63.1000 ;
	    RECT 75.0000 60.8000 75.4000 63.1000 ;
	    RECT 76.6000 60.8000 77.0000 63.1000 ;
	    RECT 77.4000 60.8000 77.8000 63.1000 ;
	    RECT 79.0000 60.8000 79.4000 64.9000 ;
	    RECT 80.6000 60.8000 81.0000 63.1000 ;
	    RECT 82.2000 60.8000 82.6000 64.9000 ;
	    RECT 84.6000 60.8000 85.0000 65.0000 ;
	    RECT 87.4000 60.8000 87.8000 63.1000 ;
	    RECT 89.0000 60.8000 89.4000 63.1000 ;
	    RECT 91.8000 60.8000 92.2000 65.1000 ;
	    RECT 94.2000 60.8000 94.6000 64.5000 ;
	    RECT 96.6000 60.8000 97.0000 65.1000 ;
	    RECT 98.2000 60.8000 98.6000 63.1000 ;
	    RECT 99.8000 60.8000 100.2000 64.9000 ;
	    RECT 102.2000 60.8000 102.6000 65.0000 ;
	    RECT 105.0000 60.8000 105.4000 63.1000 ;
	    RECT 106.6000 60.8000 107.0000 63.1000 ;
	    RECT 109.4000 60.8000 109.8000 65.1000 ;
	    RECT 112.6000 60.8000 113.0000 65.1000 ;
	    RECT 114.2000 60.8000 114.6000 65.1000 ;
	    RECT 115.8000 60.8000 116.2000 65.1000 ;
	    RECT 117.4000 60.8000 117.8000 65.1000 ;
	    RECT 119.0000 60.8000 119.4000 65.1000 ;
	    RECT 120.6000 60.8000 121.0000 65.0000 ;
	    RECT 123.4000 60.8000 123.8000 63.1000 ;
	    RECT 125.0000 60.8000 125.4000 63.1000 ;
	    RECT 127.8000 60.8000 128.2000 65.1000 ;
	    RECT 130.2000 60.8000 130.6000 64.9000 ;
	    RECT 131.8000 60.8000 132.2000 63.1000 ;
	    RECT 133.4000 60.8000 133.8000 65.0000 ;
	    RECT 136.2000 60.8000 136.6000 63.1000 ;
	    RECT 137.8000 60.8000 138.2000 63.1000 ;
	    RECT 140.6000 60.8000 141.0000 65.1000 ;
	    RECT 142.2000 60.8000 142.6000 63.1000 ;
	    RECT 143.8000 60.8000 144.2000 64.9000 ;
	    RECT 146.2000 60.8000 146.6000 65.1000 ;
	    RECT 149.0000 60.8000 149.4000 63.1000 ;
	    RECT 150.6000 60.8000 151.0000 63.1000 ;
	    RECT 153.4000 60.8000 153.8000 65.0000 ;
	    RECT 155.0000 60.8000 155.4000 63.1000 ;
	    RECT 156.6000 60.8000 157.0000 64.9000 ;
	    RECT 159.0000 60.8000 159.4000 65.0000 ;
	    RECT 161.8000 60.8000 162.2000 63.1000 ;
	    RECT 163.4000 60.8000 163.8000 63.1000 ;
	    RECT 166.2000 60.8000 166.6000 65.1000 ;
	    RECT 168.6000 60.8000 169.0000 64.5000 ;
	    RECT 171.0000 60.8000 171.4000 64.5000 ;
	    RECT 0.2000 60.2000 173.4000 60.8000 ;
	    RECT 1.4000 58.1000 1.8000 60.2000 ;
	    RECT 3.0000 57.9000 3.4000 60.2000 ;
	    RECT 4.6000 58.1000 5.0000 60.2000 ;
	    RECT 6.2000 57.9000 6.6000 60.2000 ;
	    RECT 7.0000 55.9000 7.4000 60.2000 ;
	    RECT 9.4000 57.9000 9.8000 60.2000 ;
	    RECT 10.2000 55.9000 10.6000 60.2000 ;
	    RECT 12.3000 57.9000 12.7000 60.2000 ;
	    RECT 14.2000 58.1000 14.6000 60.2000 ;
	    RECT 15.8000 57.9000 16.2000 60.2000 ;
	    RECT 17.4000 58.1000 17.8000 60.2000 ;
	    RECT 19.0000 57.9000 19.4000 60.2000 ;
	    RECT 19.8000 57.9000 20.2000 60.2000 ;
	    RECT 21.4000 58.1000 21.8000 60.2000 ;
	    RECT 23.0000 57.9000 23.4000 60.2000 ;
	    RECT 24.6000 58.1000 25.0000 60.2000 ;
	    RECT 26.2000 57.9000 26.6000 60.2000 ;
	    RECT 27.8000 58.1000 28.2000 60.2000 ;
	    RECT 30.5000 55.9000 30.9000 60.2000 ;
	    RECT 33.4000 56.5000 33.8000 60.2000 ;
	    RECT 36.6000 56.5000 37.0000 60.2000 ;
	    RECT 39.8000 56.5000 40.2000 60.2000 ;
	    RECT 43.0000 56.5000 43.4000 60.2000 ;
	    RECT 46.2000 55.9000 46.6000 60.2000 ;
	    RECT 47.8000 56.0000 48.2000 60.2000 ;
	    RECT 50.6000 57.9000 51.0000 60.2000 ;
	    RECT 52.2000 57.9000 52.6000 60.2000 ;
	    RECT 55.0000 55.9000 55.4000 60.2000 ;
	    RECT 57.4000 58.1000 57.8000 60.2000 ;
	    RECT 59.0000 57.9000 59.4000 60.2000 ;
	    RECT 62.2000 56.0000 62.6000 60.2000 ;
	    RECT 65.0000 57.9000 65.4000 60.2000 ;
	    RECT 66.6000 57.9000 67.0000 60.2000 ;
	    RECT 69.4000 55.9000 69.8000 60.2000 ;
	    RECT 71.8000 58.1000 72.2000 60.2000 ;
	    RECT 73.4000 57.9000 73.8000 60.2000 ;
	    RECT 75.0000 58.1000 75.4000 60.2000 ;
	    RECT 76.6000 57.9000 77.0000 60.2000 ;
	    RECT 77.4000 57.9000 77.8000 60.2000 ;
	    RECT 79.0000 58.1000 79.4000 60.2000 ;
	    RECT 81.4000 56.0000 81.8000 60.2000 ;
	    RECT 84.2000 57.9000 84.6000 60.2000 ;
	    RECT 85.8000 57.9000 86.2000 60.2000 ;
	    RECT 88.6000 55.9000 89.0000 60.2000 ;
	    RECT 91.0000 56.0000 91.4000 60.2000 ;
	    RECT 93.8000 57.9000 94.2000 60.2000 ;
	    RECT 95.4000 57.9000 95.8000 60.2000 ;
	    RECT 98.2000 55.9000 98.6000 60.2000 ;
	    RECT 100.6000 55.9000 101.0000 60.2000 ;
	    RECT 101.4000 55.9000 101.8000 60.2000 ;
	    RECT 103.0000 55.9000 103.4000 60.2000 ;
	    RECT 104.6000 55.9000 105.0000 60.2000 ;
	    RECT 106.2000 55.9000 106.6000 60.2000 ;
	    RECT 107.8000 55.9000 108.2000 60.2000 ;
	    RECT 109.4000 58.1000 109.8000 60.2000 ;
	    RECT 111.0000 57.9000 111.4000 60.2000 ;
	    RECT 114.2000 56.5000 114.6000 60.2000 ;
	    RECT 115.8000 57.9000 116.2000 60.2000 ;
	    RECT 117.4000 58.1000 117.8000 60.2000 ;
	    RECT 119.0000 57.9000 119.4000 60.2000 ;
	    RECT 120.6000 57.9000 121.0000 60.2000 ;
	    RECT 122.2000 57.9000 122.6000 60.2000 ;
	    RECT 123.8000 56.5000 124.2000 60.2000 ;
	    RECT 125.4000 57.9000 125.8000 60.2000 ;
	    RECT 127.0000 57.9000 127.4000 60.2000 ;
	    RECT 128.6000 57.9000 129.0000 60.2000 ;
	    RECT 129.4000 57.9000 129.8000 60.2000 ;
	    RECT 131.0000 57.9000 131.4000 60.2000 ;
	    RECT 132.6000 57.9000 133.0000 60.2000 ;
	    RECT 134.2000 55.9000 134.6000 60.2000 ;
	    RECT 135.0000 57.9000 135.4000 60.2000 ;
	    RECT 136.6000 58.1000 137.0000 60.2000 ;
	    RECT 139.5000 55.9000 139.9000 60.2000 ;
	    RECT 141.4000 57.9000 141.8000 60.2000 ;
	    RECT 143.0000 58.1000 143.4000 60.2000 ;
	    RECT 144.6000 57.9000 145.0000 60.2000 ;
	    RECT 146.2000 58.1000 146.6000 60.2000 ;
	    RECT 147.8000 57.9000 148.2000 60.2000 ;
	    RECT 149.4000 57.9000 149.8000 60.2000 ;
	    RECT 151.0000 57.9000 151.4000 60.2000 ;
	    RECT 151.8000 57.9000 152.2000 60.2000 ;
	    RECT 153.4000 57.9000 153.8000 60.2000 ;
	    RECT 154.2000 57.9000 154.6000 60.2000 ;
	    RECT 155.8000 57.9000 156.2000 60.2000 ;
	    RECT 156.6000 57.9000 157.0000 60.2000 ;
	    RECT 158.2000 57.9000 158.6000 60.2000 ;
	    RECT 159.8000 55.9000 160.2000 60.2000 ;
	    RECT 161.9000 57.9000 162.3000 60.2000 ;
	    RECT 163.0000 57.9000 163.4000 60.2000 ;
	    RECT 164.6000 56.1000 165.0000 60.2000 ;
	    RECT 166.2000 57.9000 166.6000 60.2000 ;
	    RECT 167.8000 57.9000 168.2000 60.2000 ;
	    RECT 169.4000 57.9000 169.8000 60.2000 ;
	    RECT 171.0000 56.5000 171.4000 60.2000 ;
	    RECT 0.6000 40.8000 1.0000 43.1000 ;
	    RECT 2.2000 40.8000 2.6000 42.9000 ;
	    RECT 4.9000 40.8000 5.3000 45.1000 ;
	    RECT 7.8000 40.8000 8.2000 43.1000 ;
	    RECT 8.6000 40.8000 9.0000 43.1000 ;
	    RECT 10.2000 40.8000 10.6000 43.1000 ;
	    RECT 11.0000 40.8000 11.4000 43.1000 ;
	    RECT 12.6000 40.8000 13.0000 43.1000 ;
	    RECT 13.4000 40.8000 13.8000 43.1000 ;
	    RECT 15.0000 40.8000 15.4000 43.1000 ;
	    RECT 16.6000 40.8000 17.0000 43.1000 ;
	    RECT 17.4000 40.8000 17.8000 43.1000 ;
	    RECT 19.0000 40.8000 19.4000 42.9000 ;
	    RECT 21.7000 40.8000 22.1000 45.1000 ;
	    RECT 23.8000 40.8000 24.2000 43.1000 ;
	    RECT 25.4000 40.8000 25.8000 42.9000 ;
	    RECT 27.0000 40.8000 27.4000 43.1000 ;
	    RECT 28.6000 40.8000 29.0000 43.1000 ;
	    RECT 29.4000 40.8000 29.8000 43.1000 ;
	    RECT 31.0000 40.8000 31.4000 42.9000 ;
	    RECT 32.6000 40.8000 33.0000 43.1000 ;
	    RECT 34.2000 40.8000 34.6000 42.9000 ;
	    RECT 36.9000 40.8000 37.3000 45.1000 ;
	    RECT 39.0000 40.8000 39.4000 43.1000 ;
	    RECT 40.6000 40.8000 41.0000 43.1000 ;
	    RECT 41.4000 40.8000 41.8000 43.1000 ;
	    RECT 43.0000 40.8000 43.4000 43.1000 ;
	    RECT 43.8000 40.8000 44.2000 43.1000 ;
	    RECT 45.4000 40.8000 45.8000 43.1000 ;
	    RECT 47.0000 40.8000 47.4000 43.1000 ;
	    RECT 48.6000 40.8000 49.0000 43.1000 ;
	    RECT 49.4000 40.8000 49.8000 43.1000 ;
	    RECT 51.0000 40.8000 51.4000 43.1000 ;
	    RECT 52.6000 40.8000 53.0000 43.1000 ;
	    RECT 54.7000 40.8000 55.1000 45.1000 ;
	    RECT 57.4000 40.8000 57.8000 42.9000 ;
	    RECT 59.0000 40.8000 59.4000 43.1000 ;
	    RECT 62.7000 40.8000 63.1000 45.1000 ;
	    RECT 65.4000 40.8000 65.8000 42.9000 ;
	    RECT 67.0000 40.8000 67.4000 43.1000 ;
	    RECT 67.8000 40.8000 68.2000 43.1000 ;
	    RECT 69.4000 40.8000 69.8000 42.9000 ;
	    RECT 71.0000 40.8000 71.4000 43.1000 ;
	    RECT 72.6000 40.8000 73.0000 42.9000 ;
	    RECT 75.3000 40.8000 75.7000 45.1000 ;
	    RECT 77.4000 40.8000 77.8000 43.1000 ;
	    RECT 79.0000 40.8000 79.4000 43.1000 ;
	    RECT 79.8000 40.8000 80.2000 43.1000 ;
	    RECT 81.4000 40.8000 81.8000 43.1000 ;
	    RECT 83.0000 40.8000 83.4000 43.1000 ;
	    RECT 83.8000 40.8000 84.2000 43.1000 ;
	    RECT 85.4000 40.8000 85.8000 42.9000 ;
	    RECT 88.1000 40.8000 88.5000 45.1000 ;
	    RECT 90.2000 40.8000 90.6000 43.1000 ;
	    RECT 91.8000 40.8000 92.2000 43.1000 ;
	    RECT 93.4000 40.8000 93.8000 43.1000 ;
	    RECT 95.0000 40.8000 95.4000 43.1000 ;
	    RECT 96.6000 40.8000 97.0000 42.9000 ;
	    RECT 98.2000 40.8000 98.6000 43.1000 ;
	    RECT 99.0000 40.8000 99.4000 43.1000 ;
	    RECT 100.6000 40.8000 101.0000 42.9000 ;
	    RECT 102.2000 40.8000 102.6000 43.1000 ;
	    RECT 103.8000 40.8000 104.2000 43.1000 ;
	    RECT 104.6000 40.8000 105.0000 43.1000 ;
	    RECT 106.2000 40.8000 106.6000 43.1000 ;
	    RECT 107.3000 40.8000 107.7000 43.1000 ;
	    RECT 109.4000 40.8000 109.8000 45.1000 ;
	    RECT 111.0000 40.8000 111.4000 43.1000 ;
	    RECT 113.4000 40.8000 113.8000 45.1000 ;
	    RECT 115.0000 40.8000 115.4000 45.1000 ;
	    RECT 115.8000 40.8000 116.2000 43.1000 ;
	    RECT 117.4000 40.8000 117.8000 42.9000 ;
	    RECT 120.1000 40.8000 120.5000 45.1000 ;
	    RECT 122.2000 40.8000 122.6000 43.1000 ;
	    RECT 123.8000 40.8000 124.2000 42.9000 ;
	    RECT 125.4000 40.8000 125.8000 43.1000 ;
	    RECT 127.0000 40.8000 127.4000 42.9000 ;
	    RECT 128.6000 40.8000 129.0000 43.1000 ;
	    RECT 130.2000 40.8000 130.6000 42.9000 ;
	    RECT 132.9000 40.8000 133.3000 45.1000 ;
	    RECT 136.3000 40.8000 136.7000 45.1000 ;
	    RECT 139.5000 40.8000 139.9000 45.1000 ;
	    RECT 141.4000 40.8000 141.8000 43.1000 ;
	    RECT 143.0000 40.8000 143.4000 42.9000 ;
	    RECT 144.6000 40.8000 145.0000 43.1000 ;
	    RECT 146.2000 40.8000 146.6000 43.1000 ;
	    RECT 147.0000 40.8000 147.4000 43.1000 ;
	    RECT 148.6000 40.8000 149.0000 42.9000 ;
	    RECT 150.2000 40.8000 150.6000 43.1000 ;
	    RECT 151.8000 40.8000 152.2000 42.9000 ;
	    RECT 154.7000 40.8000 155.1000 45.1000 ;
	    RECT 157.4000 40.8000 157.8000 42.9000 ;
	    RECT 159.0000 40.8000 159.4000 43.1000 ;
	    RECT 159.8000 40.8000 160.2000 43.1000 ;
	    RECT 161.4000 40.8000 161.8000 43.1000 ;
	    RECT 162.2000 40.8000 162.6000 43.1000 ;
	    RECT 163.8000 40.8000 164.2000 42.9000 ;
	    RECT 166.2000 40.8000 166.6000 42.9000 ;
	    RECT 167.8000 40.8000 168.2000 43.1000 ;
	    RECT 169.7000 40.8000 170.1000 45.1000 ;
	    RECT 0.2000 40.2000 173.4000 40.8000 ;
	    RECT 1.4000 38.1000 1.8000 40.2000 ;
	    RECT 3.0000 37.9000 3.4000 40.2000 ;
	    RECT 4.6000 38.1000 5.0000 40.2000 ;
	    RECT 6.2000 37.9000 6.6000 40.2000 ;
	    RECT 7.0000 37.9000 7.4000 40.2000 ;
	    RECT 8.6000 38.1000 9.0000 40.2000 ;
	    RECT 11.0000 38.1000 11.4000 40.2000 ;
	    RECT 12.6000 37.9000 13.0000 40.2000 ;
	    RECT 14.2000 38.1000 14.6000 40.2000 ;
	    RECT 15.8000 37.9000 16.2000 40.2000 ;
	    RECT 16.6000 37.9000 17.0000 40.2000 ;
	    RECT 18.2000 38.1000 18.6000 40.2000 ;
	    RECT 19.8000 37.9000 20.2000 40.2000 ;
	    RECT 21.4000 37.9000 21.8000 40.2000 ;
	    RECT 22.2000 37.9000 22.6000 40.2000 ;
	    RECT 23.8000 38.1000 24.2000 40.2000 ;
	    RECT 26.5000 35.9000 26.9000 40.2000 ;
	    RECT 28.6000 37.9000 29.0000 40.2000 ;
	    RECT 30.2000 38.1000 30.6000 40.2000 ;
	    RECT 32.9000 35.9000 33.3000 40.2000 ;
	    RECT 35.0000 37.9000 35.4000 40.2000 ;
	    RECT 36.6000 37.9000 37.0000 40.2000 ;
	    RECT 38.2000 37.9000 38.6000 40.2000 ;
	    RECT 39.3000 37.9000 39.7000 40.2000 ;
	    RECT 41.4000 35.9000 41.8000 40.2000 ;
	    RECT 43.0000 37.9000 43.4000 40.2000 ;
	    RECT 45.1000 35.9000 45.5000 40.2000 ;
	    RECT 47.8000 38.1000 48.2000 40.2000 ;
	    RECT 49.4000 37.9000 49.8000 40.2000 ;
	    RECT 50.2000 37.9000 50.6000 40.2000 ;
	    RECT 51.8000 37.9000 52.2000 40.2000 ;
	    RECT 53.4000 37.9000 53.8000 40.2000 ;
	    RECT 55.0000 38.1000 55.4000 40.2000 ;
	    RECT 56.6000 37.9000 57.0000 40.2000 ;
	    RECT 57.4000 37.9000 57.8000 40.2000 ;
	    RECT 59.0000 37.9000 59.4000 40.2000 ;
	    RECT 61.4000 35.9000 61.8000 40.2000 ;
	    RECT 63.8000 38.1000 64.2000 40.2000 ;
	    RECT 65.4000 37.9000 65.8000 40.2000 ;
	    RECT 67.0000 38.1000 67.4000 40.2000 ;
	    RECT 68.6000 37.9000 69.0000 40.2000 ;
	    RECT 69.4000 37.9000 69.8000 40.2000 ;
	    RECT 71.0000 38.1000 71.4000 40.2000 ;
	    RECT 73.4000 38.1000 73.8000 40.2000 ;
	    RECT 75.0000 37.9000 75.4000 40.2000 ;
	    RECT 76.1000 37.9000 76.5000 40.2000 ;
	    RECT 78.2000 35.9000 78.6000 40.2000 ;
	    RECT 79.8000 37.9000 80.2000 40.2000 ;
	    RECT 80.6000 35.9000 81.0000 40.2000 ;
	    RECT 82.2000 35.9000 82.6000 40.2000 ;
	    RECT 83.0000 37.9000 83.4000 40.2000 ;
	    RECT 84.6000 37.9000 85.0000 40.2000 ;
	    RECT 86.2000 37.9000 86.6000 40.2000 ;
	    RECT 87.0000 37.9000 87.4000 40.2000 ;
	    RECT 88.6000 37.9000 89.0000 40.2000 ;
	    RECT 90.2000 37.9000 90.6000 40.2000 ;
	    RECT 92.3000 35.9000 92.7000 40.2000 ;
	    RECT 95.0000 38.1000 95.4000 40.2000 ;
	    RECT 96.6000 37.9000 97.0000 40.2000 ;
	    RECT 98.2000 38.1000 98.6000 40.2000 ;
	    RECT 99.8000 37.9000 100.2000 40.2000 ;
	    RECT 101.7000 35.9000 102.1000 40.2000 ;
	    RECT 103.8000 37.9000 104.2000 40.2000 ;
	    RECT 106.2000 38.1000 106.6000 40.2000 ;
	    RECT 107.8000 37.9000 108.2000 40.2000 ;
	    RECT 108.6000 37.9000 109.0000 40.2000 ;
	    RECT 110.2000 38.1000 110.6000 40.2000 ;
	    RECT 114.7000 35.9000 115.1000 40.2000 ;
	    RECT 117.4000 38.1000 117.8000 40.2000 ;
	    RECT 119.0000 37.9000 119.4000 40.2000 ;
	    RECT 119.8000 37.9000 120.2000 40.2000 ;
	    RECT 121.4000 38.1000 121.8000 40.2000 ;
	    RECT 123.0000 35.9000 123.4000 40.2000 ;
	    RECT 124.6000 37.9000 125.0000 40.2000 ;
	    RECT 126.2000 38.1000 126.6000 40.2000 ;
	    RECT 127.8000 37.9000 128.2000 40.2000 ;
	    RECT 130.7000 35.9000 131.1000 40.2000 ;
	    RECT 132.6000 37.9000 133.0000 40.2000 ;
	    RECT 134.2000 37.9000 134.6000 40.2000 ;
	    RECT 135.8000 37.9000 136.2000 40.2000 ;
	    RECT 136.6000 37.9000 137.0000 40.2000 ;
	    RECT 138.2000 38.1000 138.6000 40.2000 ;
	    RECT 139.8000 37.9000 140.2000 40.2000 ;
	    RECT 141.4000 37.9000 141.8000 40.2000 ;
	    RECT 143.0000 38.1000 143.4000 40.2000 ;
	    RECT 144.6000 37.9000 145.0000 40.2000 ;
	    RECT 145.4000 37.9000 145.8000 40.2000 ;
	    RECT 147.0000 38.1000 147.4000 40.2000 ;
	    RECT 149.4000 38.1000 149.8000 40.2000 ;
	    RECT 151.0000 37.9000 151.4000 40.2000 ;
	    RECT 152.6000 35.9000 153.0000 40.2000 ;
	    RECT 153.4000 37.9000 153.8000 40.2000 ;
	    RECT 155.0000 38.1000 155.4000 40.2000 ;
	    RECT 157.4000 36.5000 157.8000 40.2000 ;
	    RECT 159.8000 36.5000 160.2000 40.2000 ;
	    RECT 161.4000 37.9000 161.8000 40.2000 ;
	    RECT 163.0000 38.1000 163.4000 40.2000 ;
	    RECT 164.6000 37.9000 165.0000 40.2000 ;
	    RECT 166.2000 38.1000 166.6000 40.2000 ;
	    RECT 167.8000 37.9000 168.2000 40.2000 ;
	    RECT 169.4000 37.9000 169.8000 40.2000 ;
	    RECT 171.0000 37.9000 171.4000 40.2000 ;
	    RECT 0.6000 20.8000 1.0000 23.1000 ;
	    RECT 2.2000 20.8000 2.6000 23.1000 ;
	    RECT 3.8000 20.8000 4.2000 23.1000 ;
	    RECT 5.7000 20.8000 6.1000 25.1000 ;
	    RECT 8.6000 20.8000 9.0000 22.9000 ;
	    RECT 10.2000 20.8000 10.6000 23.1000 ;
	    RECT 11.8000 20.8000 12.2000 24.5000 ;
	    RECT 13.4000 20.8000 13.8000 23.1000 ;
	    RECT 15.0000 20.8000 15.4000 22.9000 ;
	    RECT 16.6000 20.8000 17.0000 23.1000 ;
	    RECT 18.2000 20.8000 18.6000 22.9000 ;
	    RECT 20.6000 20.8000 21.0000 24.5000 ;
	    RECT 22.2000 20.8000 22.6000 23.1000 ;
	    RECT 23.8000 20.8000 24.2000 22.9000 ;
	    RECT 26.5000 20.8000 26.9000 25.1000 ;
	    RECT 29.4000 20.8000 29.8000 24.5000 ;
	    RECT 31.0000 20.8000 31.4000 23.1000 ;
	    RECT 32.6000 20.8000 33.0000 23.1000 ;
	    RECT 33.4000 20.8000 33.8000 23.1000 ;
	    RECT 35.0000 20.8000 35.4000 22.9000 ;
	    RECT 37.7000 20.8000 38.1000 25.1000 ;
	    RECT 40.6000 20.8000 41.0000 23.1000 ;
	    RECT 41.4000 20.8000 41.8000 23.1000 ;
	    RECT 43.0000 20.8000 43.4000 23.1000 ;
	    RECT 44.6000 20.8000 45.0000 23.1000 ;
	    RECT 45.4000 20.8000 45.8000 23.1000 ;
	    RECT 47.0000 20.8000 47.4000 23.1000 ;
	    RECT 48.6000 20.8000 49.0000 23.1000 ;
	    RECT 50.7000 20.8000 51.1000 25.1000 ;
	    RECT 53.4000 20.8000 53.8000 22.9000 ;
	    RECT 55.0000 20.8000 55.4000 23.1000 ;
	    RECT 56.6000 20.8000 57.0000 22.9000 ;
	    RECT 58.2000 20.8000 58.6000 23.1000 ;
	    RECT 59.8000 20.8000 60.2000 24.5000 ;
	    RECT 63.0000 20.8000 63.4000 23.1000 ;
	    RECT 64.6000 20.8000 65.0000 23.1000 ;
	    RECT 65.4000 20.8000 65.8000 23.1000 ;
	    RECT 67.0000 20.8000 67.4000 23.1000 ;
	    RECT 68.6000 20.8000 69.0000 24.5000 ;
	    RECT 71.5000 20.8000 71.9000 25.1000 ;
	    RECT 73.4000 20.8000 73.8000 23.1000 ;
	    RECT 75.0000 20.8000 75.4000 22.9000 ;
	    RECT 76.6000 20.8000 77.0000 23.1000 ;
	    RECT 78.2000 20.8000 78.6000 23.1000 ;
	    RECT 79.8000 20.8000 80.2000 24.5000 ;
	    RECT 81.4000 20.8000 81.8000 23.1000 ;
	    RECT 83.0000 20.8000 83.4000 22.9000 ;
	    RECT 85.9000 20.8000 86.3000 25.1000 ;
	    RECT 87.8000 20.8000 88.2000 23.1000 ;
	    RECT 89.4000 20.8000 89.8000 23.1000 ;
	    RECT 91.0000 20.8000 91.4000 23.1000 ;
	    RECT 92.6000 20.8000 93.0000 23.1000 ;
	    RECT 94.2000 20.8000 94.6000 22.9000 ;
	    RECT 95.8000 20.8000 96.2000 23.1000 ;
	    RECT 97.4000 20.8000 97.8000 22.9000 ;
	    RECT 99.0000 20.8000 99.4000 23.1000 ;
	    RECT 99.8000 20.8000 100.2000 23.1000 ;
	    RECT 101.4000 20.8000 101.8000 22.9000 ;
	    RECT 103.0000 20.8000 103.4000 23.1000 ;
	    RECT 104.6000 20.8000 105.0000 23.1000 ;
	    RECT 106.2000 20.8000 106.6000 23.1000 ;
	    RECT 107.0000 20.8000 107.4000 23.1000 ;
	    RECT 108.6000 20.8000 109.0000 22.9000 ;
	    RECT 111.0000 20.8000 111.4000 24.5000 ;
	    RECT 114.2000 20.8000 114.6000 23.1000 ;
	    RECT 115.8000 20.8000 116.2000 23.1000 ;
	    RECT 116.6000 20.8000 117.0000 23.1000 ;
	    RECT 118.2000 20.8000 118.6000 23.1000 ;
	    RECT 120.3000 20.8000 120.7000 25.1000 ;
	    RECT 123.0000 20.8000 123.4000 22.9000 ;
	    RECT 124.6000 20.8000 125.0000 23.1000 ;
	    RECT 125.4000 20.8000 125.8000 23.1000 ;
	    RECT 127.0000 20.8000 127.4000 23.1000 ;
	    RECT 129.1000 20.8000 129.5000 25.1000 ;
	    RECT 131.8000 20.8000 132.2000 22.9000 ;
	    RECT 133.4000 20.8000 133.8000 23.1000 ;
	    RECT 134.2000 20.8000 134.6000 23.1000 ;
	    RECT 135.8000 20.8000 136.2000 22.9000 ;
	    RECT 137.4000 20.8000 137.8000 23.1000 ;
	    RECT 139.0000 20.8000 139.4000 23.1000 ;
	    RECT 141.1000 20.8000 141.5000 25.1000 ;
	    RECT 143.8000 20.8000 144.2000 22.9000 ;
	    RECT 145.4000 20.8000 145.8000 23.1000 ;
	    RECT 146.2000 20.8000 146.6000 25.1000 ;
	    RECT 147.8000 20.8000 148.2000 25.1000 ;
	    RECT 148.6000 20.8000 149.0000 23.1000 ;
	    RECT 150.2000 20.8000 150.6000 23.1000 ;
	    RECT 151.0000 20.8000 151.4000 23.1000 ;
	    RECT 152.6000 20.8000 153.0000 22.9000 ;
	    RECT 154.2000 20.8000 154.6000 23.1000 ;
	    RECT 155.8000 20.8000 156.2000 23.1000 ;
	    RECT 157.4000 20.8000 157.8000 24.5000 ;
	    RECT 159.8000 20.8000 160.2000 25.0000 ;
	    RECT 162.6000 20.8000 163.0000 23.1000 ;
	    RECT 164.2000 20.8000 164.6000 23.1000 ;
	    RECT 167.0000 20.8000 167.4000 25.1000 ;
	    RECT 169.9000 20.8000 170.3000 25.1000 ;
	    RECT 0.2000 20.2000 173.4000 20.8000 ;
	    RECT 0.6000 15.9000 1.0000 20.2000 ;
	    RECT 2.2000 15.9000 2.6000 20.2000 ;
	    RECT 3.8000 18.1000 4.2000 20.2000 ;
	    RECT 5.4000 17.9000 5.8000 20.2000 ;
	    RECT 7.3000 15.9000 7.7000 20.2000 ;
	    RECT 10.2000 18.1000 10.6000 20.2000 ;
	    RECT 11.8000 17.9000 12.2000 20.2000 ;
	    RECT 13.4000 15.9000 13.8000 20.2000 ;
	    RECT 14.2000 17.9000 14.6000 20.2000 ;
	    RECT 15.8000 18.1000 16.2000 20.2000 ;
	    RECT 17.4000 17.9000 17.8000 20.2000 ;
	    RECT 19.0000 18.1000 19.4000 20.2000 ;
	    RECT 20.6000 17.9000 21.0000 20.2000 ;
	    RECT 22.2000 17.9000 22.6000 20.2000 ;
	    RECT 23.0000 17.9000 23.4000 20.2000 ;
	    RECT 24.6000 18.1000 25.0000 20.2000 ;
	    RECT 26.2000 17.9000 26.6000 20.2000 ;
	    RECT 27.8000 18.1000 28.2000 20.2000 ;
	    RECT 30.2000 16.5000 30.6000 20.2000 ;
	    RECT 31.8000 17.9000 32.2000 20.2000 ;
	    RECT 33.4000 18.1000 33.8000 20.2000 ;
	    RECT 36.1000 15.9000 36.5000 20.2000 ;
	    RECT 39.3000 15.9000 39.7000 20.2000 ;
	    RECT 42.5000 15.9000 42.9000 20.2000 ;
	    RECT 44.6000 15.9000 45.0000 20.2000 ;
	    RECT 46.7000 17.9000 47.1000 20.2000 ;
	    RECT 48.6000 17.9000 49.0000 20.2000 ;
	    RECT 50.2000 18.1000 50.6000 20.2000 ;
	    RECT 51.8000 17.9000 52.2000 20.2000 ;
	    RECT 53.7000 15.9000 54.1000 20.2000 ;
	    RECT 56.1000 17.9000 56.5000 20.2000 ;
	    RECT 58.2000 15.9000 58.6000 20.2000 ;
	    RECT 59.8000 17.9000 60.2000 20.2000 ;
	    RECT 62.2000 17.9000 62.6000 20.2000 ;
	    RECT 63.8000 15.9000 64.2000 20.2000 ;
	    RECT 65.9000 17.9000 66.3000 20.2000 ;
	    RECT 67.8000 18.1000 68.2000 20.2000 ;
	    RECT 69.4000 17.9000 69.8000 20.2000 ;
	    RECT 71.5000 15.9000 71.9000 20.2000 ;
	    RECT 73.7000 17.9000 74.1000 20.2000 ;
	    RECT 75.8000 15.9000 76.2000 20.2000 ;
	    RECT 77.4000 17.9000 77.8000 20.2000 ;
	    RECT 79.5000 15.9000 79.9000 20.2000 ;
	    RECT 81.4000 17.9000 81.8000 20.2000 ;
	    RECT 83.0000 18.1000 83.4000 20.2000 ;
	    RECT 84.6000 17.9000 85.0000 20.2000 ;
	    RECT 86.2000 18.1000 86.6000 20.2000 ;
	    RECT 88.9000 15.9000 89.3000 20.2000 ;
	    RECT 91.0000 17.9000 91.4000 20.2000 ;
	    RECT 92.6000 18.1000 93.0000 20.2000 ;
	    RECT 95.3000 15.9000 95.7000 20.2000 ;
	    RECT 97.4000 17.9000 97.8000 20.2000 ;
	    RECT 99.0000 17.9000 99.4000 20.2000 ;
	    RECT 100.6000 17.9000 101.0000 20.2000 ;
	    RECT 102.2000 18.1000 102.6000 20.2000 ;
	    RECT 103.8000 17.9000 104.2000 20.2000 ;
	    RECT 105.9000 15.9000 106.3000 20.2000 ;
	    RECT 108.6000 18.1000 109.0000 20.2000 ;
	    RECT 110.2000 17.9000 110.6000 20.2000 ;
	    RECT 113.4000 18.1000 113.8000 20.2000 ;
	    RECT 115.0000 17.9000 115.4000 20.2000 ;
	    RECT 116.9000 15.9000 117.3000 20.2000 ;
	    RECT 120.1000 15.9000 120.5000 20.2000 ;
	    RECT 123.0000 18.1000 123.4000 20.2000 ;
	    RECT 124.6000 17.9000 125.0000 20.2000 ;
	    RECT 126.2000 18.1000 126.6000 20.2000 ;
	    RECT 127.8000 17.9000 128.2000 20.2000 ;
	    RECT 129.4000 16.5000 129.8000 20.2000 ;
	    RECT 132.1000 15.9000 132.5000 20.2000 ;
	    RECT 135.3000 15.9000 135.7000 20.2000 ;
	    RECT 137.4000 17.9000 137.8000 20.2000 ;
	    RECT 139.3000 17.9000 139.7000 20.2000 ;
	    RECT 141.4000 15.9000 141.8000 20.2000 ;
	    RECT 142.5000 17.9000 142.9000 20.2000 ;
	    RECT 144.6000 15.9000 145.0000 20.2000 ;
	    RECT 146.2000 17.9000 146.6000 20.2000 ;
	    RECT 147.8000 18.1000 148.2000 20.2000 ;
	    RECT 149.4000 17.9000 149.8000 20.2000 ;
	    RECT 151.3000 15.9000 151.7000 20.2000 ;
	    RECT 153.7000 17.9000 154.1000 20.2000 ;
	    RECT 155.8000 15.9000 156.2000 20.2000 ;
	    RECT 156.6000 17.9000 157.0000 20.2000 ;
	    RECT 158.2000 17.9000 158.6000 20.2000 ;
	    RECT 159.8000 18.1000 160.2000 20.2000 ;
	    RECT 161.4000 17.9000 161.8000 20.2000 ;
	    RECT 163.0000 18.1000 163.4000 20.2000 ;
	    RECT 164.9000 17.9000 165.3000 20.2000 ;
	    RECT 167.0000 15.9000 167.4000 20.2000 ;
	    RECT 168.6000 17.9000 169.0000 20.2000 ;
	    RECT 170.2000 16.5000 170.6000 20.2000 ;
	    RECT 0.6000 0.8000 1.0000 3.1000 ;
	    RECT 2.2000 0.8000 2.6000 3.1000 ;
	    RECT 3.0000 0.8000 3.4000 3.1000 ;
	    RECT 4.6000 0.8000 5.0000 3.1000 ;
	    RECT 5.4000 0.8000 5.8000 3.1000 ;
	    RECT 7.0000 0.8000 7.4000 3.1000 ;
	    RECT 8.1000 0.8000 8.5000 3.1000 ;
	    RECT 10.2000 0.8000 10.6000 5.1000 ;
	    RECT 11.8000 0.8000 12.2000 3.1000 ;
	    RECT 13.9000 0.8000 14.3000 5.1000 ;
	    RECT 16.6000 0.8000 17.0000 3.1000 ;
	    RECT 17.4000 0.8000 17.8000 3.1000 ;
	    RECT 19.0000 0.8000 19.4000 3.1000 ;
	    RECT 20.6000 0.8000 21.0000 4.5000 ;
	    RECT 22.2000 0.8000 22.6000 3.1000 ;
	    RECT 23.8000 0.8000 24.2000 3.1000 ;
	    RECT 25.4000 0.8000 25.8000 3.1000 ;
	    RECT 26.2000 0.8000 26.6000 3.1000 ;
	    RECT 27.8000 0.8000 28.2000 3.1000 ;
	    RECT 28.6000 0.8000 29.0000 3.1000 ;
	    RECT 30.2000 0.8000 30.6000 3.1000 ;
	    RECT 31.8000 0.8000 32.2000 3.1000 ;
	    RECT 32.6000 0.8000 33.0000 3.1000 ;
	    RECT 34.2000 0.8000 34.6000 3.1000 ;
	    RECT 35.0000 0.8000 35.4000 3.1000 ;
	    RECT 36.6000 0.8000 37.0000 3.1000 ;
	    RECT 37.4000 0.8000 37.8000 3.1000 ;
	    RECT 39.0000 0.8000 39.4000 3.1000 ;
	    RECT 40.1000 0.8000 40.5000 3.1000 ;
	    RECT 42.2000 0.8000 42.6000 5.1000 ;
	    RECT 43.8000 0.8000 44.2000 3.1000 ;
	    RECT 45.4000 0.8000 45.8000 3.1000 ;
	    RECT 46.2000 0.8000 46.6000 3.1000 ;
	    RECT 47.8000 0.8000 48.2000 3.1000 ;
	    RECT 49.4000 0.8000 49.8000 3.1000 ;
	    RECT 51.0000 0.8000 51.4000 3.1000 ;
	    RECT 51.8000 0.8000 52.2000 3.1000 ;
	    RECT 53.4000 0.8000 53.8000 3.1000 ;
	    RECT 54.2000 0.8000 54.6000 3.1000 ;
	    RECT 55.8000 0.8000 56.2000 3.1000 ;
	    RECT 56.6000 0.8000 57.0000 3.1000 ;
	    RECT 58.2000 0.8000 58.6000 3.1000 ;
	    RECT 59.8000 0.8000 60.2000 4.5000 ;
	    RECT 63.0000 0.8000 63.4000 3.1000 ;
	    RECT 64.6000 0.8000 65.0000 3.1000 ;
	    RECT 65.4000 0.8000 65.8000 3.1000 ;
	    RECT 67.8000 0.8000 68.2000 3.1000 ;
	    RECT 68.6000 0.8000 69.0000 3.1000 ;
	    RECT 70.2000 0.8000 70.6000 3.1000 ;
	    RECT 71.0000 0.8000 71.4000 3.1000 ;
	    RECT 72.6000 0.8000 73.0000 3.1000 ;
	    RECT 74.2000 0.8000 74.6000 3.1000 ;
	    RECT 75.0000 0.8000 75.4000 3.1000 ;
	    RECT 76.6000 0.8000 77.0000 3.1000 ;
	    RECT 78.2000 0.8000 78.6000 3.1000 ;
	    RECT 79.8000 0.8000 80.2000 4.5000 ;
	    RECT 81.4000 0.8000 81.8000 3.1000 ;
	    RECT 83.0000 0.8000 83.4000 3.1000 ;
	    RECT 84.6000 0.8000 85.0000 3.1000 ;
	    RECT 85.4000 0.8000 85.8000 3.1000 ;
	    RECT 87.0000 0.8000 87.4000 3.1000 ;
	    RECT 88.6000 0.8000 89.0000 3.1000 ;
	    RECT 89.4000 0.8000 89.8000 3.1000 ;
	    RECT 91.0000 0.8000 91.4000 3.1000 ;
	    RECT 92.6000 0.8000 93.0000 3.1000 ;
	    RECT 93.4000 0.8000 93.8000 3.1000 ;
	    RECT 95.0000 0.8000 95.4000 3.1000 ;
	    RECT 95.8000 0.8000 96.2000 3.1000 ;
	    RECT 97.7000 0.8000 98.1000 3.1000 ;
	    RECT 99.8000 0.8000 100.2000 5.1000 ;
	    RECT 100.6000 0.8000 101.0000 3.1000 ;
	    RECT 102.2000 0.8000 102.6000 3.1000 ;
	    RECT 103.0000 0.8000 103.4000 3.1000 ;
	    RECT 104.6000 0.8000 105.0000 3.1000 ;
	    RECT 106.2000 0.8000 106.6000 3.1000 ;
	    RECT 107.0000 0.8000 107.4000 3.1000 ;
	    RECT 108.6000 0.8000 109.0000 3.1000 ;
	    RECT 110.2000 0.8000 110.6000 3.1000 ;
	    RECT 112.6000 0.8000 113.0000 3.1000 ;
	    RECT 114.2000 0.8000 114.6000 3.1000 ;
	    RECT 115.3000 0.8000 115.7000 3.1000 ;
	    RECT 117.4000 0.8000 117.8000 5.1000 ;
	    RECT 119.0000 0.8000 119.4000 3.1000 ;
	    RECT 120.6000 0.8000 121.0000 4.5000 ;
	    RECT 122.2000 0.8000 122.6000 3.1000 ;
	    RECT 123.8000 0.8000 124.2000 3.1000 ;
	    RECT 124.6000 0.8000 125.0000 3.1000 ;
	    RECT 126.2000 0.8000 126.6000 3.1000 ;
	    RECT 127.8000 0.8000 128.2000 3.1000 ;
	    RECT 128.6000 0.8000 129.0000 3.1000 ;
	    RECT 130.2000 0.8000 130.6000 3.1000 ;
	    RECT 131.8000 0.8000 132.2000 3.1000 ;
	    RECT 133.4000 0.8000 133.8000 3.1000 ;
	    RECT 134.2000 0.8000 134.6000 3.1000 ;
	    RECT 135.8000 0.8000 136.2000 3.1000 ;
	    RECT 137.4000 0.8000 137.8000 3.1000 ;
	    RECT 138.2000 0.8000 138.6000 3.1000 ;
	    RECT 139.8000 0.8000 140.2000 3.1000 ;
	    RECT 140.6000 0.8000 141.0000 3.1000 ;
	    RECT 142.2000 0.8000 142.6000 3.1000 ;
	    RECT 143.0000 0.8000 143.4000 3.1000 ;
	    RECT 144.6000 0.8000 145.0000 3.1000 ;
	    RECT 146.2000 0.8000 146.6000 3.1000 ;
	    RECT 147.0000 0.8000 147.4000 3.1000 ;
	    RECT 148.6000 0.8000 149.0000 3.1000 ;
	    RECT 149.4000 0.8000 149.8000 3.1000 ;
	    RECT 151.0000 0.8000 151.4000 3.1000 ;
	    RECT 153.1000 0.8000 153.5000 5.1000 ;
	    RECT 156.3000 0.8000 156.7000 5.1000 ;
	    RECT 159.0000 0.8000 159.4000 5.1000 ;
	    RECT 159.8000 0.8000 160.2000 5.1000 ;
	    RECT 161.4000 0.8000 161.8000 5.1000 ;
	    RECT 163.0000 0.8000 163.4000 5.1000 ;
	    RECT 164.6000 0.8000 165.0000 5.1000 ;
	    RECT 166.2000 0.8000 166.6000 5.1000 ;
	    RECT 167.8000 0.8000 168.2000 4.5000 ;
	    RECT 169.4000 0.8000 169.8000 3.1000 ;
	    RECT 171.0000 0.8000 171.4000 4.9000 ;
	    RECT 0.2000 0.2000 173.4000 0.8000 ;
         LAYER metal2 ;
	    RECT 60.0000 160.3000 61.6000 160.7000 ;
	    RECT 60.0000 140.3000 61.6000 140.7000 ;
	    RECT 60.0000 120.3000 61.6000 120.7000 ;
	    RECT 60.0000 100.3000 61.6000 100.7000 ;
	    RECT 60.0000 80.3000 61.6000 80.7000 ;
	    RECT 60.0000 60.3000 61.6000 60.7000 ;
	    RECT 60.0000 40.3000 61.6000 40.7000 ;
	    RECT 60.0000 20.3000 61.6000 20.7000 ;
	    RECT 60.0000 0.3000 61.6000 0.7000 ;
         LAYER metal3 ;
	    RECT 60.0000 160.3000 61.6000 160.7000 ;
	    RECT 60.0000 140.3000 61.6000 140.7000 ;
	    RECT 60.0000 120.3000 61.6000 120.7000 ;
	    RECT 60.0000 100.3000 61.6000 100.7000 ;
	    RECT 60.0000 80.3000 61.6000 80.7000 ;
	    RECT 60.0000 60.3000 61.6000 60.7000 ;
	    RECT 60.0000 40.3000 61.6000 40.7000 ;
	    RECT 60.0000 20.3000 61.6000 20.7000 ;
	    RECT 60.0000 0.3000 61.6000 0.7000 ;
         LAYER metal4 ;
	    RECT 60.0000 160.3000 61.6000 160.7000 ;
	    RECT 60.0000 140.3000 61.6000 140.7000 ;
	    RECT 60.0000 120.3000 61.6000 120.7000 ;
	    RECT 60.0000 100.3000 61.6000 100.7000 ;
	    RECT 60.0000 80.3000 61.6000 80.7000 ;
	    RECT 60.0000 60.3000 61.6000 60.7000 ;
	    RECT 60.0000 40.3000 61.6000 40.7000 ;
	    RECT 60.0000 20.3000 61.6000 20.7000 ;
	    RECT 60.0000 0.3000 61.6000 0.7000 ;
         LAYER metal5 ;
	    RECT 60.0000 160.7000 60.6000 160.8000 ;
	    RECT 61.0000 160.7000 61.6000 160.8000 ;
	    RECT 60.0000 160.2000 61.6000 160.7000 ;
	    RECT 60.0000 140.7000 60.6000 140.8000 ;
	    RECT 61.0000 140.7000 61.6000 140.8000 ;
	    RECT 60.0000 140.2000 61.6000 140.7000 ;
	    RECT 60.0000 120.7000 60.6000 120.8000 ;
	    RECT 61.0000 120.7000 61.6000 120.8000 ;
	    RECT 60.0000 120.2000 61.6000 120.7000 ;
	    RECT 60.0000 100.7000 60.6000 100.8000 ;
	    RECT 61.0000 100.7000 61.6000 100.8000 ;
	    RECT 60.0000 100.2000 61.6000 100.7000 ;
	    RECT 60.0000 80.7000 60.6000 80.8000 ;
	    RECT 61.0000 80.7000 61.6000 80.8000 ;
	    RECT 60.0000 80.2000 61.6000 80.7000 ;
	    RECT 60.0000 60.7000 60.6000 60.8000 ;
	    RECT 61.0000 60.7000 61.6000 60.8000 ;
	    RECT 60.0000 60.2000 61.6000 60.7000 ;
	    RECT 60.0000 40.7000 60.6000 40.8000 ;
	    RECT 61.0000 40.7000 61.6000 40.8000 ;
	    RECT 60.0000 40.2000 61.6000 40.7000 ;
	    RECT 60.0000 20.7000 60.6000 20.8000 ;
	    RECT 61.0000 20.7000 61.6000 20.8000 ;
	    RECT 60.0000 20.2000 61.6000 20.7000 ;
	    RECT 60.0000 0.7000 60.6000 0.8000 ;
	    RECT 61.0000 0.7000 61.6000 0.8000 ;
	    RECT 60.0000 0.2000 61.6000 0.7000 ;
         LAYER metal6 ;
	    RECT 60.0000 -3.0000 61.6000 164.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 0.6000 150.8000 1.0000 152.1000 ;
	    RECT 3.8000 150.8000 4.2000 153.1000 ;
	    RECT 4.6000 150.8000 5.0000 153.1000 ;
	    RECT 7.8000 150.8000 8.2000 152.1000 ;
	    RECT 9.4000 150.8000 9.8000 152.7000 ;
	    RECT 13.4000 150.8000 13.8000 153.1000 ;
	    RECT 14.2000 150.8000 14.6000 153.1000 ;
	    RECT 17.4000 150.8000 17.8000 153.1000 ;
	    RECT 19.0000 150.8000 19.4000 153.1000 ;
	    RECT 21.4000 150.8000 21.8000 153.1000 ;
	    RECT 24.6000 150.8000 25.0000 152.1000 ;
	    RECT 25.4000 150.8000 25.8000 153.1000 ;
	    RECT 27.8000 150.8000 28.2000 152.1000 ;
	    RECT 30.2000 150.8000 30.6000 152.1000 ;
	    RECT 31.0000 150.8000 31.4000 152.1000 ;
	    RECT 33.4000 150.8000 33.8000 152.7000 ;
	    RECT 37.4000 150.8000 37.8000 153.1000 ;
	    RECT 39.8000 150.8000 40.2000 153.1000 ;
	    RECT 41.4000 150.8000 41.8000 153.1000 ;
	    RECT 43.0000 150.8000 43.4000 153.1000 ;
	    RECT 45.4000 150.8000 45.8000 153.1000 ;
	    RECT 48.6000 150.8000 49.0000 152.1000 ;
	    RECT 51.0000 150.8000 51.4000 153.1000 ;
	    RECT 51.8000 150.8000 52.2000 153.1000 ;
	    RECT 55.0000 150.8000 55.4000 153.1000 ;
	    RECT 56.6000 150.8000 57.0000 152.1000 ;
	    RECT 59.0000 150.8000 59.4000 152.7000 ;
	    RECT 64.6000 150.8000 65.0000 153.1000 ;
	    RECT 65.4000 150.8000 65.8000 153.1000 ;
	    RECT 68.6000 150.8000 69.0000 152.1000 ;
	    RECT 71.0000 150.8000 71.4000 153.1000 ;
	    RECT 71.8000 150.8000 72.2000 153.1000 ;
	    RECT 75.0000 150.8000 75.4000 152.1000 ;
	    RECT 75.8000 150.8000 76.2000 152.1000 ;
	    RECT 77.4000 150.8000 77.8000 152.1000 ;
	    RECT 79.8000 150.8000 80.2000 153.1000 ;
	    RECT 81.4000 150.8000 81.8000 153.0000 ;
	    RECT 84.2000 150.8000 84.6000 152.1000 ;
	    RECT 85.8000 150.8000 86.3000 152.1000 ;
	    RECT 88.6000 150.8000 89.0000 153.1000 ;
	    RECT 91.0000 150.8000 91.4000 153.1000 ;
	    RECT 92.6000 150.8000 93.0000 152.7000 ;
	    RECT 96.6000 150.8000 97.0000 152.7000 ;
	    RECT 99.8000 150.8000 100.2000 152.1000 ;
	    RECT 101.4000 150.8000 101.8000 152.1000 ;
	    RECT 102.2000 150.8000 102.6000 153.1000 ;
	    RECT 104.6000 150.8000 105.0000 152.1000 ;
	    RECT 106.7000 150.8000 107.1000 153.1000 ;
	    RECT 109.4000 150.8000 109.8000 153.1000 ;
	    RECT 110.2000 150.8000 110.6000 152.1000 ;
	    RECT 111.8000 150.8000 112.2000 152.1000 ;
	    RECT 114.2000 150.8000 114.6000 152.1000 ;
	    RECT 115.8000 150.8000 116.2000 153.1000 ;
	    RECT 118.4000 150.8000 118.8000 153.1000 ;
	    RECT 121.4000 150.8000 121.8000 153.1000 ;
	    RECT 123.0000 150.8000 123.4000 152.1000 ;
	    RECT 124.6000 150.8000 125.0000 151.9000 ;
	    RECT 128.6000 150.8000 129.0000 152.1000 ;
	    RECT 131.8000 150.8000 132.2000 152.7000 ;
	    RECT 133.4000 150.8000 133.8000 152.1000 ;
	    RECT 135.5000 150.8000 135.9000 153.1000 ;
	    RECT 138.2000 150.8000 138.6000 152.7000 ;
	    RECT 139.8000 150.8000 140.2000 152.1000 ;
	    RECT 141.4000 150.8000 141.8000 152.1000 ;
	    RECT 142.2000 150.8000 142.6000 152.1000 ;
	    RECT 144.3000 150.8000 144.7000 153.1000 ;
	    RECT 147.0000 150.8000 147.4000 153.1000 ;
	    RECT 147.8000 150.8000 148.2000 154.1000 ;
	    RECT 153.4000 150.8000 153.8000 154.1000 ;
	    RECT 154.2000 150.8000 154.6000 153.1000 ;
	    RECT 157.4000 150.8000 157.8000 152.7000 ;
	    RECT 159.8000 150.8000 160.2000 153.1000 ;
	    RECT 163.0000 150.8000 163.4000 153.1000 ;
	    RECT 165.7000 150.8000 166.2000 152.1000 ;
	    RECT 167.4000 150.8000 167.8000 152.1000 ;
	    RECT 170.2000 150.8000 170.6000 153.0000 ;
	    RECT 0.2000 150.2000 173.4000 150.8000 ;
	    RECT 3.0000 146.9000 3.4000 150.2000 ;
	    RECT 4.6000 148.1000 5.0000 150.2000 ;
	    RECT 6.2000 148.9000 6.6000 150.2000 ;
	    RECT 8.6000 148.3000 9.0000 150.2000 ;
	    RECT 11.0000 148.9000 11.4000 150.2000 ;
	    RECT 12.6000 147.9000 13.0000 150.2000 ;
	    RECT 15.8000 148.3000 16.2000 150.2000 ;
	    RECT 18.2000 148.9000 18.6000 150.2000 ;
	    RECT 19.8000 148.9000 20.2000 150.2000 ;
	    RECT 20.6000 146.9000 21.0000 150.2000 ;
	    RECT 24.6000 148.1000 25.0000 150.2000 ;
	    RECT 26.2000 148.9000 26.6000 150.2000 ;
	    RECT 28.6000 148.3000 29.0000 150.2000 ;
	    RECT 31.0000 148.9000 31.4000 150.2000 ;
	    RECT 33.4000 148.3000 33.8000 150.2000 ;
	    RECT 35.8000 148.9000 36.2000 150.2000 ;
	    RECT 37.4000 148.3000 37.8000 150.2000 ;
	    RECT 40.6000 147.9000 41.0000 150.2000 ;
	    RECT 42.2000 148.9000 42.6000 150.2000 ;
	    RECT 44.6000 148.3000 45.0000 150.2000 ;
	    RECT 47.0000 148.9000 47.4000 150.2000 ;
	    RECT 48.6000 148.1000 49.0000 150.2000 ;
	    RECT 50.2000 148.9000 50.6000 150.2000 ;
	    RECT 54.2000 146.9000 54.6000 150.2000 ;
	    RECT 55.0000 148.9000 55.4000 150.2000 ;
	    RECT 59.0000 146.9000 59.4000 150.2000 ;
	    RECT 61.4000 148.9000 61.8000 150.2000 ;
	    RECT 63.0000 148.1000 63.4000 150.2000 ;
	    RECT 64.6000 146.9000 65.0000 150.2000 ;
	    RECT 67.8000 146.9000 68.2000 150.2000 ;
	    RECT 71.0000 148.9000 71.4000 150.2000 ;
	    RECT 72.9000 147.9000 73.3000 150.2000 ;
	    RECT 75.0000 148.9000 75.4000 150.2000 ;
	    RECT 75.8000 148.9000 76.2000 150.2000 ;
	    RECT 77.4000 148.9000 77.8000 150.2000 ;
	    RECT 78.2000 147.9000 78.6000 150.2000 ;
	    RECT 80.6000 146.9000 81.0000 150.2000 ;
	    RECT 83.8000 148.9000 84.2000 150.2000 ;
	    RECT 85.4000 147.9000 85.8000 150.2000 ;
	    RECT 87.2000 147.9000 87.6000 150.2000 ;
	    RECT 90.2000 147.9000 90.6000 150.2000 ;
	    RECT 91.8000 147.9000 92.2000 150.2000 ;
	    RECT 95.0000 146.9000 95.4000 150.2000 ;
	    RECT 95.8000 147.9000 96.2000 150.2000 ;
	    RECT 98.2000 148.9000 98.6000 150.2000 ;
	    RECT 99.8000 148.9000 100.2000 150.2000 ;
	    RECT 103.0000 146.9000 103.4000 150.2000 ;
	    RECT 103.8000 147.9000 104.2000 150.2000 ;
	    RECT 105.4000 147.9000 105.8000 150.2000 ;
	    RECT 107.8000 148.3000 108.2000 150.2000 ;
	    RECT 111.0000 148.3000 111.4000 150.2000 ;
	    RECT 116.6000 146.9000 117.0000 150.2000 ;
	    RECT 118.2000 148.3000 118.6000 150.2000 ;
	    RECT 122.2000 148.3000 122.6000 150.2000 ;
	    RECT 123.8000 146.9000 124.2000 150.2000 ;
	    RECT 127.0000 148.9000 127.4000 150.2000 ;
	    RECT 129.1000 147.9000 129.5000 150.2000 ;
	    RECT 131.8000 148.3000 132.2000 150.2000 ;
	    RECT 136.6000 149.1000 137.0000 150.2000 ;
	    RECT 138.2000 148.9000 138.6000 150.2000 ;
	    RECT 140.6000 148.3000 141.0000 150.2000 ;
	    RECT 143.0000 147.9000 143.4000 150.2000 ;
	    RECT 146.0000 147.9000 146.4000 150.2000 ;
	    RECT 147.0000 147.9000 147.4000 150.2000 ;
	    RECT 150.0000 147.9000 150.4000 150.2000 ;
	    RECT 151.0000 148.9000 151.4000 150.2000 ;
	    RECT 152.6000 148.9000 153.0000 150.2000 ;
	    RECT 153.4000 146.9000 153.8000 150.2000 ;
	    RECT 157.4000 148.3000 157.8000 150.2000 ;
	    RECT 159.8000 148.9000 160.2000 150.2000 ;
	    RECT 161.4000 148.9000 161.8000 150.2000 ;
	    RECT 163.0000 147.9000 163.4000 150.2000 ;
	    RECT 165.7000 148.9000 166.2000 150.2000 ;
	    RECT 167.4000 148.9000 167.8000 150.2000 ;
	    RECT 170.2000 148.0000 170.6000 150.2000 ;
	    RECT 1.4000 130.8000 1.8000 133.1000 ;
	    RECT 3.0000 130.8000 3.4000 133.1000 ;
	    RECT 5.4000 130.8000 5.8000 132.1000 ;
	    RECT 7.0000 130.8000 7.4000 132.9000 ;
	    RECT 8.6000 130.8000 9.0000 134.1000 ;
	    RECT 11.8000 130.8000 12.2000 133.1000 ;
	    RECT 15.8000 130.8000 16.2000 133.1000 ;
	    RECT 18.2000 130.8000 18.6000 133.1000 ;
	    RECT 20.6000 130.8000 21.0000 133.1000 ;
	    RECT 21.4000 130.8000 21.8000 133.1000 ;
	    RECT 24.6000 130.8000 25.0000 133.1000 ;
	    RECT 27.0000 130.8000 27.4000 132.1000 ;
	    RECT 29.4000 130.8000 29.8000 133.1000 ;
	    RECT 30.2000 130.8000 30.6000 133.1000 ;
	    RECT 32.6000 130.8000 33.0000 132.1000 ;
	    RECT 34.2000 130.8000 34.6000 132.9000 ;
	    RECT 35.8000 130.8000 36.2000 133.1000 ;
	    RECT 38.2000 130.8000 38.6000 132.1000 ;
	    RECT 40.6000 130.8000 41.0000 132.7000 ;
	    RECT 43.0000 130.8000 43.4000 133.1000 ;
	    RECT 45.4000 130.8000 45.8000 132.1000 ;
	    RECT 47.8000 130.8000 48.2000 132.7000 ;
	    RECT 51.8000 130.8000 52.2000 133.1000 ;
	    RECT 54.2000 130.8000 54.6000 133.1000 ;
	    RECT 56.6000 130.8000 57.0000 132.7000 ;
	    RECT 59.8000 130.8000 60.2000 133.1000 ;
	    RECT 63.8000 130.8000 64.2000 133.1000 ;
	    RECT 64.6000 130.8000 65.0000 132.1000 ;
	    RECT 66.2000 130.8000 66.6000 132.9000 ;
	    RECT 69.4000 130.8000 69.8000 133.1000 ;
	    RECT 70.2000 130.8000 70.6000 133.1000 ;
	    RECT 72.6000 130.8000 73.0000 132.1000 ;
	    RECT 74.2000 130.8000 74.6000 132.9000 ;
	    RECT 78.2000 130.8000 78.6000 134.1000 ;
	    RECT 80.6000 130.8000 81.0000 133.1000 ;
	    RECT 83.0000 130.8000 83.4000 132.7000 ;
	    RECT 84.6000 130.8000 85.0000 132.1000 ;
	    RECT 86.2000 130.8000 86.6000 132.1000 ;
	    RECT 87.8000 130.8000 88.2000 132.7000 ;
	    RECT 90.2000 130.8000 90.6000 133.1000 ;
	    RECT 91.8000 130.8000 92.2000 134.1000 ;
	    RECT 95.0000 130.8000 95.4000 134.1000 ;
	    RECT 100.6000 130.8000 101.0000 134.1000 ;
	    RECT 103.8000 130.8000 104.2000 134.1000 ;
	    RECT 104.6000 130.8000 105.0000 132.1000 ;
	    RECT 106.2000 130.8000 106.6000 132.1000 ;
	    RECT 107.8000 130.8000 108.2000 132.1000 ;
	    RECT 108.9000 130.8000 109.3000 133.1000 ;
	    RECT 111.0000 130.8000 111.4000 132.1000 ;
	    RECT 113.4000 130.8000 113.8000 132.1000 ;
	    RECT 115.5000 130.8000 115.9000 133.1000 ;
	    RECT 116.6000 130.8000 117.0000 132.1000 ;
	    RECT 118.2000 130.8000 118.6000 132.1000 ;
	    RECT 119.8000 130.8000 120.2000 132.1000 ;
	    RECT 121.4000 130.8000 121.8000 132.1000 ;
	    RECT 122.2000 130.8000 122.6000 133.1000 ;
	    RECT 124.6000 130.8000 125.0000 134.1000 ;
	    RECT 128.6000 130.8000 129.0000 132.7000 ;
	    RECT 131.0000 130.8000 131.4000 132.1000 ;
	    RECT 132.6000 130.8000 133.0000 132.1000 ;
	    RECT 134.2000 130.8000 134.6000 132.7000 ;
	    RECT 139.0000 130.8000 139.4000 132.7000 ;
	    RECT 142.2000 130.8000 142.6000 132.7000 ;
	    RECT 143.8000 130.8000 144.2000 132.1000 ;
	    RECT 145.4000 130.8000 145.8000 132.1000 ;
	    RECT 148.6000 130.8000 149.0000 134.1000 ;
	    RECT 151.0000 130.8000 151.4000 133.1000 ;
	    RECT 153.4000 130.8000 153.8000 132.7000 ;
	    RECT 156.1000 130.8000 156.5000 133.0000 ;
	    RECT 158.2000 130.8000 158.6000 134.1000 ;
	    RECT 161.4000 130.8000 161.8000 132.1000 ;
	    RECT 163.0000 130.8000 163.4000 132.1000 ;
	    RECT 165.1000 130.8000 165.5000 133.1000 ;
	    RECT 167.0000 130.8000 167.4000 132.7000 ;
	    RECT 170.2000 130.8000 170.6000 132.7000 ;
	    RECT 0.2000 130.2000 173.4000 130.8000 ;
	    RECT 0.6000 127.9000 1.0000 130.2000 ;
	    RECT 2.2000 127.9000 2.6000 130.2000 ;
	    RECT 5.4000 126.9000 5.8000 130.2000 ;
	    RECT 6.2000 127.9000 6.6000 130.2000 ;
	    RECT 7.8000 127.9000 8.2000 130.2000 ;
	    RECT 8.6000 126.9000 9.0000 130.2000 ;
	    RECT 11.8000 126.9000 12.2000 130.2000 ;
	    RECT 17.4000 126.9000 17.8000 130.2000 ;
	    RECT 20.6000 126.9000 21.0000 130.2000 ;
	    RECT 22.2000 128.1000 22.6000 130.2000 ;
	    RECT 23.8000 128.9000 24.2000 130.2000 ;
	    RECT 24.6000 128.9000 25.0000 130.2000 ;
	    RECT 26.2000 128.1000 26.6000 130.2000 ;
	    RECT 30.2000 126.9000 30.6000 130.2000 ;
	    RECT 33.4000 126.9000 33.8000 130.2000 ;
	    RECT 34.2000 126.9000 34.6000 130.2000 ;
	    RECT 39.0000 127.9000 39.4000 130.2000 ;
	    RECT 40.6000 128.9000 41.0000 130.2000 ;
	    RECT 43.0000 127.9000 43.4000 130.2000 ;
	    RECT 43.8000 128.9000 44.2000 130.2000 ;
	    RECT 45.4000 128.1000 45.8000 130.2000 ;
	    RECT 49.4000 126.9000 49.8000 130.2000 ;
	    RECT 50.2000 128.9000 50.6000 130.2000 ;
	    RECT 51.8000 128.1000 52.2000 130.2000 ;
	    RECT 55.8000 126.9000 56.2000 130.2000 ;
	    RECT 57.4000 127.9000 57.8000 130.2000 ;
	    RECT 63.0000 126.9000 63.4000 130.2000 ;
	    RECT 63.8000 128.9000 64.2000 130.2000 ;
	    RECT 65.4000 128.1000 65.8000 130.2000 ;
	    RECT 67.0000 126.9000 67.4000 130.2000 ;
	    RECT 70.2000 126.9000 70.6000 130.2000 ;
	    RECT 73.4000 127.9000 73.8000 130.2000 ;
	    RECT 76.6000 128.9000 77.0000 130.2000 ;
	    RECT 77.4000 126.9000 77.8000 130.2000 ;
	    RECT 80.6000 127.9000 81.0000 130.2000 ;
	    RECT 82.2000 127.9000 82.6000 130.2000 ;
	    RECT 84.6000 127.9000 85.0000 130.2000 ;
	    RECT 86.2000 128.0000 86.6000 130.2000 ;
	    RECT 89.0000 128.9000 89.4000 130.2000 ;
	    RECT 90.6000 128.9000 91.1000 130.2000 ;
	    RECT 93.4000 127.9000 93.8000 130.2000 ;
	    RECT 95.0000 128.9000 95.4000 130.2000 ;
	    RECT 96.6000 127.9000 97.0000 130.2000 ;
	    RECT 100.6000 127.9000 101.0000 130.2000 ;
	    RECT 101.4000 127.9000 101.8000 130.2000 ;
	    RECT 104.6000 128.0000 105.0000 130.2000 ;
	    RECT 107.4000 128.9000 107.8000 130.2000 ;
	    RECT 109.0000 128.9000 109.5000 130.2000 ;
	    RECT 111.8000 127.9000 112.2000 130.2000 ;
	    RECT 115.0000 127.9000 115.4000 130.2000 ;
	    RECT 117.4000 128.9000 117.8000 130.2000 ;
	    RECT 120.1000 128.0000 120.5000 130.2000 ;
	    RECT 123.0000 127.9000 123.4000 130.2000 ;
	    RECT 126.2000 128.3000 126.6000 130.2000 ;
	    RECT 128.1000 127.9000 128.5000 130.2000 ;
	    RECT 130.2000 128.9000 130.6000 130.2000 ;
	    RECT 131.0000 128.9000 131.4000 130.2000 ;
	    RECT 133.1000 127.9000 133.5000 130.2000 ;
	    RECT 134.2000 128.9000 134.6000 130.2000 ;
	    RECT 135.8000 128.9000 136.2000 130.2000 ;
	    RECT 137.4000 128.9000 137.8000 130.2000 ;
	    RECT 138.2000 127.9000 138.6000 130.2000 ;
	    RECT 140.8000 127.9000 141.2000 130.2000 ;
	    RECT 143.8000 127.9000 144.2000 130.2000 ;
	    RECT 146.2000 127.9000 146.6000 130.2000 ;
	    RECT 147.0000 128.9000 147.4000 130.2000 ;
	    RECT 149.1000 127.9000 149.5000 130.2000 ;
	    RECT 150.2000 127.9000 150.6000 130.2000 ;
	    RECT 152.8000 127.9000 153.2000 130.2000 ;
	    RECT 155.8000 127.9000 156.2000 130.2000 ;
	    RECT 158.2000 127.9000 158.6000 130.2000 ;
	    RECT 160.6000 127.9000 161.0000 130.2000 ;
	    RECT 163.0000 127.9000 163.4000 130.2000 ;
	    RECT 164.6000 127.9000 165.0000 130.2000 ;
	    RECT 167.3000 128.9000 167.8000 130.2000 ;
	    RECT 169.0000 128.9000 169.4000 130.2000 ;
	    RECT 171.8000 128.0000 172.2000 130.2000 ;
	    RECT 0.6000 110.8000 1.0000 112.1000 ;
	    RECT 2.2000 110.8000 2.6000 112.9000 ;
	    RECT 3.8000 110.8000 4.2000 113.1000 ;
	    RECT 7.0000 110.8000 7.4000 112.1000 ;
	    RECT 7.8000 110.8000 8.2000 112.1000 ;
	    RECT 11.0000 110.8000 11.4000 113.1000 ;
	    RECT 14.2000 110.8000 14.6000 114.1000 ;
	    RECT 15.8000 110.8000 16.2000 112.9000 ;
	    RECT 17.4000 110.8000 17.8000 112.1000 ;
	    RECT 19.0000 110.8000 19.4000 113.1000 ;
	    RECT 20.6000 110.8000 21.0000 112.1000 ;
	    RECT 23.8000 110.8000 24.2000 113.1000 ;
	    RECT 24.6000 110.8000 25.0000 112.1000 ;
	    RECT 26.2000 110.8000 26.6000 112.9000 ;
	    RECT 27.8000 110.8000 28.2000 114.1000 ;
	    RECT 31.0000 110.8000 31.4000 112.1000 ;
	    RECT 32.6000 110.8000 33.0000 112.1000 ;
	    RECT 34.2000 110.8000 34.6000 114.1000 ;
	    RECT 39.0000 110.8000 39.4000 113.1000 ;
	    RECT 40.6000 110.8000 41.0000 113.1000 ;
	    RECT 42.2000 110.8000 42.6000 112.1000 ;
	    RECT 43.8000 110.8000 44.2000 112.9000 ;
	    RECT 47.8000 110.8000 48.2000 114.1000 ;
	    RECT 48.6000 110.8000 49.0000 112.1000 ;
	    RECT 50.2000 110.8000 50.6000 112.9000 ;
	    RECT 51.8000 110.8000 52.2000 113.1000 ;
	    RECT 55.0000 110.8000 55.4000 112.1000 ;
	    RECT 55.8000 110.8000 56.2000 114.1000 ;
	    RECT 59.8000 110.8000 60.2000 113.1000 ;
	    RECT 63.8000 110.8000 64.2000 113.1000 ;
	    RECT 67.8000 110.8000 68.2000 114.1000 ;
	    RECT 71.0000 110.8000 71.4000 114.1000 ;
	    RECT 72.6000 110.8000 73.0000 113.0000 ;
	    RECT 75.4000 110.8000 75.8000 112.1000 ;
	    RECT 77.0000 110.8000 77.5000 112.1000 ;
	    RECT 79.8000 110.8000 80.2000 113.1000 ;
	    RECT 82.2000 110.8000 82.6000 113.1000 ;
	    RECT 84.9000 110.8000 85.4000 112.1000 ;
	    RECT 86.6000 110.8000 87.0000 112.1000 ;
	    RECT 89.4000 110.8000 89.8000 113.0000 ;
	    RECT 91.8000 110.8000 92.2000 113.0000 ;
	    RECT 94.6000 110.8000 95.0000 112.1000 ;
	    RECT 96.2000 110.8000 96.7000 112.1000 ;
	    RECT 99.0000 110.8000 99.4000 113.1000 ;
	    RECT 101.4000 110.8000 101.8000 113.0000 ;
	    RECT 104.2000 110.8000 104.6000 112.1000 ;
	    RECT 105.8000 110.8000 106.3000 112.1000 ;
	    RECT 108.6000 110.8000 109.0000 113.1000 ;
	    RECT 112.6000 110.8000 113.0000 113.1000 ;
	    RECT 115.3000 110.8000 115.8000 112.1000 ;
	    RECT 117.0000 110.8000 117.4000 112.1000 ;
	    RECT 119.8000 110.8000 120.2000 113.0000 ;
	    RECT 123.0000 110.8000 123.4000 112.7000 ;
	    RECT 124.6000 110.8000 125.0000 112.1000 ;
	    RECT 126.2000 110.8000 126.6000 112.1000 ;
	    RECT 128.3000 110.8000 128.7000 113.0000 ;
	    RECT 130.2000 110.8000 130.6000 112.1000 ;
	    RECT 131.8000 110.8000 132.2000 112.1000 ;
	    RECT 133.4000 110.8000 133.8000 112.7000 ;
	    RECT 137.4000 110.8000 137.8000 113.1000 ;
	    RECT 139.0000 110.8000 139.4000 112.7000 ;
	    RECT 142.7000 110.8000 143.1000 113.0000 ;
	    RECT 145.4000 110.8000 145.8000 112.7000 ;
	    RECT 149.4000 110.8000 149.8000 112.7000 ;
	    RECT 152.6000 110.8000 153.0000 113.1000 ;
	    RECT 154.2000 110.8000 154.6000 113.1000 ;
	    RECT 155.0000 110.8000 155.4000 113.1000 ;
	    RECT 157.4000 110.8000 157.8000 113.1000 ;
	    RECT 159.8000 110.8000 160.2000 112.7000 ;
	    RECT 163.8000 110.8000 164.2000 113.1000 ;
	    RECT 166.5000 110.8000 167.0000 112.1000 ;
	    RECT 168.2000 110.8000 168.6000 112.1000 ;
	    RECT 171.0000 110.8000 171.4000 113.0000 ;
	    RECT 0.2000 110.2000 173.4000 110.8000 ;
	    RECT 0.6000 108.9000 1.0000 110.2000 ;
	    RECT 2.2000 106.9000 2.6000 110.2000 ;
	    RECT 7.0000 107.9000 7.4000 110.2000 ;
	    RECT 10.2000 106.9000 10.6000 110.2000 ;
	    RECT 11.8000 108.1000 12.2000 110.2000 ;
	    RECT 13.4000 108.9000 13.8000 110.2000 ;
	    RECT 16.6000 106.9000 17.0000 110.2000 ;
	    RECT 18.2000 107.9000 18.6000 110.2000 ;
	    RECT 19.8000 108.9000 20.2000 110.2000 ;
	    RECT 21.4000 108.1000 21.8000 110.2000 ;
	    RECT 25.4000 106.9000 25.8000 110.2000 ;
	    RECT 27.0000 107.9000 27.4000 110.2000 ;
	    RECT 27.8000 106.9000 28.2000 110.2000 ;
	    RECT 31.0000 107.9000 31.4000 110.2000 ;
	    RECT 34.2000 108.9000 34.6000 110.2000 ;
	    RECT 37.4000 106.9000 37.8000 110.2000 ;
	    RECT 40.6000 106.9000 41.0000 110.2000 ;
	    RECT 41.4000 108.9000 41.8000 110.2000 ;
	    RECT 43.0000 108.1000 43.4000 110.2000 ;
	    RECT 45.4000 108.9000 45.8000 110.2000 ;
	    RECT 47.8000 107.9000 48.2000 110.2000 ;
	    RECT 51.0000 106.9000 51.4000 110.2000 ;
	    RECT 51.8000 108.9000 52.2000 110.2000 ;
	    RECT 53.4000 108.1000 53.8000 110.2000 ;
	    RECT 55.0000 106.9000 55.4000 110.2000 ;
	    RECT 58.2000 107.9000 58.6000 110.2000 ;
	    RECT 64.6000 106.9000 65.0000 110.2000 ;
	    RECT 67.8000 106.9000 68.2000 110.2000 ;
	    RECT 71.0000 106.9000 71.4000 110.2000 ;
	    RECT 71.8000 107.9000 72.2000 110.2000 ;
	    RECT 73.4000 107.9000 73.8000 110.2000 ;
	    RECT 74.2000 107.9000 74.6000 110.2000 ;
	    RECT 76.6000 107.9000 77.0000 110.2000 ;
	    RECT 79.8000 106.9000 80.2000 110.2000 ;
	    RECT 83.0000 106.9000 83.4000 110.2000 ;
	    RECT 83.8000 106.9000 84.2000 110.2000 ;
	    RECT 87.0000 106.9000 87.4000 110.2000 ;
	    RECT 92.6000 106.9000 93.0000 110.2000 ;
	    RECT 94.2000 107.9000 94.6000 110.2000 ;
	    RECT 96.9000 108.9000 97.4000 110.2000 ;
	    RECT 98.6000 108.9000 99.0000 110.2000 ;
	    RECT 101.4000 108.0000 101.8000 110.2000 ;
	    RECT 104.1000 108.0000 104.5000 110.2000 ;
	    RECT 107.5000 108.0000 107.9000 110.2000 ;
	    RECT 111.8000 108.0000 112.2000 110.2000 ;
	    RECT 114.6000 108.9000 115.0000 110.2000 ;
	    RECT 116.2000 108.9000 116.7000 110.2000 ;
	    RECT 119.0000 107.9000 119.4000 110.2000 ;
	    RECT 121.7000 108.0000 122.1000 110.2000 ;
	    RECT 125.1000 108.0000 125.5000 110.2000 ;
	    RECT 129.4000 108.3000 129.8000 110.2000 ;
	    RECT 131.0000 108.9000 131.4000 110.2000 ;
	    RECT 132.6000 107.9000 133.0000 110.2000 ;
	    RECT 135.6000 107.9000 136.0000 110.2000 ;
	    RECT 138.2000 107.9000 138.6000 110.2000 ;
	    RECT 139.0000 107.9000 139.4000 110.2000 ;
	    RECT 142.2000 108.9000 142.6000 110.2000 ;
	    RECT 143.8000 107.9000 144.2000 110.2000 ;
	    RECT 146.5000 108.9000 147.0000 110.2000 ;
	    RECT 148.2000 108.9000 148.6000 110.2000 ;
	    RECT 151.0000 108.0000 151.4000 110.2000 ;
	    RECT 153.4000 108.0000 153.8000 110.2000 ;
	    RECT 156.2000 108.9000 156.6000 110.2000 ;
	    RECT 157.8000 108.9000 158.3000 110.2000 ;
	    RECT 160.6000 107.9000 161.0000 110.2000 ;
	    RECT 163.0000 107.9000 163.4000 110.2000 ;
	    RECT 165.7000 108.9000 166.2000 110.2000 ;
	    RECT 167.4000 108.9000 167.8000 110.2000 ;
	    RECT 170.2000 108.0000 170.6000 110.2000 ;
	    RECT 1.4000 90.8000 1.8000 93.1000 ;
	    RECT 3.0000 90.8000 3.4000 92.1000 ;
	    RECT 6.2000 90.8000 6.6000 93.1000 ;
	    RECT 7.0000 90.8000 7.4000 92.1000 ;
	    RECT 8.6000 90.8000 9.0000 92.9000 ;
	    RECT 12.6000 90.8000 13.0000 94.1000 ;
	    RECT 13.4000 90.8000 13.8000 92.1000 ;
	    RECT 15.0000 90.8000 15.4000 92.9000 ;
	    RECT 16.6000 90.8000 17.0000 93.1000 ;
	    RECT 19.0000 90.8000 19.4000 92.1000 ;
	    RECT 23.0000 90.8000 23.4000 94.1000 ;
	    RECT 24.6000 90.8000 25.0000 93.1000 ;
	    RECT 26.2000 90.8000 26.6000 94.1000 ;
	    RECT 29.4000 90.8000 29.8000 94.1000 ;
	    RECT 33.4000 90.8000 33.8000 92.9000 ;
	    RECT 35.0000 90.8000 35.4000 92.1000 ;
	    RECT 38.2000 90.8000 38.6000 94.1000 ;
	    RECT 39.0000 90.8000 39.4000 92.1000 ;
	    RECT 42.2000 90.8000 42.6000 93.1000 ;
	    RECT 43.0000 90.8000 43.4000 92.1000 ;
	    RECT 44.6000 90.8000 45.0000 92.9000 ;
	    RECT 48.6000 90.8000 49.0000 94.1000 ;
	    RECT 49.4000 90.8000 49.8000 92.1000 ;
	    RECT 52.6000 90.8000 53.0000 93.1000 ;
	    RECT 53.4000 90.8000 53.8000 92.1000 ;
	    RECT 55.0000 90.8000 55.4000 92.9000 ;
	    RECT 56.6000 90.8000 57.0000 94.1000 ;
	    RECT 62.2000 90.8000 62.6000 92.1000 ;
	    RECT 63.0000 90.8000 63.4000 92.1000 ;
	    RECT 66.2000 90.8000 66.6000 93.1000 ;
	    RECT 67.0000 90.8000 67.4000 92.1000 ;
	    RECT 68.6000 90.8000 69.0000 92.9000 ;
	    RECT 72.6000 90.8000 73.0000 94.1000 ;
	    RECT 75.8000 90.8000 76.2000 94.1000 ;
	    RECT 76.6000 90.8000 77.0000 92.1000 ;
	    RECT 78.2000 90.8000 78.6000 92.9000 ;
	    RECT 79.8000 90.8000 80.2000 92.1000 ;
	    RECT 81.4000 90.8000 81.8000 94.1000 ;
	    RECT 86.2000 90.8000 86.6000 93.1000 ;
	    RECT 87.0000 90.8000 87.4000 94.1000 ;
	    RECT 90.2000 90.8000 90.6000 94.1000 ;
	    RECT 93.4000 90.8000 93.8000 92.1000 ;
	    RECT 95.0000 90.8000 95.4000 92.9000 ;
	    RECT 99.0000 90.8000 99.4000 94.1000 ;
	    RECT 100.1000 90.8000 100.5000 93.1000 ;
	    RECT 102.2000 90.8000 102.6000 92.1000 ;
	    RECT 103.0000 90.8000 103.4000 92.1000 ;
	    RECT 105.1000 90.8000 105.5000 93.1000 ;
	    RECT 106.5000 90.8000 106.9000 93.1000 ;
	    RECT 108.6000 90.8000 109.0000 92.1000 ;
	    RECT 109.7000 90.8000 110.1000 93.1000 ;
	    RECT 111.8000 90.8000 112.2000 92.1000 ;
	    RECT 114.5000 90.8000 114.9000 93.1000 ;
	    RECT 116.6000 90.8000 117.0000 92.1000 ;
	    RECT 118.2000 90.8000 118.6000 93.1000 ;
	    RECT 120.9000 90.8000 121.4000 92.1000 ;
	    RECT 122.6000 90.8000 123.0000 92.1000 ;
	    RECT 125.4000 90.8000 125.8000 93.0000 ;
	    RECT 127.8000 90.8000 128.2000 93.0000 ;
	    RECT 130.6000 90.8000 131.0000 92.1000 ;
	    RECT 132.2000 90.8000 132.7000 92.1000 ;
	    RECT 135.0000 90.8000 135.4000 93.1000 ;
	    RECT 138.2000 90.8000 138.6000 93.1000 ;
	    RECT 139.8000 90.8000 140.2000 92.1000 ;
	    RECT 141.4000 90.8000 141.8000 93.1000 ;
	    RECT 143.8000 90.8000 144.2000 93.0000 ;
	    RECT 146.6000 90.8000 147.0000 92.1000 ;
	    RECT 148.2000 90.8000 148.7000 92.1000 ;
	    RECT 151.0000 90.8000 151.4000 93.1000 ;
	    RECT 152.6000 90.8000 153.0000 93.1000 ;
	    RECT 154.2000 90.8000 154.6000 93.1000 ;
	    RECT 155.8000 90.8000 156.2000 93.1000 ;
	    RECT 157.4000 90.8000 157.8000 93.1000 ;
	    RECT 159.0000 90.8000 159.4000 93.1000 ;
	    RECT 160.6000 90.8000 161.0000 93.1000 ;
	    RECT 163.3000 90.8000 163.8000 92.1000 ;
	    RECT 165.0000 90.8000 165.4000 92.1000 ;
	    RECT 167.8000 90.8000 168.2000 93.0000 ;
	    RECT 170.5000 90.8000 170.9000 93.0000 ;
	    RECT 0.2000 90.2000 173.4000 90.8000 ;
	    RECT 0.6000 88.9000 1.0000 90.2000 ;
	    RECT 2.2000 87.9000 2.6000 90.2000 ;
	    RECT 5.4000 88.9000 5.8000 90.2000 ;
	    RECT 6.2000 88.9000 6.6000 90.2000 ;
	    RECT 7.8000 88.1000 8.2000 90.2000 ;
	    RECT 11.8000 86.9000 12.2000 90.2000 ;
	    RECT 15.0000 86.9000 15.4000 90.2000 ;
	    RECT 15.8000 88.9000 16.2000 90.2000 ;
	    RECT 17.4000 87.9000 17.8000 90.2000 ;
	    RECT 19.8000 88.9000 20.2000 90.2000 ;
	    RECT 21.4000 88.1000 21.8000 90.2000 ;
	    RECT 23.0000 86.9000 23.4000 90.2000 ;
	    RECT 26.2000 86.9000 26.6000 90.2000 ;
	    RECT 31.8000 86.9000 32.2000 90.2000 ;
	    RECT 34.2000 87.9000 34.6000 90.2000 ;
	    RECT 35.8000 88.1000 36.2000 90.2000 ;
	    RECT 37.4000 88.9000 37.8000 90.2000 ;
	    RECT 38.2000 87.9000 38.6000 90.2000 ;
	    RECT 40.6000 86.9000 41.0000 90.2000 ;
	    RECT 43.8000 86.9000 44.2000 90.2000 ;
	    RECT 47.0000 88.9000 47.4000 90.2000 ;
	    RECT 48.6000 87.9000 49.0000 90.2000 ;
	    RECT 51.0000 88.9000 51.4000 90.2000 ;
	    RECT 52.6000 88.1000 53.0000 90.2000 ;
	    RECT 56.6000 86.9000 57.0000 90.2000 ;
	    RECT 57.4000 88.9000 57.8000 90.2000 ;
	    RECT 59.0000 88.1000 59.4000 90.2000 ;
	    RECT 62.2000 88.9000 62.6000 90.2000 ;
	    RECT 64.6000 87.9000 65.0000 90.2000 ;
	    RECT 66.2000 87.9000 66.6000 90.2000 ;
	    RECT 70.2000 87.9000 70.6000 90.2000 ;
	    RECT 73.4000 86.9000 73.8000 90.2000 ;
	    RECT 76.6000 86.9000 77.0000 90.2000 ;
	    RECT 79.8000 86.9000 80.2000 90.2000 ;
	    RECT 80.6000 86.9000 81.0000 90.2000 ;
	    RECT 83.8000 88.9000 84.2000 90.2000 ;
	    RECT 85.4000 88.1000 85.8000 90.2000 ;
	    RECT 87.0000 87.9000 87.4000 90.2000 ;
	    RECT 91.0000 87.9000 91.4000 90.2000 ;
	    RECT 94.2000 86.9000 94.6000 90.2000 ;
	    RECT 97.4000 86.9000 97.8000 90.2000 ;
	    RECT 100.6000 86.9000 101.0000 90.2000 ;
	    RECT 102.2000 87.9000 102.6000 90.2000 ;
	    RECT 104.9000 88.9000 105.4000 90.2000 ;
	    RECT 106.6000 88.9000 107.0000 90.2000 ;
	    RECT 109.4000 88.0000 109.8000 90.2000 ;
	    RECT 113.4000 87.9000 113.8000 90.2000 ;
	    RECT 115.0000 87.9000 115.4000 90.2000 ;
	    RECT 117.7000 88.0000 118.1000 90.2000 ;
	    RECT 120.6000 88.0000 121.0000 90.2000 ;
	    RECT 123.4000 88.9000 123.8000 90.2000 ;
	    RECT 125.0000 88.9000 125.5000 90.2000 ;
	    RECT 127.8000 87.9000 128.2000 90.2000 ;
	    RECT 130.7000 88.0000 131.1000 90.2000 ;
	    RECT 133.4000 87.9000 133.8000 90.2000 ;
	    RECT 136.1000 88.9000 136.6000 90.2000 ;
	    RECT 137.8000 88.9000 138.2000 90.2000 ;
	    RECT 140.6000 88.0000 141.0000 90.2000 ;
	    RECT 142.2000 88.9000 142.6000 90.2000 ;
	    RECT 144.3000 87.9000 144.7000 90.2000 ;
	    RECT 145.4000 87.9000 145.8000 90.2000 ;
	    RECT 147.0000 87.9000 147.4000 90.2000 ;
	    RECT 148.6000 87.9000 149.0000 90.2000 ;
	    RECT 150.2000 87.9000 150.6000 90.2000 ;
	    RECT 151.8000 87.9000 152.2000 90.2000 ;
	    RECT 153.4000 88.0000 153.8000 90.2000 ;
	    RECT 156.2000 88.9000 156.6000 90.2000 ;
	    RECT 157.8000 88.9000 158.3000 90.2000 ;
	    RECT 160.6000 87.9000 161.0000 90.2000 ;
	    RECT 163.5000 88.0000 163.9000 90.2000 ;
	    RECT 166.5000 88.0000 166.9000 90.2000 ;
	    RECT 169.4000 87.9000 169.8000 90.2000 ;
	    RECT 172.6000 87.9000 173.0000 90.2000 ;
	    RECT 2.2000 70.8000 2.6000 73.1000 ;
	    RECT 3.8000 70.8000 4.2000 72.9000 ;
	    RECT 5.4000 70.8000 5.8000 72.1000 ;
	    RECT 7.0000 70.8000 7.4000 73.1000 ;
	    RECT 9.4000 70.8000 9.8000 73.1000 ;
	    RECT 11.8000 70.8000 12.2000 72.1000 ;
	    RECT 14.2000 70.8000 14.6000 73.1000 ;
	    RECT 15.0000 70.8000 15.4000 72.1000 ;
	    RECT 16.6000 70.8000 17.0000 72.9000 ;
	    RECT 18.2000 70.8000 18.6000 73.1000 ;
	    RECT 21.4000 70.8000 21.8000 72.1000 ;
	    RECT 22.2000 70.8000 22.6000 73.1000 ;
	    RECT 25.4000 70.8000 25.8000 72.1000 ;
	    RECT 26.2000 70.8000 26.6000 72.1000 ;
	    RECT 29.4000 70.8000 29.8000 73.1000 ;
	    RECT 31.0000 70.8000 31.4000 72.9000 ;
	    RECT 32.6000 70.8000 33.0000 72.1000 ;
	    RECT 34.2000 70.8000 34.6000 72.1000 ;
	    RECT 35.8000 70.8000 36.2000 72.1000 ;
	    RECT 37.4000 70.8000 37.8000 72.7000 ;
	    RECT 40.6000 70.8000 41.0000 73.1000 ;
	    RECT 41.4000 70.8000 41.8000 72.1000 ;
	    RECT 44.6000 70.8000 45.0000 73.1000 ;
	    RECT 45.4000 70.8000 45.8000 72.1000 ;
	    RECT 47.0000 70.8000 47.4000 72.9000 ;
	    RECT 51.0000 70.8000 51.4000 74.1000 ;
	    RECT 51.8000 70.8000 52.2000 72.1000 ;
	    RECT 53.4000 70.8000 53.8000 72.9000 ;
	    RECT 55.8000 70.8000 56.2000 73.1000 ;
	    RECT 59.8000 70.8000 60.2000 74.1000 ;
	    RECT 64.6000 70.8000 65.0000 74.1000 ;
	    RECT 66.2000 70.8000 66.6000 73.1000 ;
	    RECT 70.2000 70.8000 70.6000 74.1000 ;
	    RECT 73.4000 70.8000 73.8000 74.1000 ;
	    RECT 75.0000 70.8000 75.4000 72.9000 ;
	    RECT 76.6000 70.8000 77.0000 72.1000 ;
	    RECT 77.4000 70.8000 77.8000 72.1000 ;
	    RECT 79.0000 70.8000 79.4000 72.9000 ;
	    RECT 80.6000 70.8000 81.0000 74.1000 ;
	    RECT 83.8000 70.8000 84.2000 72.1000 ;
	    RECT 85.4000 70.8000 85.8000 72.1000 ;
	    RECT 88.1000 70.8000 88.5000 73.0000 ;
	    RECT 91.5000 70.8000 91.9000 73.0000 ;
	    RECT 95.8000 70.8000 96.2000 74.1000 ;
	    RECT 96.9000 70.8000 97.3000 73.1000 ;
	    RECT 99.0000 70.8000 99.4000 72.1000 ;
	    RECT 100.1000 70.8000 100.5000 73.1000 ;
	    RECT 102.2000 70.8000 102.6000 72.1000 ;
	    RECT 103.0000 70.8000 103.4000 73.1000 ;
	    RECT 104.6000 70.8000 105.0000 73.1000 ;
	    RECT 106.2000 70.8000 106.6000 73.1000 ;
	    RECT 107.8000 70.8000 108.2000 73.1000 ;
	    RECT 109.4000 70.8000 109.8000 73.1000 ;
	    RECT 111.0000 70.8000 111.4000 73.1000 ;
	    RECT 115.0000 70.8000 115.4000 73.1000 ;
	    RECT 117.7000 70.8000 118.2000 72.1000 ;
	    RECT 119.4000 70.8000 119.8000 72.1000 ;
	    RECT 122.2000 70.8000 122.6000 73.0000 ;
	    RECT 125.1000 70.8000 125.5000 73.0000 ;
	    RECT 127.8000 70.8000 128.2000 73.1000 ;
	    RECT 130.5000 70.8000 131.0000 72.1000 ;
	    RECT 132.2000 70.8000 132.6000 72.1000 ;
	    RECT 135.0000 70.8000 135.4000 73.0000 ;
	    RECT 136.9000 70.8000 137.3000 73.1000 ;
	    RECT 139.0000 70.8000 139.4000 72.1000 ;
	    RECT 140.6000 70.8000 141.0000 73.1000 ;
	    RECT 142.2000 70.8000 142.6000 73.1000 ;
	    RECT 144.1000 70.8000 144.5000 73.1000 ;
	    RECT 146.2000 70.8000 146.6000 72.1000 ;
	    RECT 147.3000 70.8000 147.7000 73.1000 ;
	    RECT 149.4000 70.8000 149.8000 72.1000 ;
	    RECT 150.2000 70.8000 150.6000 72.1000 ;
	    RECT 152.3000 70.8000 152.7000 73.1000 ;
	    RECT 154.2000 70.8000 154.6000 73.1000 ;
	    RECT 156.9000 70.8000 157.4000 72.1000 ;
	    RECT 158.6000 70.8000 159.0000 72.1000 ;
	    RECT 161.4000 70.8000 161.8000 73.0000 ;
	    RECT 163.8000 70.8000 164.2000 73.1000 ;
	    RECT 166.5000 70.8000 167.0000 72.1000 ;
	    RECT 168.2000 70.8000 168.6000 72.1000 ;
	    RECT 171.0000 70.8000 171.4000 73.0000 ;
	    RECT 0.2000 70.2000 173.4000 70.8000 ;
	    RECT 3.0000 66.9000 3.4000 70.2000 ;
	    RECT 3.8000 67.9000 4.2000 70.2000 ;
	    RECT 5.4000 68.9000 5.8000 70.2000 ;
	    RECT 7.0000 68.1000 7.4000 70.2000 ;
	    RECT 8.6000 66.9000 9.0000 70.2000 ;
	    RECT 11.8000 66.9000 12.2000 70.2000 ;
	    RECT 17.4000 66.9000 17.8000 70.2000 ;
	    RECT 18.2000 66.9000 18.6000 70.2000 ;
	    RECT 23.0000 67.9000 23.4000 70.2000 ;
	    RECT 26.2000 66.9000 26.6000 70.2000 ;
	    RECT 27.0000 68.9000 27.4000 70.2000 ;
	    RECT 28.6000 68.1000 29.0000 70.2000 ;
	    RECT 30.2000 66.9000 30.6000 70.2000 ;
	    RECT 33.4000 67.9000 33.8000 70.2000 ;
	    RECT 36.6000 68.9000 37.0000 70.2000 ;
	    RECT 37.4000 67.9000 37.8000 70.2000 ;
	    RECT 41.4000 67.9000 41.8000 70.2000 ;
	    RECT 42.2000 68.9000 42.6000 70.2000 ;
	    RECT 44.6000 68.3000 45.0000 70.2000 ;
	    RECT 48.6000 67.9000 49.0000 70.2000 ;
	    RECT 49.4000 68.9000 49.8000 70.2000 ;
	    RECT 52.6000 68.3000 53.0000 70.2000 ;
	    RECT 54.2000 68.9000 54.6000 70.2000 ;
	    RECT 55.8000 67.9000 56.2000 70.2000 ;
	    RECT 59.8000 67.9000 60.2000 70.2000 ;
	    RECT 62.2000 68.9000 62.6000 70.2000 ;
	    RECT 65.4000 67.9000 65.8000 70.2000 ;
	    RECT 66.2000 67.9000 66.6000 70.2000 ;
	    RECT 69.4000 68.9000 69.8000 70.2000 ;
	    RECT 71.0000 68.1000 71.4000 70.2000 ;
	    RECT 72.6000 68.9000 73.0000 70.2000 ;
	    RECT 73.4000 68.9000 73.8000 70.2000 ;
	    RECT 76.6000 67.9000 77.0000 70.2000 ;
	    RECT 78.7000 68.0000 79.1000 70.2000 ;
	    RECT 81.9000 68.0000 82.3000 70.2000 ;
	    RECT 84.6000 67.9000 85.0000 70.2000 ;
	    RECT 87.3000 68.9000 87.8000 70.2000 ;
	    RECT 89.0000 68.9000 89.4000 70.2000 ;
	    RECT 91.8000 68.0000 92.2000 70.2000 ;
	    RECT 93.7000 67.9000 94.1000 70.2000 ;
	    RECT 95.8000 68.9000 96.2000 70.2000 ;
	    RECT 96.6000 67.9000 97.0000 70.2000 ;
	    RECT 99.5000 68.0000 99.9000 70.2000 ;
	    RECT 102.2000 67.9000 102.6000 70.2000 ;
	    RECT 104.9000 68.9000 105.4000 70.2000 ;
	    RECT 106.6000 68.9000 107.0000 70.2000 ;
	    RECT 109.4000 68.0000 109.8000 70.2000 ;
	    RECT 112.6000 67.9000 113.0000 70.2000 ;
	    RECT 114.2000 67.9000 114.6000 70.2000 ;
	    RECT 115.8000 67.9000 116.2000 70.2000 ;
	    RECT 117.4000 67.9000 117.8000 70.2000 ;
	    RECT 119.0000 67.9000 119.4000 70.2000 ;
	    RECT 120.6000 67.9000 121.0000 70.2000 ;
	    RECT 123.3000 68.9000 123.8000 70.2000 ;
	    RECT 125.0000 68.9000 125.4000 70.2000 ;
	    RECT 127.8000 68.0000 128.2000 70.2000 ;
	    RECT 130.5000 68.0000 130.9000 70.2000 ;
	    RECT 133.4000 67.9000 133.8000 70.2000 ;
	    RECT 136.1000 68.9000 136.6000 70.2000 ;
	    RECT 137.8000 68.9000 138.2000 70.2000 ;
	    RECT 140.6000 68.0000 141.0000 70.2000 ;
	    RECT 143.5000 68.0000 143.9000 70.2000 ;
	    RECT 146.2000 68.0000 146.6000 70.2000 ;
	    RECT 149.0000 68.9000 149.4000 70.2000 ;
	    RECT 150.6000 68.9000 151.1000 70.2000 ;
	    RECT 153.4000 67.9000 153.8000 70.2000 ;
	    RECT 156.3000 68.0000 156.7000 70.2000 ;
	    RECT 159.0000 67.9000 159.4000 70.2000 ;
	    RECT 161.7000 68.9000 162.2000 70.2000 ;
	    RECT 163.4000 68.9000 163.8000 70.2000 ;
	    RECT 166.2000 68.0000 166.6000 70.2000 ;
	    RECT 168.6000 67.9000 169.0000 70.2000 ;
	    RECT 171.0000 67.9000 171.4000 70.2000 ;
	    RECT 3.0000 50.8000 3.4000 54.1000 ;
	    RECT 6.2000 50.8000 6.6000 54.1000 ;
	    RECT 7.0000 50.8000 7.4000 53.1000 ;
	    RECT 9.4000 50.8000 9.8000 52.1000 ;
	    RECT 11.0000 50.8000 11.4000 52.7000 ;
	    RECT 15.8000 50.8000 16.2000 54.1000 ;
	    RECT 19.0000 50.8000 19.4000 54.1000 ;
	    RECT 19.8000 50.8000 20.2000 54.1000 ;
	    RECT 23.0000 50.8000 23.4000 54.1000 ;
	    RECT 26.2000 50.8000 26.6000 54.1000 ;
	    RECT 30.2000 50.8000 30.6000 52.9000 ;
	    RECT 31.8000 50.8000 32.2000 52.1000 ;
	    RECT 32.9000 50.8000 33.3000 53.1000 ;
	    RECT 35.0000 50.8000 35.4000 52.1000 ;
	    RECT 36.1000 50.8000 36.5000 53.1000 ;
	    RECT 38.2000 50.8000 38.6000 52.1000 ;
	    RECT 39.3000 50.8000 39.7000 53.1000 ;
	    RECT 41.4000 50.8000 41.8000 52.1000 ;
	    RECT 42.5000 50.8000 42.9000 53.1000 ;
	    RECT 44.6000 50.8000 45.0000 52.1000 ;
	    RECT 46.2000 50.8000 46.6000 53.1000 ;
	    RECT 47.8000 50.8000 48.2000 53.1000 ;
	    RECT 50.5000 50.8000 51.0000 52.1000 ;
	    RECT 52.2000 50.8000 52.6000 52.1000 ;
	    RECT 55.0000 50.8000 55.4000 53.0000 ;
	    RECT 59.0000 50.8000 59.4000 54.1000 ;
	    RECT 62.2000 50.8000 62.6000 53.1000 ;
	    RECT 64.9000 50.8000 65.4000 52.1000 ;
	    RECT 66.6000 50.8000 67.0000 52.1000 ;
	    RECT 69.4000 50.8000 69.8000 53.0000 ;
	    RECT 73.4000 50.8000 73.8000 54.1000 ;
	    RECT 76.6000 50.8000 77.0000 54.1000 ;
	    RECT 77.4000 50.8000 77.8000 54.1000 ;
	    RECT 81.4000 50.8000 81.8000 53.1000 ;
	    RECT 84.1000 50.8000 84.6000 52.1000 ;
	    RECT 85.8000 50.8000 86.2000 52.1000 ;
	    RECT 88.6000 50.8000 89.0000 53.0000 ;
	    RECT 91.0000 50.8000 91.4000 53.1000 ;
	    RECT 93.7000 50.8000 94.2000 52.1000 ;
	    RECT 95.4000 50.8000 95.8000 52.1000 ;
	    RECT 98.2000 50.8000 98.6000 53.0000 ;
	    RECT 100.6000 50.8000 101.0000 53.1000 ;
	    RECT 101.4000 50.8000 101.8000 53.1000 ;
	    RECT 103.0000 50.8000 103.4000 53.1000 ;
	    RECT 104.6000 50.8000 105.0000 53.1000 ;
	    RECT 106.2000 50.8000 106.6000 53.1000 ;
	    RECT 107.8000 50.8000 108.2000 53.1000 ;
	    RECT 111.0000 50.8000 111.4000 54.1000 ;
	    RECT 114.2000 50.8000 114.6000 53.1000 ;
	    RECT 115.8000 50.8000 116.2000 54.1000 ;
	    RECT 119.0000 50.8000 119.4000 52.1000 ;
	    RECT 122.2000 50.8000 122.6000 53.1000 ;
	    RECT 123.8000 50.8000 124.2000 53.1000 ;
	    RECT 125.4000 50.8000 125.8000 53.1000 ;
	    RECT 128.6000 50.8000 129.0000 52.1000 ;
	    RECT 129.4000 50.8000 129.8000 53.1000 ;
	    RECT 132.6000 50.8000 133.0000 52.1000 ;
	    RECT 134.2000 50.8000 134.6000 53.1000 ;
	    RECT 135.0000 50.8000 135.4000 54.1000 ;
	    RECT 138.2000 50.8000 138.6000 52.1000 ;
	    RECT 139.8000 50.8000 140.2000 52.9000 ;
	    RECT 141.4000 50.8000 141.8000 54.1000 ;
	    RECT 144.6000 50.8000 145.0000 54.1000 ;
	    RECT 147.8000 50.8000 148.2000 53.1000 ;
	    RECT 151.0000 50.8000 151.4000 52.1000 ;
	    RECT 151.8000 50.8000 152.2000 53.1000 ;
	    RECT 154.2000 50.8000 154.6000 53.1000 ;
	    RECT 156.6000 50.8000 157.0000 52.1000 ;
	    RECT 158.2000 50.8000 158.6000 52.1000 ;
	    RECT 160.6000 50.8000 161.0000 52.7000 ;
	    RECT 164.3000 50.8000 164.7000 53.0000 ;
	    RECT 166.2000 50.8000 166.6000 52.1000 ;
	    RECT 169.4000 50.8000 169.8000 53.1000 ;
	    RECT 171.0000 50.8000 171.4000 53.1000 ;
	    RECT 0.2000 50.2000 173.4000 50.8000 ;
	    RECT 0.6000 46.9000 1.0000 50.2000 ;
	    RECT 4.6000 48.1000 5.0000 50.2000 ;
	    RECT 6.2000 48.9000 6.6000 50.2000 ;
	    RECT 7.8000 48.9000 8.2000 50.2000 ;
	    RECT 10.2000 47.9000 10.6000 50.2000 ;
	    RECT 11.0000 47.9000 11.4000 50.2000 ;
	    RECT 13.4000 48.9000 13.8000 50.2000 ;
	    RECT 15.0000 47.9000 15.4000 50.2000 ;
	    RECT 17.4000 46.9000 17.8000 50.2000 ;
	    RECT 21.4000 48.1000 21.8000 50.2000 ;
	    RECT 23.0000 48.9000 23.4000 50.2000 ;
	    RECT 23.8000 46.9000 24.2000 50.2000 ;
	    RECT 27.0000 47.9000 27.4000 50.2000 ;
	    RECT 29.4000 46.9000 29.8000 50.2000 ;
	    RECT 32.6000 46.9000 33.0000 50.2000 ;
	    RECT 36.6000 48.1000 37.0000 50.2000 ;
	    RECT 38.2000 48.9000 38.6000 50.2000 ;
	    RECT 39.0000 47.9000 39.4000 50.2000 ;
	    RECT 41.4000 47.9000 41.8000 50.2000 ;
	    RECT 43.8000 47.9000 44.2000 50.2000 ;
	    RECT 47.0000 48.9000 47.4000 50.2000 ;
	    RECT 48.6000 48.9000 49.0000 50.2000 ;
	    RECT 49.4000 48.9000 49.8000 50.2000 ;
	    RECT 52.6000 47.9000 53.0000 50.2000 ;
	    RECT 53.4000 48.9000 53.8000 50.2000 ;
	    RECT 55.0000 48.1000 55.4000 50.2000 ;
	    RECT 59.0000 46.9000 59.4000 50.2000 ;
	    RECT 61.4000 48.9000 61.8000 50.2000 ;
	    RECT 63.0000 48.1000 63.4000 50.2000 ;
	    RECT 67.0000 46.9000 67.4000 50.2000 ;
	    RECT 67.8000 46.9000 68.2000 50.2000 ;
	    RECT 71.0000 46.9000 71.4000 50.2000 ;
	    RECT 75.0000 48.1000 75.4000 50.2000 ;
	    RECT 76.6000 48.9000 77.0000 50.2000 ;
	    RECT 77.4000 47.9000 77.8000 50.2000 ;
	    RECT 79.8000 48.9000 80.2000 50.2000 ;
	    RECT 83.0000 47.9000 83.4000 50.2000 ;
	    RECT 83.8000 46.9000 84.2000 50.2000 ;
	    RECT 87.8000 48.1000 88.2000 50.2000 ;
	    RECT 89.4000 48.9000 89.8000 50.2000 ;
	    RECT 90.2000 47.9000 90.6000 50.2000 ;
	    RECT 93.4000 48.9000 93.8000 50.2000 ;
	    RECT 95.0000 48.9000 95.4000 50.2000 ;
	    RECT 98.2000 46.9000 98.6000 50.2000 ;
	    RECT 99.0000 46.9000 99.4000 50.2000 ;
	    RECT 103.8000 47.9000 104.2000 50.2000 ;
	    RECT 104.6000 47.9000 105.0000 50.2000 ;
	    RECT 108.6000 48.3000 109.0000 50.2000 ;
	    RECT 111.0000 48.9000 111.4000 50.2000 ;
	    RECT 113.4000 47.9000 113.8000 50.2000 ;
	    RECT 115.0000 47.9000 115.4000 50.2000 ;
	    RECT 115.8000 46.9000 116.2000 50.2000 ;
	    RECT 119.8000 48.1000 120.2000 50.2000 ;
	    RECT 121.4000 48.9000 121.8000 50.2000 ;
	    RECT 122.2000 46.9000 122.6000 50.2000 ;
	    RECT 125.4000 46.9000 125.8000 50.2000 ;
	    RECT 128.6000 46.9000 129.0000 50.2000 ;
	    RECT 132.6000 48.1000 133.0000 50.2000 ;
	    RECT 134.2000 48.9000 134.6000 50.2000 ;
	    RECT 135.0000 48.9000 135.4000 50.2000 ;
	    RECT 136.6000 48.1000 137.0000 50.2000 ;
	    RECT 138.2000 48.9000 138.6000 50.2000 ;
	    RECT 139.8000 48.1000 140.2000 50.2000 ;
	    RECT 141.4000 46.9000 141.8000 50.2000 ;
	    RECT 146.2000 47.9000 146.6000 50.2000 ;
	    RECT 147.0000 46.9000 147.4000 50.2000 ;
	    RECT 150.2000 46.9000 150.6000 50.2000 ;
	    RECT 153.4000 48.9000 153.8000 50.2000 ;
	    RECT 155.0000 48.1000 155.4000 50.2000 ;
	    RECT 159.0000 46.9000 159.4000 50.2000 ;
	    RECT 159.8000 47.9000 160.2000 50.2000 ;
	    RECT 162.2000 46.9000 162.6000 50.2000 ;
	    RECT 167.8000 46.9000 168.2000 50.2000 ;
	    RECT 169.4000 48.1000 169.8000 50.2000 ;
	    RECT 171.0000 48.9000 171.4000 50.2000 ;
	    RECT 3.0000 30.8000 3.4000 34.1000 ;
	    RECT 6.2000 30.8000 6.6000 34.1000 ;
	    RECT 7.0000 30.8000 7.4000 34.1000 ;
	    RECT 12.6000 30.8000 13.0000 34.1000 ;
	    RECT 15.8000 30.8000 16.2000 34.1000 ;
	    RECT 16.6000 30.8000 17.0000 34.1000 ;
	    RECT 19.8000 30.8000 20.2000 33.1000 ;
	    RECT 22.2000 30.8000 22.6000 34.1000 ;
	    RECT 26.2000 30.8000 26.6000 32.9000 ;
	    RECT 27.8000 30.8000 28.2000 32.1000 ;
	    RECT 28.6000 30.8000 29.0000 34.1000 ;
	    RECT 32.6000 30.8000 33.0000 32.9000 ;
	    RECT 34.2000 30.8000 34.6000 32.1000 ;
	    RECT 35.0000 30.8000 35.4000 33.1000 ;
	    RECT 38.2000 30.8000 38.6000 32.1000 ;
	    RECT 40.6000 30.8000 41.0000 32.7000 ;
	    RECT 43.0000 30.8000 43.4000 32.1000 ;
	    RECT 43.8000 30.8000 44.2000 32.1000 ;
	    RECT 45.4000 30.8000 45.8000 32.9000 ;
	    RECT 49.4000 30.8000 49.8000 34.1000 ;
	    RECT 50.2000 30.8000 50.6000 32.1000 ;
	    RECT 53.4000 30.8000 53.8000 33.1000 ;
	    RECT 56.6000 30.8000 57.0000 34.1000 ;
	    RECT 59.0000 30.8000 59.4000 33.1000 ;
	    RECT 61.4000 30.8000 61.8000 33.1000 ;
	    RECT 65.4000 30.8000 65.8000 34.1000 ;
	    RECT 68.6000 30.8000 69.0000 34.1000 ;
	    RECT 69.4000 30.8000 69.8000 34.1000 ;
	    RECT 75.0000 30.8000 75.4000 34.1000 ;
	    RECT 77.4000 30.8000 77.8000 32.7000 ;
	    RECT 79.8000 30.8000 80.2000 32.1000 ;
	    RECT 80.6000 30.8000 81.0000 33.1000 ;
	    RECT 82.2000 30.8000 82.6000 33.1000 ;
	    RECT 83.0000 30.8000 83.4000 32.1000 ;
	    RECT 86.2000 30.8000 86.6000 33.1000 ;
	    RECT 87.0000 30.8000 87.4000 32.1000 ;
	    RECT 88.6000 30.8000 89.0000 33.1000 ;
	    RECT 91.0000 30.8000 91.4000 32.1000 ;
	    RECT 92.6000 30.8000 93.0000 32.9000 ;
	    RECT 96.6000 30.8000 97.0000 34.1000 ;
	    RECT 99.8000 30.8000 100.2000 34.1000 ;
	    RECT 101.4000 30.8000 101.8000 32.9000 ;
	    RECT 103.0000 30.8000 103.4000 32.1000 ;
	    RECT 103.8000 30.8000 104.2000 32.1000 ;
	    RECT 107.8000 30.8000 108.2000 34.1000 ;
	    RECT 108.6000 30.8000 109.0000 34.1000 ;
	    RECT 113.4000 30.8000 113.8000 32.1000 ;
	    RECT 115.0000 30.8000 115.4000 32.9000 ;
	    RECT 119.0000 30.8000 119.4000 34.1000 ;
	    RECT 119.8000 30.8000 120.2000 34.1000 ;
	    RECT 123.0000 30.8000 123.4000 33.1000 ;
	    RECT 124.6000 30.8000 125.0000 34.1000 ;
	    RECT 127.8000 30.8000 128.2000 32.1000 ;
	    RECT 129.4000 30.8000 129.8000 32.1000 ;
	    RECT 131.0000 30.8000 131.4000 32.9000 ;
	    RECT 132.6000 30.8000 133.0000 32.1000 ;
	    RECT 135.8000 30.8000 136.2000 33.1000 ;
	    RECT 136.6000 30.8000 137.0000 34.1000 ;
	    RECT 141.4000 30.8000 141.8000 33.1000 ;
	    RECT 144.6000 30.8000 145.0000 34.1000 ;
	    RECT 145.4000 30.8000 145.8000 34.1000 ;
	    RECT 151.0000 30.8000 151.4000 34.1000 ;
	    RECT 152.6000 30.8000 153.0000 33.1000 ;
	    RECT 153.4000 30.8000 153.8000 34.1000 ;
	    RECT 157.4000 30.8000 157.8000 33.1000 ;
	    RECT 159.8000 30.8000 160.2000 33.1000 ;
	    RECT 161.4000 30.8000 161.8000 34.1000 ;
	    RECT 164.6000 30.8000 165.0000 34.1000 ;
	    RECT 167.8000 30.8000 168.2000 32.1000 ;
	    RECT 171.0000 30.8000 171.4000 33.1000 ;
	    RECT 0.2000 30.2000 173.4000 30.8000 ;
	    RECT 0.6000 28.9000 1.0000 30.2000 ;
	    RECT 3.8000 27.9000 4.2000 30.2000 ;
	    RECT 5.4000 28.1000 5.8000 30.2000 ;
	    RECT 7.0000 28.9000 7.4000 30.2000 ;
	    RECT 10.2000 26.9000 10.6000 30.2000 ;
	    RECT 11.8000 27.9000 12.2000 30.2000 ;
	    RECT 13.4000 26.9000 13.8000 30.2000 ;
	    RECT 16.6000 26.9000 17.0000 30.2000 ;
	    RECT 20.6000 27.9000 21.0000 30.2000 ;
	    RECT 22.2000 26.9000 22.6000 30.2000 ;
	    RECT 26.2000 28.1000 26.6000 30.2000 ;
	    RECT 27.8000 28.9000 28.2000 30.2000 ;
	    RECT 29.4000 27.9000 29.8000 30.2000 ;
	    RECT 31.0000 27.9000 31.4000 30.2000 ;
	    RECT 33.4000 26.9000 33.8000 30.2000 ;
	    RECT 37.4000 28.1000 37.8000 30.2000 ;
	    RECT 39.0000 28.9000 39.4000 30.2000 ;
	    RECT 40.6000 28.9000 41.0000 30.2000 ;
	    RECT 41.4000 28.9000 41.8000 30.2000 ;
	    RECT 44.6000 27.9000 45.0000 30.2000 ;
	    RECT 45.4000 28.9000 45.8000 30.2000 ;
	    RECT 48.6000 27.9000 49.0000 30.2000 ;
	    RECT 49.4000 28.9000 49.8000 30.2000 ;
	    RECT 51.0000 28.1000 51.4000 30.2000 ;
	    RECT 55.0000 26.9000 55.4000 30.2000 ;
	    RECT 58.2000 26.9000 58.6000 30.2000 ;
	    RECT 59.8000 27.9000 60.2000 30.2000 ;
	    RECT 64.6000 27.9000 65.0000 30.2000 ;
	    RECT 67.0000 27.9000 67.4000 30.2000 ;
	    RECT 68.6000 27.9000 69.0000 30.2000 ;
	    RECT 70.2000 28.9000 70.6000 30.2000 ;
	    RECT 71.8000 28.1000 72.2000 30.2000 ;
	    RECT 73.4000 26.9000 73.8000 30.2000 ;
	    RECT 78.2000 27.9000 78.6000 30.2000 ;
	    RECT 79.8000 27.9000 80.2000 30.2000 ;
	    RECT 81.4000 26.9000 81.8000 30.2000 ;
	    RECT 84.6000 28.9000 85.0000 30.2000 ;
	    RECT 86.2000 28.1000 86.6000 30.2000 ;
	    RECT 87.8000 28.9000 88.2000 30.2000 ;
	    RECT 89.4000 27.9000 89.8000 30.2000 ;
	    RECT 92.6000 28.9000 93.0000 30.2000 ;
	    RECT 95.8000 26.9000 96.2000 30.2000 ;
	    RECT 99.0000 26.9000 99.4000 30.2000 ;
	    RECT 99.8000 26.9000 100.2000 30.2000 ;
	    RECT 103.0000 28.9000 103.4000 30.2000 ;
	    RECT 106.2000 27.9000 106.6000 30.2000 ;
	    RECT 107.0000 26.9000 107.4000 30.2000 ;
	    RECT 111.0000 27.9000 111.4000 30.2000 ;
	    RECT 115.8000 27.9000 116.2000 30.2000 ;
	    RECT 118.2000 27.9000 118.6000 30.2000 ;
	    RECT 119.0000 28.9000 119.4000 30.2000 ;
	    RECT 120.6000 28.1000 121.0000 30.2000 ;
	    RECT 124.6000 26.9000 125.0000 30.2000 ;
	    RECT 125.4000 27.9000 125.8000 30.2000 ;
	    RECT 127.8000 28.9000 128.2000 30.2000 ;
	    RECT 129.4000 28.1000 129.8000 30.2000 ;
	    RECT 133.4000 26.9000 133.8000 30.2000 ;
	    RECT 134.2000 26.9000 134.6000 30.2000 ;
	    RECT 137.4000 27.9000 137.8000 30.2000 ;
	    RECT 139.8000 28.9000 140.2000 30.2000 ;
	    RECT 141.4000 28.1000 141.8000 30.2000 ;
	    RECT 145.4000 26.9000 145.8000 30.2000 ;
	    RECT 146.2000 27.9000 146.6000 30.2000 ;
	    RECT 147.8000 27.9000 148.2000 30.2000 ;
	    RECT 148.6000 27.9000 149.0000 30.2000 ;
	    RECT 151.0000 26.9000 151.4000 30.2000 ;
	    RECT 154.2000 27.9000 154.6000 30.2000 ;
	    RECT 157.4000 27.9000 157.8000 30.2000 ;
	    RECT 159.8000 27.9000 160.2000 30.2000 ;
	    RECT 162.5000 28.9000 163.0000 30.2000 ;
	    RECT 164.2000 28.9000 164.6000 30.2000 ;
	    RECT 167.0000 28.0000 167.4000 30.2000 ;
	    RECT 168.6000 28.9000 169.0000 30.2000 ;
	    RECT 170.2000 28.1000 170.6000 30.2000 ;
	    RECT 0.6000 10.8000 1.0000 13.1000 ;
	    RECT 2.2000 10.8000 2.6000 13.1000 ;
	    RECT 5.4000 10.8000 5.8000 14.1000 ;
	    RECT 7.0000 10.8000 7.4000 12.9000 ;
	    RECT 8.6000 10.8000 9.0000 12.1000 ;
	    RECT 11.8000 10.8000 12.2000 14.1000 ;
	    RECT 13.4000 10.8000 13.8000 13.1000 ;
	    RECT 14.2000 10.8000 14.6000 14.1000 ;
	    RECT 17.4000 10.8000 17.8000 14.1000 ;
	    RECT 20.6000 10.8000 21.0000 13.1000 ;
	    RECT 23.0000 10.8000 23.4000 14.1000 ;
	    RECT 26.2000 10.8000 26.6000 14.1000 ;
	    RECT 30.2000 10.8000 30.6000 13.1000 ;
	    RECT 31.8000 10.8000 32.2000 14.1000 ;
	    RECT 35.8000 10.8000 36.2000 12.9000 ;
	    RECT 37.4000 10.8000 37.8000 12.1000 ;
	    RECT 39.0000 10.8000 39.4000 12.9000 ;
	    RECT 40.6000 10.8000 41.0000 12.1000 ;
	    RECT 42.2000 10.8000 42.6000 12.9000 ;
	    RECT 43.8000 10.8000 44.2000 12.1000 ;
	    RECT 45.4000 10.8000 45.8000 12.7000 ;
	    RECT 48.6000 10.8000 49.0000 12.1000 ;
	    RECT 51.8000 10.8000 52.2000 14.1000 ;
	    RECT 53.4000 10.8000 53.8000 12.9000 ;
	    RECT 55.0000 10.8000 55.4000 12.1000 ;
	    RECT 57.4000 10.8000 57.8000 12.7000 ;
	    RECT 59.8000 10.8000 60.2000 12.1000 ;
	    RECT 62.2000 10.8000 62.6000 12.1000 ;
	    RECT 64.6000 10.8000 65.0000 12.7000 ;
	    RECT 69.4000 10.8000 69.8000 14.1000 ;
	    RECT 70.2000 10.8000 70.6000 12.1000 ;
	    RECT 71.8000 10.8000 72.2000 12.9000 ;
	    RECT 75.0000 10.8000 75.4000 12.7000 ;
	    RECT 77.4000 10.8000 77.8000 12.1000 ;
	    RECT 78.2000 10.8000 78.6000 12.1000 ;
	    RECT 79.8000 10.8000 80.2000 12.9000 ;
	    RECT 81.4000 10.8000 81.8000 14.1000 ;
	    RECT 84.6000 10.8000 85.0000 14.1000 ;
	    RECT 88.6000 10.8000 89.0000 12.9000 ;
	    RECT 90.2000 10.8000 90.6000 12.1000 ;
	    RECT 91.0000 10.8000 91.4000 14.1000 ;
	    RECT 95.0000 10.8000 95.4000 12.9000 ;
	    RECT 96.6000 10.8000 97.0000 12.1000 ;
	    RECT 97.4000 10.8000 97.8000 13.1000 ;
	    RECT 100.6000 10.8000 101.0000 12.1000 ;
	    RECT 103.8000 10.8000 104.2000 14.1000 ;
	    RECT 104.6000 10.8000 105.0000 12.1000 ;
	    RECT 106.2000 10.8000 106.6000 12.9000 ;
	    RECT 110.2000 10.8000 110.6000 14.1000 ;
	    RECT 115.0000 10.8000 115.4000 14.1000 ;
	    RECT 116.6000 10.8000 117.0000 12.9000 ;
	    RECT 118.2000 10.8000 118.6000 12.1000 ;
	    RECT 119.8000 10.8000 120.2000 12.9000 ;
	    RECT 121.4000 10.8000 121.8000 12.1000 ;
	    RECT 124.6000 10.8000 125.0000 14.1000 ;
	    RECT 127.8000 10.8000 128.2000 14.1000 ;
	    RECT 129.4000 10.8000 129.8000 13.1000 ;
	    RECT 131.8000 10.8000 132.2000 12.9000 ;
	    RECT 133.4000 10.8000 133.8000 12.1000 ;
	    RECT 135.0000 10.8000 135.4000 12.9000 ;
	    RECT 136.6000 10.8000 137.0000 12.1000 ;
	    RECT 137.4000 10.8000 137.8000 12.1000 ;
	    RECT 140.6000 10.8000 141.0000 12.7000 ;
	    RECT 143.8000 10.8000 144.2000 12.7000 ;
	    RECT 146.2000 10.8000 146.6000 12.1000 ;
	    RECT 149.4000 10.8000 149.8000 14.1000 ;
	    RECT 151.0000 10.8000 151.4000 12.9000 ;
	    RECT 152.6000 10.8000 153.0000 12.1000 ;
	    RECT 155.0000 10.8000 155.4000 12.7000 ;
	    RECT 156.6000 10.8000 157.0000 12.1000 ;
	    RECT 158.2000 10.8000 158.6000 14.1000 ;
	    RECT 161.4000 10.8000 161.8000 14.1000 ;
	    RECT 166.2000 10.8000 166.6000 12.7000 ;
	    RECT 168.6000 10.8000 169.0000 12.1000 ;
	    RECT 170.2000 10.8000 170.6000 13.1000 ;
	    RECT 0.2000 10.2000 173.4000 10.8000 ;
	    RECT 0.6000 7.9000 1.0000 10.2000 ;
	    RECT 3.0000 7.9000 3.4000 10.2000 ;
	    RECT 5.4000 7.9000 5.8000 10.2000 ;
	    RECT 9.4000 8.3000 9.8000 10.2000 ;
	    RECT 11.8000 8.9000 12.2000 10.2000 ;
	    RECT 12.6000 8.9000 13.0000 10.2000 ;
	    RECT 14.2000 8.1000 14.6000 10.2000 ;
	    RECT 16.6000 8.9000 17.0000 10.2000 ;
	    RECT 19.0000 7.9000 19.4000 10.2000 ;
	    RECT 20.6000 7.9000 21.0000 10.2000 ;
	    RECT 22.2000 7.9000 22.6000 10.2000 ;
	    RECT 25.4000 8.9000 25.8000 10.2000 ;
	    RECT 26.2000 7.9000 26.6000 10.2000 ;
	    RECT 28.6000 7.9000 29.0000 10.2000 ;
	    RECT 31.8000 8.9000 32.2000 10.2000 ;
	    RECT 32.6000 7.9000 33.0000 10.2000 ;
	    RECT 35.0000 7.9000 35.4000 10.2000 ;
	    RECT 37.4000 7.9000 37.8000 10.2000 ;
	    RECT 41.4000 8.3000 41.8000 10.2000 ;
	    RECT 43.8000 8.9000 44.2000 10.2000 ;
	    RECT 45.4000 8.9000 45.8000 10.2000 ;
	    RECT 46.2000 7.9000 46.6000 10.2000 ;
	    RECT 49.4000 8.9000 49.8000 10.2000 ;
	    RECT 51.0000 8.9000 51.4000 10.2000 ;
	    RECT 53.4000 7.9000 53.8000 10.2000 ;
	    RECT 54.2000 7.9000 54.6000 10.2000 ;
	    RECT 58.2000 7.9000 58.6000 10.2000 ;
	    RECT 59.8000 7.9000 60.2000 10.2000 ;
	    RECT 63.0000 7.9000 63.4000 10.2000 ;
	    RECT 65.4000 8.9000 65.8000 10.2000 ;
	    RECT 67.8000 8.9000 68.2000 10.2000 ;
	    RECT 70.2000 7.9000 70.6000 10.2000 ;
	    RECT 71.0000 7.9000 71.4000 10.2000 ;
	    RECT 74.2000 8.9000 74.6000 10.2000 ;
	    RECT 75.0000 7.9000 75.4000 10.2000 ;
	    RECT 78.2000 8.9000 78.6000 10.2000 ;
	    RECT 79.8000 7.9000 80.2000 10.2000 ;
	    RECT 81.4000 8.9000 81.8000 10.2000 ;
	    RECT 84.6000 7.9000 85.0000 10.2000 ;
	    RECT 85.4000 8.9000 85.8000 10.2000 ;
	    RECT 88.6000 7.9000 89.0000 10.2000 ;
	    RECT 89.4000 7.9000 89.8000 10.2000 ;
	    RECT 92.6000 8.9000 93.0000 10.2000 ;
	    RECT 93.4000 7.9000 93.8000 10.2000 ;
	    RECT 95.8000 8.9000 96.2000 10.2000 ;
	    RECT 99.0000 8.3000 99.4000 10.2000 ;
	    RECT 102.2000 7.9000 102.6000 10.2000 ;
	    RECT 103.0000 7.9000 103.4000 10.2000 ;
	    RECT 106.2000 8.9000 106.6000 10.2000 ;
	    RECT 107.0000 8.9000 107.4000 10.2000 ;
	    RECT 110.2000 7.9000 110.6000 10.2000 ;
	    RECT 112.6000 7.9000 113.0000 10.2000 ;
	    RECT 116.6000 8.3000 117.0000 10.2000 ;
	    RECT 119.0000 8.9000 119.4000 10.2000 ;
	    RECT 120.6000 7.9000 121.0000 10.2000 ;
	    RECT 122.2000 7.9000 122.6000 10.2000 ;
	    RECT 124.6000 7.9000 125.0000 10.2000 ;
	    RECT 127.8000 8.9000 128.2000 10.2000 ;
	    RECT 128.6000 8.9000 129.0000 10.2000 ;
	    RECT 130.2000 8.9000 130.6000 10.2000 ;
	    RECT 133.4000 7.9000 133.8000 10.2000 ;
	    RECT 134.2000 8.9000 134.6000 10.2000 ;
	    RECT 137.4000 7.9000 137.8000 10.2000 ;
	    RECT 139.8000 7.9000 140.2000 10.2000 ;
	    RECT 142.2000 7.9000 142.6000 10.2000 ;
	    RECT 143.0000 8.9000 143.4000 10.2000 ;
	    RECT 146.2000 7.9000 146.6000 10.2000 ;
	    RECT 148.6000 7.9000 149.0000 10.2000 ;
	    RECT 151.0000 7.9000 151.4000 10.2000 ;
	    RECT 151.8000 8.9000 152.2000 10.2000 ;
	    RECT 153.4000 8.1000 153.8000 10.2000 ;
	    RECT 155.0000 8.9000 155.4000 10.2000 ;
	    RECT 156.6000 8.1000 157.0000 10.2000 ;
	    RECT 159.0000 7.9000 159.4000 10.2000 ;
	    RECT 159.8000 7.9000 160.2000 10.2000 ;
	    RECT 161.4000 7.9000 161.8000 10.2000 ;
	    RECT 163.0000 7.9000 163.4000 10.2000 ;
	    RECT 164.6000 7.9000 165.0000 10.2000 ;
	    RECT 166.2000 7.9000 166.6000 10.2000 ;
	    RECT 167.8000 7.9000 168.2000 10.2000 ;
	    RECT 170.7000 8.0000 171.1000 10.2000 ;
         LAYER metal2 ;
	    RECT 111.2000 150.3000 112.8000 150.7000 ;
	    RECT 111.2000 130.3000 112.8000 130.7000 ;
	    RECT 111.2000 110.3000 112.8000 110.7000 ;
	    RECT 111.2000 90.3000 112.8000 90.7000 ;
	    RECT 111.2000 70.3000 112.8000 70.7000 ;
	    RECT 111.2000 50.3000 112.8000 50.7000 ;
	    RECT 111.2000 30.3000 112.8000 30.7000 ;
	    RECT 111.2000 10.3000 112.8000 10.7000 ;
         LAYER metal3 ;
	    RECT 111.2000 150.3000 112.8000 150.7000 ;
	    RECT 111.2000 130.3000 112.8000 130.7000 ;
	    RECT 111.2000 110.3000 112.8000 110.7000 ;
	    RECT 111.2000 90.3000 112.8000 90.7000 ;
	    RECT 111.2000 70.3000 112.8000 70.7000 ;
	    RECT 111.2000 50.3000 112.8000 50.7000 ;
	    RECT 111.2000 30.3000 112.8000 30.7000 ;
	    RECT 111.2000 10.3000 112.8000 10.7000 ;
         LAYER metal4 ;
	    RECT 111.2000 150.3000 112.8000 150.7000 ;
	    RECT 111.2000 130.3000 112.8000 130.7000 ;
	    RECT 111.2000 110.3000 112.8000 110.7000 ;
	    RECT 111.2000 90.3000 112.8000 90.7000 ;
	    RECT 111.2000 70.3000 112.8000 70.7000 ;
	    RECT 111.2000 50.3000 112.8000 50.7000 ;
	    RECT 111.2000 30.3000 112.8000 30.7000 ;
	    RECT 111.2000 10.3000 112.8000 10.7000 ;
         LAYER metal5 ;
	    RECT 111.2000 150.7000 111.8000 150.8000 ;
	    RECT 112.2000 150.7000 112.8000 150.8000 ;
	    RECT 111.2000 150.2000 112.8000 150.7000 ;
	    RECT 111.2000 130.7000 111.8000 130.8000 ;
	    RECT 112.2000 130.7000 112.8000 130.8000 ;
	    RECT 111.2000 130.2000 112.8000 130.7000 ;
	    RECT 111.2000 110.7000 111.8000 110.8000 ;
	    RECT 112.2000 110.7000 112.8000 110.8000 ;
	    RECT 111.2000 110.2000 112.8000 110.7000 ;
	    RECT 111.2000 90.7000 111.8000 90.8000 ;
	    RECT 112.2000 90.7000 112.8000 90.8000 ;
	    RECT 111.2000 90.2000 112.8000 90.7000 ;
	    RECT 111.2000 70.7000 111.8000 70.8000 ;
	    RECT 112.2000 70.7000 112.8000 70.8000 ;
	    RECT 111.2000 70.2000 112.8000 70.7000 ;
	    RECT 111.2000 50.7000 111.8000 50.8000 ;
	    RECT 112.2000 50.7000 112.8000 50.8000 ;
	    RECT 111.2000 50.2000 112.8000 50.7000 ;
	    RECT 111.2000 30.7000 111.8000 30.8000 ;
	    RECT 112.2000 30.7000 112.8000 30.8000 ;
	    RECT 111.2000 30.2000 112.8000 30.7000 ;
	    RECT 111.2000 10.7000 111.8000 10.8000 ;
	    RECT 112.2000 10.7000 112.8000 10.8000 ;
	    RECT 111.2000 10.2000 112.8000 10.7000 ;
         LAYER metal6 ;
	    RECT 111.2000 -3.0000 112.8000 164.0000 ;
      END
   END gnd
   PIN CLK
      PORT
         LAYER metal1 ;
	    RECT 158.5000 94.1000 159.4000 94.5000 ;
	    RECT 159.0000 93.8000 159.4000 94.1000 ;
	    RECT 145.4000 86.9000 145.8000 87.2000 ;
	    RECT 145.4000 86.5000 146.3000 86.9000 ;
	    RECT 108.9000 74.1000 109.8000 74.5000 ;
	    RECT 109.4000 73.8000 109.8000 74.1000 ;
	    RECT 111.0000 67.1000 111.4000 67.2000 ;
	    RECT 112.6000 67.1000 113.0000 67.2000 ;
	    RECT 111.0000 66.9000 113.0000 67.1000 ;
	    RECT 111.0000 66.8000 113.5000 66.9000 ;
	    RECT 112.6000 66.5000 113.5000 66.8000 ;
	    RECT 107.3000 54.1000 108.2000 54.5000 ;
	    RECT 107.8000 53.8000 108.2000 54.1000 ;
	    RECT 166.2000 6.9000 166.6000 7.2000 ;
	    RECT 165.7000 6.5000 166.6000 6.9000 ;
         LAYER metal2 ;
	    RECT 159.0000 93.8000 159.4000 94.2000 ;
	    RECT 159.0000 91.2000 159.3000 93.8000 ;
	    RECT 145.4000 90.8000 145.8000 91.2000 ;
	    RECT 159.0000 90.8000 159.4000 91.2000 ;
	    RECT 145.4000 87.2000 145.7000 90.8000 ;
	    RECT 145.4000 86.8000 145.8000 87.2000 ;
	    RECT 145.4000 84.2000 145.7000 86.8000 ;
	    RECT 109.4000 83.8000 109.8000 84.2000 ;
	    RECT 145.4000 83.8000 145.8000 84.2000 ;
	    RECT 109.4000 74.2000 109.7000 83.8000 ;
	    RECT 109.4000 73.8000 109.8000 74.2000 ;
	    RECT 109.4000 64.2000 109.7000 73.8000 ;
	    RECT 111.0000 66.8000 111.4000 67.2000 ;
	    RECT 111.0000 64.2000 111.3000 66.8000 ;
	    RECT 109.4000 63.8000 109.8000 64.2000 ;
	    RECT 111.0000 63.8000 111.4000 64.2000 ;
	    RECT 109.4000 58.2000 109.7000 63.8000 ;
	    RECT 107.8000 57.8000 108.2000 58.2000 ;
	    RECT 109.4000 57.8000 109.8000 58.2000 ;
	    RECT 107.8000 54.2000 108.1000 57.8000 ;
	    RECT 107.8000 53.8000 108.2000 54.2000 ;
	    RECT 166.2000 7.8000 166.6000 8.2000 ;
	    RECT 166.2000 7.2000 166.5000 7.8000 ;
	    RECT 166.2000 6.8000 166.6000 7.2000 ;
         LAYER metal3 ;
	    RECT 145.4000 91.1000 145.8000 91.2000 ;
	    RECT 159.0000 91.1000 159.4000 91.2000 ;
	    RECT 163.8000 91.1000 164.2000 91.2000 ;
	    RECT 145.4000 90.8000 164.2000 91.1000 ;
	    RECT 109.4000 84.1000 109.8000 84.2000 ;
	    RECT 145.4000 84.1000 145.8000 84.2000 ;
	    RECT 109.4000 83.8000 145.8000 84.1000 ;
	    RECT 163.8000 66.1000 164.2000 66.2000 ;
	    RECT 166.2000 66.1000 166.6000 66.2000 ;
	    RECT 175.8000 66.1000 176.2000 66.2000 ;
	    RECT 163.8000 65.8000 176.2000 66.1000 ;
	    RECT 109.4000 64.1000 109.8000 64.2000 ;
	    RECT 111.0000 64.1000 111.4000 64.2000 ;
	    RECT 109.4000 63.8000 111.4000 64.1000 ;
	    RECT 107.8000 58.1000 108.2000 58.2000 ;
	    RECT 109.4000 58.1000 109.8000 58.2000 ;
	    RECT 107.8000 57.8000 109.8000 58.1000 ;
	    RECT 166.2000 7.8000 166.6000 8.2000 ;
	    RECT 166.2000 7.2000 166.5000 7.8000 ;
	    RECT 166.2000 6.8000 166.6000 7.2000 ;
         LAYER metal4 ;
	    RECT 163.8000 90.8000 164.2000 91.2000 ;
	    RECT 163.8000 66.2000 164.1000 90.8000 ;
	    RECT 163.8000 65.8000 164.2000 66.2000 ;
	    RECT 166.2000 65.8000 166.6000 66.2000 ;
	    RECT 166.2000 7.2000 166.5000 65.8000 ;
	    RECT 166.2000 6.8000 166.6000 7.2000 ;
      END
   END CLK
   PIN DATA_A[31]
      PORT
         LAYER metal1 ;
	    RECT 21.4000 63.8000 21.8000 65.2000 ;
	    RECT 39.0000 65.1000 39.4000 65.2000 ;
	    RECT 39.8000 65.1000 40.2000 65.2000 ;
	    RECT 39.0000 64.8000 40.2000 65.1000 ;
	    RECT 39.0000 64.4000 39.4000 64.8000 ;
	    RECT 39.8000 64.4000 40.2000 64.8000 ;
	    RECT 47.0000 64.4000 47.4000 65.2000 ;
         LAYER metal2 ;
	    RECT 47.0000 65.8000 47.4000 66.2000 ;
	    RECT 47.0000 65.2000 47.3000 65.8000 ;
	    RECT 0.6000 64.8000 1.0000 65.2000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 39.0000 65.1000 39.4000 65.2000 ;
	    RECT 38.2000 64.8000 39.4000 65.1000 ;
	    RECT 47.0000 64.8000 47.4000 65.2000 ;
	    RECT 0.6000 63.2000 0.9000 64.8000 ;
	    RECT 21.4000 63.8000 21.8000 64.2000 ;
	    RECT 21.4000 63.2000 21.7000 63.8000 ;
	    RECT 0.6000 62.8000 1.0000 63.2000 ;
	    RECT 21.4000 62.8000 21.8000 63.2000 ;
         LAYER metal3 ;
	    RECT 47.0000 65.8000 47.4000 66.2000 ;
	    RECT -2.6000 65.1000 -2.2000 65.2000 ;
	    RECT 0.6000 65.1000 1.0000 65.2000 ;
	    RECT -2.6000 64.8000 1.0000 65.1000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 39.0000 65.1000 39.4000 65.2000 ;
	    RECT 47.0000 65.1000 47.3000 65.8000 ;
	    RECT 38.2000 64.8000 47.3000 65.1000 ;
	    RECT 0.6000 63.1000 1.0000 63.2000 ;
	    RECT 21.4000 63.1000 21.8000 63.2000 ;
	    RECT 23.8000 63.1000 24.2000 63.2000 ;
	    RECT 0.6000 62.8000 24.2000 63.1000 ;
         LAYER metal4 ;
	    RECT 23.8000 64.8000 24.2000 65.2000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 39.0000 65.1000 39.4000 65.2000 ;
	    RECT 38.2000 64.8000 39.4000 65.1000 ;
	    RECT 23.8000 63.2000 24.1000 64.8000 ;
	    RECT 23.8000 62.8000 24.2000 63.2000 ;
         LAYER metal5 ;
	    RECT 23.8000 65.1000 24.2000 65.2000 ;
	    RECT 38.2000 65.1000 38.6000 65.2000 ;
	    RECT 23.8000 64.8000 38.6000 65.1000 ;
      END
   END DATA_A[31]
   PIN DATA_A[30]
      PORT
         LAYER metal1 ;
	    RECT 37.4000 156.8000 37.8000 157.2000 ;
	    RECT 6.2000 155.8000 6.6000 156.6000 ;
	    RECT 11.8000 155.8000 12.2000 156.6000 ;
	    RECT 35.8000 155.8000 36.2000 156.6000 ;
	    RECT 37.4000 156.1000 37.7000 156.8000 ;
	    RECT 38.2000 156.1000 38.6000 156.6000 ;
	    RECT 37.4000 155.8000 38.6000 156.1000 ;
         LAYER metal2 ;
	    RECT 6.2000 163.8000 6.6000 164.2000 ;
	    RECT 6.2000 159.2000 6.5000 163.8000 ;
	    RECT 6.2000 158.8000 6.6000 159.2000 ;
	    RECT 11.8000 158.8000 12.2000 159.2000 ;
	    RECT 35.8000 158.8000 36.2000 159.2000 ;
	    RECT 6.2000 156.2000 6.5000 158.8000 ;
	    RECT 11.8000 156.2000 12.1000 158.8000 ;
	    RECT 35.8000 156.2000 36.1000 158.8000 ;
	    RECT 37.4000 156.8000 37.8000 157.2000 ;
	    RECT 37.4000 156.2000 37.7000 156.8000 ;
	    RECT 6.2000 155.8000 6.6000 156.2000 ;
	    RECT 11.8000 155.8000 12.2000 156.2000 ;
	    RECT 35.8000 156.1000 36.2000 156.2000 ;
	    RECT 36.6000 156.1000 37.0000 156.2000 ;
	    RECT 35.8000 155.8000 37.0000 156.1000 ;
	    RECT 37.4000 155.8000 37.8000 156.2000 ;
         LAYER metal3 ;
	    RECT 6.2000 159.1000 6.6000 159.2000 ;
	    RECT 11.8000 159.1000 12.2000 159.2000 ;
	    RECT 35.8000 159.1000 36.2000 159.2000 ;
	    RECT 6.2000 158.8000 36.2000 159.1000 ;
	    RECT 36.6000 156.1000 37.0000 156.2000 ;
	    RECT 37.4000 156.1000 37.8000 156.2000 ;
	    RECT 36.6000 155.8000 37.8000 156.1000 ;
      END
   END DATA_A[30]
   PIN DATA_A[29]
      PORT
         LAYER metal1 ;
	    RECT 27.8000 157.1000 28.2000 157.2000 ;
	    RECT 27.0000 156.8000 28.2000 157.1000 ;
	    RECT 27.0000 155.8000 27.4000 156.8000 ;
	    RECT 44.6000 155.8000 45.0000 156.6000 ;
	    RECT 44.6000 135.8000 45.0000 136.6000 ;
	    RECT 50.2000 135.8000 50.6000 136.6000 ;
         LAYER metal2 ;
	    RECT 44.6000 163.8000 45.0000 164.2000 ;
	    RECT 44.6000 161.2000 44.9000 163.8000 ;
	    RECT 27.8000 160.8000 28.2000 161.2000 ;
	    RECT 44.6000 160.8000 45.0000 161.2000 ;
	    RECT 27.8000 157.2000 28.1000 160.8000 ;
	    RECT 27.8000 156.8000 28.2000 157.2000 ;
	    RECT 44.6000 156.2000 44.9000 160.8000 ;
	    RECT 44.6000 155.8000 45.0000 156.2000 ;
	    RECT 44.6000 136.8000 45.0000 137.2000 ;
	    RECT 50.2000 136.8000 50.6000 137.2000 ;
	    RECT 44.6000 136.2000 44.9000 136.8000 ;
	    RECT 50.2000 136.2000 50.5000 136.8000 ;
	    RECT 44.6000 135.8000 45.0000 136.2000 ;
	    RECT 50.2000 135.8000 50.6000 136.2000 ;
         LAYER metal3 ;
	    RECT 27.8000 161.1000 28.2000 161.2000 ;
	    RECT 44.6000 161.1000 45.0000 161.2000 ;
	    RECT 27.8000 160.8000 45.0000 161.1000 ;
	    RECT 44.6000 137.1000 45.0000 137.2000 ;
	    RECT 50.2000 137.1000 50.6000 137.2000 ;
	    RECT 44.6000 136.8000 50.6000 137.1000 ;
	    RECT 44.6000 136.2000 44.9000 136.8000 ;
	    RECT 44.6000 135.8000 45.0000 136.2000 ;
         LAYER metal4 ;
	    RECT 44.6000 160.8000 45.0000 161.2000 ;
	    RECT 44.6000 136.2000 44.9000 160.8000 ;
	    RECT 44.6000 135.8000 45.0000 136.2000 ;
      END
   END DATA_A[29]
   PIN DATA_A[28]
      PORT
         LAYER metal1 ;
	    RECT 15.8000 155.8000 16.2000 156.6000 ;
	    RECT 20.6000 155.8000 21.0000 156.6000 ;
	    RECT 53.4000 155.8000 53.8000 156.6000 ;
	    RECT 63.0000 155.8000 63.4000 156.6000 ;
	    RECT 15.8000 155.2000 16.1000 155.8000 ;
	    RECT 15.8000 154.8000 16.2000 155.2000 ;
         LAYER metal2 ;
	    RECT 64.6000 163.8000 65.0000 164.2000 ;
	    RECT 64.6000 158.2000 64.9000 163.8000 ;
	    RECT 53.4000 157.8000 53.8000 158.2000 ;
	    RECT 63.0000 157.8000 63.4000 158.2000 ;
	    RECT 64.6000 157.8000 65.0000 158.2000 ;
	    RECT 20.6000 156.8000 21.0000 157.2000 ;
	    RECT 20.6000 156.2000 20.9000 156.8000 ;
	    RECT 53.4000 156.2000 53.7000 157.8000 ;
	    RECT 63.0000 156.2000 63.3000 157.8000 ;
	    RECT 15.8000 155.8000 16.2000 156.2000 ;
	    RECT 20.6000 155.8000 21.0000 156.2000 ;
	    RECT 53.4000 155.8000 53.8000 156.2000 ;
	    RECT 63.0000 155.8000 63.4000 156.2000 ;
	    RECT 15.8000 155.2000 16.1000 155.8000 ;
	    RECT 15.8000 154.8000 16.2000 155.2000 ;
         LAYER metal3 ;
	    RECT 53.4000 158.1000 53.8000 158.2000 ;
	    RECT 63.0000 158.1000 63.4000 158.2000 ;
	    RECT 64.6000 158.1000 65.0000 158.2000 ;
	    RECT 20.6000 157.8000 65.0000 158.1000 ;
	    RECT 20.6000 157.2000 20.9000 157.8000 ;
	    RECT 20.6000 156.8000 21.0000 157.2000 ;
	    RECT 15.8000 156.1000 16.2000 156.2000 ;
	    RECT 20.6000 156.1000 20.9000 156.8000 ;
	    RECT 15.8000 155.8000 20.9000 156.1000 ;
      END
   END DATA_A[28]
   PIN DATA_A[27]
      PORT
         LAYER metal1 ;
	    RECT 21.4000 73.8000 21.8000 74.2000 ;
	    RECT 21.4000 73.2000 21.7000 73.8000 ;
	    RECT 21.4000 72.4000 21.8000 73.2000 ;
	    RECT 26.2000 72.4000 26.6000 73.2000 ;
	    RECT 83.8000 72.4000 84.2000 73.2000 ;
	    RECT 69.4000 67.8000 69.8000 68.6000 ;
         LAYER metal2 ;
	    RECT 11.0000 77.8000 11.4000 78.2000 ;
	    RECT 11.0000 73.2000 11.3000 77.8000 ;
	    RECT 21.4000 73.8000 21.8000 74.2000 ;
	    RECT 69.4000 73.8000 69.8000 74.2000 ;
	    RECT 83.8000 73.8000 84.2000 74.2000 ;
	    RECT 21.4000 73.2000 21.7000 73.8000 ;
	    RECT 11.0000 72.8000 11.4000 73.2000 ;
	    RECT 21.4000 72.8000 21.8000 73.2000 ;
	    RECT 26.2000 73.1000 26.6000 73.2000 ;
	    RECT 27.0000 73.1000 27.4000 73.2000 ;
	    RECT 26.2000 72.8000 27.4000 73.1000 ;
	    RECT 69.4000 68.2000 69.7000 73.8000 ;
	    RECT 83.8000 73.2000 84.1000 73.8000 ;
	    RECT 83.8000 72.8000 84.2000 73.2000 ;
	    RECT 69.4000 67.8000 69.8000 68.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 78.1000 -2.2000 78.2000 ;
	    RECT 11.0000 78.1000 11.4000 78.2000 ;
	    RECT -2.6000 77.8000 11.4000 78.1000 ;
	    RECT 69.4000 74.1000 69.8000 74.2000 ;
	    RECT 83.8000 74.1000 84.2000 74.2000 ;
	    RECT 27.0000 73.8000 84.2000 74.1000 ;
	    RECT 27.0000 73.2000 27.3000 73.8000 ;
	    RECT 11.0000 73.1000 11.4000 73.2000 ;
	    RECT 21.4000 73.1000 21.8000 73.2000 ;
	    RECT 27.0000 73.1000 27.4000 73.2000 ;
	    RECT 11.0000 72.8000 27.4000 73.1000 ;
      END
   END DATA_A[27]
   PIN DATA_A[26]
      PORT
         LAYER metal1 ;
	    RECT 55.0000 112.4000 55.4000 113.2000 ;
	    RECT 34.2000 107.8000 34.6000 108.6000 ;
	    RECT 54.2000 67.8000 54.6000 68.6000 ;
	    RECT 7.8000 47.8000 8.2000 48.6000 ;
         LAYER metal2 ;
	    RECT 55.0000 112.8000 55.4000 113.2000 ;
	    RECT 55.0000 112.2000 55.3000 112.8000 ;
	    RECT 55.0000 111.8000 55.4000 112.2000 ;
	    RECT 33.4000 108.1000 33.8000 108.2000 ;
	    RECT 34.2000 108.1000 34.6000 108.2000 ;
	    RECT 33.4000 107.8000 34.6000 108.1000 ;
	    RECT 54.2000 74.8000 54.6000 75.2000 ;
	    RECT 54.2000 68.2000 54.5000 74.8000 ;
	    RECT 54.2000 67.8000 54.6000 68.2000 ;
	    RECT 7.8000 48.8000 8.2000 49.2000 ;
	    RECT 7.8000 48.2000 8.1000 48.8000 ;
	    RECT 7.8000 47.8000 8.2000 48.2000 ;
         LAYER metal3 ;
	    RECT 55.0000 111.8000 55.4000 112.2000 ;
	    RECT 55.0000 111.2000 55.3000 111.8000 ;
	    RECT 55.0000 110.8000 55.4000 111.2000 ;
	    RECT 33.4000 108.1000 33.8000 108.2000 ;
	    RECT 55.0000 108.1000 55.4000 108.2000 ;
	    RECT 33.4000 107.8000 55.4000 108.1000 ;
	    RECT 54.2000 75.1000 54.6000 75.2000 ;
	    RECT 55.0000 75.1000 55.4000 75.2000 ;
	    RECT 54.2000 74.8000 55.4000 75.1000 ;
	    RECT -2.6000 58.1000 -2.2000 58.2000 ;
	    RECT 0.6000 58.1000 1.0000 58.2000 ;
	    RECT -2.6000 57.8000 1.0000 58.1000 ;
	    RECT 7.8000 49.8000 8.2000 50.2000 ;
	    RECT 7.8000 49.2000 8.1000 49.8000 ;
	    RECT 7.8000 48.8000 8.2000 49.2000 ;
         LAYER metal4 ;
	    RECT 55.0000 110.8000 55.4000 111.2000 ;
	    RECT 55.0000 108.2000 55.3000 110.8000 ;
	    RECT 55.0000 107.8000 55.4000 108.2000 ;
	    RECT 55.0000 75.2000 55.3000 107.8000 ;
	    RECT 55.0000 74.8000 55.4000 75.2000 ;
	    RECT 55.0000 58.2000 55.3000 74.8000 ;
	    RECT 0.6000 58.1000 1.0000 58.2000 ;
	    RECT 1.4000 58.1000 1.8000 58.2000 ;
	    RECT 0.6000 57.8000 1.8000 58.1000 ;
	    RECT 7.8000 57.8000 8.2000 58.2000 ;
	    RECT 55.0000 57.8000 55.4000 58.2000 ;
	    RECT 7.8000 50.2000 8.1000 57.8000 ;
	    RECT 7.8000 49.8000 8.2000 50.2000 ;
         LAYER metal5 ;
	    RECT 1.4000 58.1000 1.8000 58.2000 ;
	    RECT 7.8000 58.1000 8.2000 58.2000 ;
	    RECT 55.0000 58.1000 55.4000 58.2000 ;
	    RECT 1.4000 57.8000 55.4000 58.1000 ;
      END
   END DATA_A[26]
   PIN DATA_A[25]
      PORT
         LAYER metal1 ;
	    RECT 34.2000 72.4000 34.6000 73.2000 ;
	    RECT 85.4000 72.4000 85.8000 73.2000 ;
	    RECT 73.4000 67.8000 73.8000 68.6000 ;
	    RECT 13.4000 47.8000 13.8000 48.6000 ;
         LAYER metal2 ;
	    RECT 34.2000 73.1000 34.6000 73.2000 ;
	    RECT 35.0000 73.1000 35.4000 73.2000 ;
	    RECT 34.2000 72.8000 35.4000 73.1000 ;
	    RECT 85.4000 72.8000 85.8000 73.2000 ;
	    RECT 85.4000 71.2000 85.7000 72.8000 ;
	    RECT 73.4000 70.8000 73.8000 71.2000 ;
	    RECT 85.4000 70.8000 85.8000 71.2000 ;
	    RECT 73.4000 68.2000 73.7000 70.8000 ;
	    RECT 73.4000 67.8000 73.8000 68.2000 ;
	    RECT 73.4000 63.2000 73.7000 67.8000 ;
	    RECT 73.4000 62.8000 73.8000 63.2000 ;
	    RECT 13.4000 59.8000 13.8000 60.2000 ;
	    RECT 13.4000 52.2000 13.7000 59.8000 ;
	    RECT 13.4000 51.8000 13.8000 52.2000 ;
	    RECT 13.4000 48.2000 13.7000 51.8000 ;
	    RECT 13.4000 47.8000 13.8000 48.2000 ;
         LAYER metal3 ;
	    RECT 34.2000 73.1000 34.6000 73.2000 ;
	    RECT 35.0000 73.1000 35.4000 73.2000 ;
	    RECT 34.2000 72.8000 35.4000 73.1000 ;
	    RECT 73.4000 71.1000 73.8000 71.2000 ;
	    RECT 85.4000 71.1000 85.8000 71.2000 ;
	    RECT 73.4000 70.8000 85.8000 71.1000 ;
	    RECT 34.2000 63.1000 34.6000 63.2000 ;
	    RECT 73.4000 63.1000 73.8000 63.2000 ;
	    RECT 34.2000 62.8000 73.8000 63.1000 ;
	    RECT 13.4000 60.1000 13.8000 60.2000 ;
	    RECT 34.2000 60.1000 34.6000 60.2000 ;
	    RECT 13.4000 59.8000 34.6000 60.1000 ;
	    RECT -2.6000 56.1000 -2.2000 56.2000 ;
	    RECT 0.6000 56.1000 1.0000 56.2000 ;
	    RECT -2.6000 55.8000 1.0000 56.1000 ;
	    RECT 0.6000 52.1000 1.0000 52.2000 ;
	    RECT 13.4000 52.1000 13.8000 52.2000 ;
	    RECT 0.6000 51.8000 13.8000 52.1000 ;
         LAYER metal4 ;
	    RECT 34.2000 72.8000 34.6000 73.2000 ;
	    RECT 34.2000 63.2000 34.5000 72.8000 ;
	    RECT 34.2000 62.8000 34.6000 63.2000 ;
	    RECT 34.2000 60.2000 34.5000 62.8000 ;
	    RECT 34.2000 59.8000 34.6000 60.2000 ;
	    RECT 0.6000 55.8000 1.0000 56.2000 ;
	    RECT 0.6000 52.2000 0.9000 55.8000 ;
	    RECT 0.6000 51.8000 1.0000 52.2000 ;
      END
   END DATA_A[25]
   PIN DATA_A[24]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 107.8000 1.0000 108.6000 ;
	    RECT 45.4000 107.8000 45.8000 108.6000 ;
	    RECT 63.0000 92.4000 63.4000 93.2000 ;
	    RECT 5.4000 87.8000 5.8000 88.6000 ;
         LAYER metal2 ;
	    RECT 0.6000 109.8000 1.0000 110.2000 ;
	    RECT 6.2000 109.8000 6.6000 110.2000 ;
	    RECT 0.6000 108.2000 0.9000 109.8000 ;
	    RECT 0.6000 107.8000 1.0000 108.2000 ;
	    RECT 6.2000 102.2000 6.5000 109.8000 ;
	    RECT 45.4000 107.8000 45.8000 108.2000 ;
	    RECT 45.4000 102.2000 45.7000 107.8000 ;
	    RECT 6.2000 101.8000 6.6000 102.2000 ;
	    RECT 45.4000 101.8000 45.8000 102.2000 ;
	    RECT 63.0000 101.8000 63.4000 102.2000 ;
	    RECT 6.2000 95.1000 6.5000 101.8000 ;
	    RECT 5.4000 94.8000 6.5000 95.1000 ;
	    RECT 5.4000 88.2000 5.7000 94.8000 ;
	    RECT 63.0000 93.2000 63.3000 101.8000 ;
	    RECT 63.0000 92.8000 63.4000 93.2000 ;
	    RECT 5.4000 87.8000 5.8000 88.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 110.1000 -2.2000 110.2000 ;
	    RECT 0.6000 110.1000 1.0000 110.2000 ;
	    RECT 6.2000 110.1000 6.6000 110.2000 ;
	    RECT -2.6000 109.8000 6.6000 110.1000 ;
	    RECT 6.2000 102.1000 6.6000 102.2000 ;
	    RECT 45.4000 102.1000 45.8000 102.2000 ;
	    RECT 63.0000 102.1000 63.4000 102.2000 ;
	    RECT 6.2000 101.8000 63.4000 102.1000 ;
      END
   END DATA_A[24]
   PIN DATA_A[23]
      PORT
         LAYER metal1 ;
	    RECT 49.4000 92.4000 49.8000 93.2000 ;
	    RECT 15.8000 87.8000 16.2000 88.6000 ;
	    RECT 47.0000 87.8000 47.4000 88.6000 ;
	    RECT 11.8000 72.4000 12.2000 73.2000 ;
         LAYER metal2 ;
	    RECT 49.4000 92.8000 49.8000 93.2000 ;
	    RECT 49.4000 90.2000 49.7000 92.8000 ;
	    RECT 47.0000 89.8000 47.4000 90.2000 ;
	    RECT 49.4000 89.8000 49.8000 90.2000 ;
	    RECT 47.0000 88.2000 47.3000 89.8000 ;
	    RECT 11.8000 87.8000 12.2000 88.2000 ;
	    RECT 15.0000 88.1000 15.4000 88.2000 ;
	    RECT 15.8000 88.1000 16.2000 88.2000 ;
	    RECT 15.0000 87.8000 16.2000 88.1000 ;
	    RECT 47.0000 87.8000 47.4000 88.2000 ;
	    RECT 11.8000 83.2000 12.1000 87.8000 ;
	    RECT 15.8000 84.2000 16.1000 87.8000 ;
	    RECT 47.0000 84.2000 47.3000 87.8000 ;
	    RECT 15.8000 83.8000 16.2000 84.2000 ;
	    RECT 47.0000 83.8000 47.4000 84.2000 ;
	    RECT 11.8000 82.8000 12.2000 83.2000 ;
	    RECT 11.8000 73.2000 12.1000 82.8000 ;
	    RECT 11.8000 72.8000 12.2000 73.2000 ;
         LAYER metal3 ;
	    RECT 47.0000 90.1000 47.4000 90.2000 ;
	    RECT 49.4000 90.1000 49.8000 90.2000 ;
	    RECT 47.0000 89.8000 49.8000 90.1000 ;
	    RECT 11.8000 88.1000 12.2000 88.2000 ;
	    RECT 15.0000 88.1000 15.4000 88.2000 ;
	    RECT 11.8000 87.8000 15.4000 88.1000 ;
	    RECT 15.8000 84.1000 16.2000 84.2000 ;
	    RECT 47.0000 84.1000 47.4000 84.2000 ;
	    RECT 15.8000 83.8000 47.4000 84.1000 ;
	    RECT 11.8000 83.1000 12.2000 83.2000 ;
	    RECT -0.2000 82.8000 12.2000 83.1000 ;
	    RECT -2.6000 82.1000 -2.2000 82.2000 ;
	    RECT -0.2000 82.1000 0.1000 82.8000 ;
	    RECT -2.6000 81.8000 0.1000 82.1000 ;
      END
   END DATA_A[23]
   PIN DATA_A[22]
      PORT
         LAYER metal1 ;
	    RECT 0.6000 152.4000 1.0000 153.2000 ;
	    RECT 48.6000 152.4000 49.0000 153.2000 ;
	    RECT 18.2000 147.8000 18.6000 148.6000 ;
	    RECT 50.2000 147.8000 50.6000 148.6000 ;
         LAYER metal2 ;
	    RECT 0.6000 152.8000 1.0000 153.2000 ;
	    RECT 48.6000 152.8000 49.0000 153.2000 ;
	    RECT 0.6000 152.2000 0.9000 152.8000 ;
	    RECT 0.6000 151.8000 1.0000 152.2000 ;
	    RECT 18.2000 151.8000 18.6000 152.2000 ;
	    RECT 0.6000 146.2000 0.9000 151.8000 ;
	    RECT 18.2000 148.2000 18.5000 151.8000 ;
	    RECT 48.6000 149.2000 48.9000 152.8000 ;
	    RECT 48.6000 148.8000 49.0000 149.2000 ;
	    RECT 50.2000 148.8000 50.6000 149.2000 ;
	    RECT 50.2000 148.2000 50.5000 148.8000 ;
	    RECT 18.2000 147.8000 18.6000 148.2000 ;
	    RECT 50.2000 147.8000 50.6000 148.2000 ;
	    RECT 0.6000 145.8000 1.0000 146.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 152.1000 1.0000 152.2000 ;
	    RECT 18.2000 152.1000 18.6000 152.2000 ;
	    RECT 36.6000 152.1000 37.0000 152.2000 ;
	    RECT 0.6000 151.8000 37.0000 152.1000 ;
	    RECT 36.6000 149.1000 37.0000 149.2000 ;
	    RECT 48.6000 149.1000 49.0000 149.2000 ;
	    RECT 50.2000 149.1000 50.6000 149.2000 ;
	    RECT 36.6000 148.8000 50.6000 149.1000 ;
	    RECT -2.6000 146.1000 -2.2000 146.2000 ;
	    RECT 0.6000 146.1000 1.0000 146.2000 ;
	    RECT -2.6000 145.8000 1.0000 146.1000 ;
         LAYER metal4 ;
	    RECT 36.6000 151.8000 37.0000 152.2000 ;
	    RECT 36.6000 149.2000 36.9000 151.8000 ;
	    RECT 36.6000 148.8000 37.0000 149.2000 ;
      END
   END DATA_A[22]
   PIN DATA_A[21]
      PORT
         LAYER metal1 ;
	    RECT 75.0000 152.4000 75.4000 153.2000 ;
	    RECT 27.0000 132.4000 27.4000 133.2000 ;
	    RECT 40.6000 127.8000 41.0000 128.6000 ;
	    RECT 76.6000 127.8000 77.0000 128.6000 ;
         LAYER metal2 ;
	    RECT 76.6000 163.8000 77.0000 164.2000 ;
	    RECT 76.6000 153.2000 76.9000 163.8000 ;
	    RECT 74.2000 153.1000 74.6000 153.2000 ;
	    RECT 75.0000 153.1000 75.4000 153.2000 ;
	    RECT 74.2000 152.8000 75.4000 153.1000 ;
	    RECT 76.6000 152.8000 77.0000 153.2000 ;
	    RECT 27.0000 132.8000 27.4000 133.2000 ;
	    RECT 27.0000 128.2000 27.3000 132.8000 ;
	    RECT 40.6000 130.8000 41.0000 131.2000 ;
	    RECT 76.6000 130.8000 77.0000 131.2000 ;
	    RECT 40.6000 128.2000 40.9000 130.8000 ;
	    RECT 76.6000 128.2000 76.9000 130.8000 ;
	    RECT 27.0000 127.8000 27.4000 128.2000 ;
	    RECT 39.8000 128.1000 40.2000 128.2000 ;
	    RECT 40.6000 128.1000 41.0000 128.2000 ;
	    RECT 39.8000 127.8000 41.0000 128.1000 ;
	    RECT 76.6000 127.8000 77.0000 128.2000 ;
         LAYER metal3 ;
	    RECT 74.2000 153.1000 74.6000 153.2000 ;
	    RECT 76.6000 153.1000 77.0000 153.2000 ;
	    RECT 74.2000 152.8000 77.0000 153.1000 ;
	    RECT 74.2000 152.2000 74.5000 152.8000 ;
	    RECT 74.2000 151.8000 74.6000 152.2000 ;
	    RECT 40.6000 131.1000 41.0000 131.2000 ;
	    RECT 74.2000 131.1000 74.6000 131.2000 ;
	    RECT 76.6000 131.1000 77.0000 131.2000 ;
	    RECT 40.6000 130.8000 77.0000 131.1000 ;
	    RECT 27.0000 128.1000 27.4000 128.2000 ;
	    RECT 39.8000 128.1000 40.2000 128.2000 ;
	    RECT 27.0000 127.8000 40.2000 128.1000 ;
         LAYER metal4 ;
	    RECT 74.2000 151.8000 74.6000 152.2000 ;
	    RECT 74.2000 131.2000 74.5000 151.8000 ;
	    RECT 74.2000 130.8000 74.6000 131.2000 ;
      END
   END DATA_A[21]
   PIN DATA_A[20]
      PORT
         LAYER metal1 ;
	    RECT 24.6000 152.4000 25.0000 153.2000 ;
	    RECT 68.6000 152.4000 69.0000 153.2000 ;
	    RECT 31.0000 147.8000 31.4000 148.6000 ;
	    RECT 71.0000 147.8000 71.4000 148.6000 ;
         LAYER metal2 ;
	    RECT 72.6000 163.8000 73.0000 164.2000 ;
	    RECT 72.6000 157.2000 72.9000 163.8000 ;
	    RECT 24.6000 156.8000 25.0000 157.2000 ;
	    RECT 68.6000 156.8000 69.0000 157.2000 ;
	    RECT 72.6000 156.8000 73.0000 157.2000 ;
	    RECT 24.6000 153.2000 24.9000 156.8000 ;
	    RECT 68.6000 153.2000 68.9000 156.8000 ;
	    RECT 24.6000 152.8000 25.0000 153.2000 ;
	    RECT 68.6000 152.8000 69.0000 153.2000 ;
	    RECT 24.6000 148.2000 24.9000 152.8000 ;
	    RECT 68.6000 148.2000 68.9000 152.8000 ;
	    RECT 24.6000 147.8000 25.0000 148.2000 ;
	    RECT 30.2000 148.1000 30.6000 148.2000 ;
	    RECT 31.0000 148.1000 31.4000 148.2000 ;
	    RECT 30.2000 147.8000 31.4000 148.1000 ;
	    RECT 68.6000 147.8000 69.0000 148.2000 ;
	    RECT 70.2000 148.1000 70.6000 148.2000 ;
	    RECT 71.0000 148.1000 71.4000 148.2000 ;
	    RECT 70.2000 147.8000 71.4000 148.1000 ;
         LAYER metal3 ;
	    RECT 24.6000 157.1000 25.0000 157.2000 ;
	    RECT 68.6000 157.1000 69.0000 157.2000 ;
	    RECT 72.6000 157.1000 73.0000 157.2000 ;
	    RECT 24.6000 156.8000 73.0000 157.1000 ;
	    RECT 24.6000 148.1000 25.0000 148.2000 ;
	    RECT 30.2000 148.1000 30.6000 148.2000 ;
	    RECT 24.6000 147.8000 30.6000 148.1000 ;
	    RECT 68.6000 148.1000 69.0000 148.2000 ;
	    RECT 70.2000 148.1000 70.6000 148.2000 ;
	    RECT 68.6000 147.8000 70.6000 148.1000 ;
      END
   END DATA_A[20]
   PIN DATA_A[19]
      PORT
         LAYER metal1 ;
	    RECT 3.0000 92.4000 3.4000 93.2000 ;
	    RECT 39.0000 92.4000 39.4000 93.2000 ;
	    RECT 25.4000 72.4000 25.8000 73.2000 ;
	    RECT 41.4000 72.4000 41.8000 73.2000 ;
         LAYER metal2 ;
	    RECT 3.0000 92.8000 3.4000 93.2000 ;
	    RECT 39.0000 92.8000 39.4000 93.2000 ;
	    RECT 3.0000 92.2000 3.3000 92.8000 ;
	    RECT 3.0000 91.8000 3.4000 92.2000 ;
	    RECT 39.0000 85.2000 39.3000 92.8000 ;
	    RECT 39.0000 84.8000 39.4000 85.2000 ;
	    RECT 41.4000 84.8000 41.8000 85.2000 ;
	    RECT 41.4000 77.2000 41.7000 84.8000 ;
	    RECT 25.4000 76.8000 25.8000 77.2000 ;
	    RECT 41.4000 76.8000 41.8000 77.2000 ;
	    RECT 25.4000 73.2000 25.7000 76.8000 ;
	    RECT 41.4000 73.2000 41.7000 76.8000 ;
	    RECT 25.4000 72.8000 25.8000 73.2000 ;
	    RECT 41.4000 72.8000 41.8000 73.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 97.1000 -2.2000 97.2000 ;
	    RECT 0.6000 97.1000 1.0000 97.2000 ;
	    RECT -2.6000 96.8000 1.0000 97.1000 ;
	    RECT 0.6000 93.1000 1.0000 93.2000 ;
	    RECT 7.0000 93.1000 7.4000 93.2000 ;
	    RECT 0.6000 92.8000 7.4000 93.1000 ;
	    RECT 3.0000 92.2000 3.3000 92.8000 ;
	    RECT 3.0000 91.8000 3.4000 92.2000 ;
	    RECT 39.0000 85.1000 39.4000 85.2000 ;
	    RECT 41.4000 85.1000 41.8000 85.2000 ;
	    RECT 39.0000 84.8000 41.8000 85.1000 ;
	    RECT 7.0000 77.1000 7.4000 77.2000 ;
	    RECT 25.4000 77.1000 25.8000 77.2000 ;
	    RECT 41.4000 77.1000 41.8000 77.2000 ;
	    RECT 7.0000 76.8000 41.8000 77.1000 ;
         LAYER metal4 ;
	    RECT 0.6000 96.8000 1.0000 97.2000 ;
	    RECT 0.6000 93.2000 0.9000 96.8000 ;
	    RECT 0.6000 92.8000 1.0000 93.2000 ;
	    RECT 7.0000 92.8000 7.4000 93.2000 ;
	    RECT 7.0000 77.2000 7.3000 92.8000 ;
	    RECT 7.0000 76.8000 7.4000 77.2000 ;
      END
   END DATA_A[19]
   PIN DATA_A[18]
      PORT
         LAYER metal1 ;
	    RECT 19.0000 92.4000 19.4000 93.2000 ;
	    RECT 62.2000 92.4000 62.6000 93.2000 ;
	    RECT 0.6000 87.8000 1.0000 88.6000 ;
	    RECT 62.2000 87.8000 62.6000 88.6000 ;
         LAYER metal2 ;
	    RECT 19.0000 92.8000 19.4000 93.2000 ;
	    RECT 62.2000 92.8000 62.6000 93.2000 ;
	    RECT 19.0000 92.2000 19.3000 92.8000 ;
	    RECT 62.2000 92.2000 62.5000 92.8000 ;
	    RECT 19.0000 91.8000 19.4000 92.2000 ;
	    RECT 62.2000 91.8000 62.6000 92.2000 ;
	    RECT 19.0000 90.2000 19.3000 91.8000 ;
	    RECT 0.6000 89.8000 1.0000 90.2000 ;
	    RECT 19.0000 89.8000 19.4000 90.2000 ;
	    RECT 0.6000 88.2000 0.9000 89.8000 ;
	    RECT 62.2000 88.2000 62.5000 91.8000 ;
	    RECT 0.6000 87.8000 1.0000 88.2000 ;
	    RECT 62.2000 87.8000 62.6000 88.2000 ;
         LAYER metal3 ;
	    RECT 19.0000 92.1000 19.4000 92.2000 ;
	    RECT 62.2000 92.1000 62.6000 92.2000 ;
	    RECT 19.0000 91.8000 62.6000 92.1000 ;
	    RECT -2.6000 90.1000 -2.2000 90.2000 ;
	    RECT 0.6000 90.1000 1.0000 90.2000 ;
	    RECT 19.0000 90.1000 19.4000 90.2000 ;
	    RECT -2.6000 89.8000 19.4000 90.1000 ;
      END
   END DATA_A[18]
   PIN DATA_A[17]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 112.4000 21.0000 113.2000 ;
	    RECT 79.8000 92.4000 80.2000 93.2000 ;
	    RECT 36.6000 67.8000 37.0000 68.6000 ;
	    RECT 62.2000 67.8000 62.6000 68.6000 ;
         LAYER metal2 ;
	    RECT 20.6000 113.1000 21.0000 113.2000 ;
	    RECT 21.4000 113.1000 21.8000 113.2000 ;
	    RECT 20.6000 112.8000 21.8000 113.1000 ;
	    RECT 20.6000 109.2000 20.9000 112.8000 ;
	    RECT 1.4000 108.8000 1.8000 109.2000 ;
	    RECT 20.6000 108.8000 21.0000 109.2000 ;
	    RECT 1.4000 106.2000 1.7000 108.8000 ;
	    RECT 1.4000 105.8000 1.8000 106.2000 ;
	    RECT 79.8000 92.8000 80.2000 93.2000 ;
	    RECT 79.8000 90.2000 80.1000 92.8000 ;
	    RECT 79.8000 89.8000 80.2000 90.2000 ;
	    RECT 36.6000 71.8000 37.0000 72.2000 ;
	    RECT 36.6000 68.2000 36.9000 71.8000 ;
	    RECT 62.2000 68.8000 62.6000 69.2000 ;
	    RECT 62.2000 68.2000 62.5000 68.8000 ;
	    RECT 36.6000 67.8000 37.0000 68.2000 ;
	    RECT 62.2000 67.8000 62.6000 68.2000 ;
         LAYER metal3 ;
	    RECT 21.4000 113.1000 21.8000 113.2000 ;
	    RECT 28.6000 113.1000 29.0000 113.2000 ;
	    RECT 21.4000 112.8000 29.0000 113.1000 ;
	    RECT 1.4000 109.1000 1.8000 109.2000 ;
	    RECT 20.6000 109.1000 21.0000 109.2000 ;
	    RECT 1.4000 108.8000 21.0000 109.1000 ;
	    RECT -2.6000 106.1000 -2.2000 106.2000 ;
	    RECT 1.4000 106.1000 1.8000 106.2000 ;
	    RECT -2.6000 105.8000 1.8000 106.1000 ;
	    RECT 68.6000 90.1000 69.0000 90.2000 ;
	    RECT 79.8000 90.1000 80.2000 90.2000 ;
	    RECT 68.6000 89.8000 80.2000 90.1000 ;
	    RECT 28.6000 72.1000 29.0000 72.2000 ;
	    RECT 36.6000 72.1000 37.0000 72.2000 ;
	    RECT 54.2000 72.1000 54.6000 72.2000 ;
	    RECT 28.6000 71.8000 54.6000 72.1000 ;
	    RECT 54.2000 69.1000 54.6000 69.2000 ;
	    RECT 62.2000 69.1000 62.6000 69.2000 ;
	    RECT 68.6000 69.1000 69.0000 69.2000 ;
	    RECT 54.2000 68.8000 69.0000 69.1000 ;
         LAYER metal4 ;
	    RECT 28.6000 112.8000 29.0000 113.2000 ;
	    RECT 28.6000 72.2000 28.9000 112.8000 ;
	    RECT 68.6000 89.8000 69.0000 90.2000 ;
	    RECT 28.6000 71.8000 29.0000 72.2000 ;
	    RECT 54.2000 71.8000 54.6000 72.2000 ;
	    RECT 54.2000 69.2000 54.5000 71.8000 ;
	    RECT 68.6000 69.2000 68.9000 89.8000 ;
	    RECT 54.2000 68.8000 54.6000 69.2000 ;
	    RECT 68.6000 68.8000 69.0000 69.2000 ;
      END
   END DATA_A[17]
   PIN DATA_A[16]
      PORT
         LAYER metal1 ;
	    RECT 7.0000 113.1000 7.4000 113.2000 ;
	    RECT 7.8000 113.1000 8.2000 113.2000 ;
	    RECT 7.0000 112.8000 8.2000 113.1000 ;
	    RECT 7.0000 112.4000 7.4000 112.8000 ;
	    RECT 7.8000 112.4000 8.2000 112.8000 ;
	    RECT 31.0000 112.4000 31.4000 113.2000 ;
	    RECT 32.6000 112.4000 33.0000 113.2000 ;
         LAYER metal2 ;
	    RECT 7.0000 113.8000 7.4000 114.2000 ;
	    RECT 31.0000 113.8000 31.4000 114.2000 ;
	    RECT 32.6000 113.8000 33.0000 114.2000 ;
	    RECT 7.0000 113.2000 7.3000 113.8000 ;
	    RECT 31.0000 113.2000 31.3000 113.8000 ;
	    RECT 32.6000 113.2000 32.9000 113.8000 ;
	    RECT 7.0000 112.8000 7.4000 113.2000 ;
	    RECT 31.0000 112.8000 31.4000 113.2000 ;
	    RECT 32.6000 112.8000 33.0000 113.2000 ;
         LAYER metal3 ;
	    RECT 7.0000 114.1000 7.4000 114.2000 ;
	    RECT 31.0000 114.1000 31.4000 114.2000 ;
	    RECT 32.6000 114.1000 33.0000 114.2000 ;
	    RECT -2.6000 113.8000 33.0000 114.1000 ;
	    RECT -2.6000 113.2000 -2.3000 113.8000 ;
	    RECT -2.6000 112.8000 -2.2000 113.2000 ;
      END
   END DATA_A[16]
   PIN DATA_A[15]
      PORT
         LAYER metal1 ;
	    RECT 35.8000 72.4000 36.2000 73.2000 ;
	    RECT 42.2000 67.8000 42.6000 68.6000 ;
	    RECT 49.4000 67.8000 49.8000 68.6000 ;
	    RECT 9.4000 52.4000 9.8000 53.2000 ;
         LAYER metal2 ;
	    RECT 35.8000 72.8000 36.2000 73.2000 ;
	    RECT 35.8000 69.2000 36.1000 72.8000 ;
	    RECT 35.8000 68.8000 36.2000 69.2000 ;
	    RECT 42.2000 68.8000 42.6000 69.2000 ;
	    RECT 49.4000 68.8000 49.8000 69.2000 ;
	    RECT 42.2000 68.2000 42.5000 68.8000 ;
	    RECT 49.4000 68.2000 49.7000 68.8000 ;
	    RECT 42.2000 67.8000 42.6000 68.2000 ;
	    RECT 49.4000 67.8000 49.8000 68.2000 ;
	    RECT 8.6000 53.1000 9.0000 53.2000 ;
	    RECT 9.4000 53.1000 9.8000 53.2000 ;
	    RECT 8.6000 52.8000 9.8000 53.1000 ;
         LAYER metal3 ;
	    RECT 14.2000 69.1000 14.6000 69.2000 ;
	    RECT 35.8000 69.1000 36.2000 69.2000 ;
	    RECT 42.2000 69.1000 42.6000 69.2000 ;
	    RECT 49.4000 69.1000 49.8000 69.2000 ;
	    RECT 14.2000 68.8000 49.8000 69.1000 ;
	    RECT -2.6000 53.8000 -2.2000 54.2000 ;
	    RECT -2.6000 53.1000 -2.3000 53.8000 ;
	    RECT 8.6000 53.1000 9.0000 53.2000 ;
	    RECT 14.2000 53.1000 14.6000 53.2000 ;
	    RECT -2.6000 52.8000 14.6000 53.1000 ;
         LAYER metal4 ;
	    RECT 14.2000 68.8000 14.6000 69.2000 ;
	    RECT 14.2000 53.2000 14.5000 68.8000 ;
	    RECT 14.2000 52.8000 14.6000 53.2000 ;
      END
   END DATA_A[15]
   PIN DATA_A[14]
      PORT
         LAYER metal1 ;
	    RECT 31.0000 153.8000 31.4000 154.2000 ;
	    RECT 31.0000 153.2000 31.3000 153.8000 ;
	    RECT 7.8000 152.4000 8.2000 153.2000 ;
	    RECT 27.8000 152.4000 28.2000 153.2000 ;
	    RECT 31.0000 152.4000 31.4000 153.2000 ;
	    RECT 11.0000 147.8000 11.4000 148.6000 ;
         LAYER metal2 ;
	    RECT 31.0000 153.8000 31.4000 154.2000 ;
	    RECT 31.0000 153.2000 31.3000 153.8000 ;
	    RECT 7.8000 153.1000 8.2000 153.2000 ;
	    RECT 8.6000 153.1000 9.0000 153.2000 ;
	    RECT 7.8000 152.8000 9.0000 153.1000 ;
	    RECT 11.0000 152.8000 11.4000 153.2000 ;
	    RECT 27.8000 153.1000 28.2000 153.2000 ;
	    RECT 28.6000 153.1000 29.0000 153.2000 ;
	    RECT 27.8000 152.8000 29.0000 153.1000 ;
	    RECT 31.0000 152.8000 31.4000 153.2000 ;
	    RECT 11.0000 148.2000 11.3000 152.8000 ;
	    RECT 11.0000 147.8000 11.4000 148.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 153.1000 -2.2000 153.2000 ;
	    RECT 8.6000 153.1000 9.0000 153.2000 ;
	    RECT 11.0000 153.1000 11.4000 153.2000 ;
	    RECT 28.6000 153.1000 29.0000 153.2000 ;
	    RECT 31.0000 153.1000 31.4000 153.2000 ;
	    RECT -2.6000 152.8000 31.4000 153.1000 ;
      END
   END DATA_A[14]
   PIN DATA_A[13]
      PORT
         LAYER metal1 ;
	    RECT 30.2000 152.4000 30.6000 153.2000 ;
	    RECT 42.2000 147.8000 42.6000 148.6000 ;
	    RECT 38.2000 132.4000 38.6000 133.2000 ;
	    RECT 45.4000 132.4000 45.8000 133.2000 ;
         LAYER metal2 ;
	    RECT 29.4000 163.8000 29.8000 164.2000 ;
	    RECT 29.4000 163.1000 29.7000 163.8000 ;
	    RECT 29.4000 162.8000 30.5000 163.1000 ;
	    RECT 30.2000 153.2000 30.5000 162.8000 ;
	    RECT 30.2000 152.8000 30.6000 153.2000 ;
	    RECT 30.2000 151.2000 30.5000 152.8000 ;
	    RECT 30.2000 150.8000 30.6000 151.2000 ;
	    RECT 42.2000 150.8000 42.6000 151.2000 ;
	    RECT 45.4000 150.8000 45.8000 151.2000 ;
	    RECT 42.2000 148.2000 42.5000 150.8000 ;
	    RECT 42.2000 147.8000 42.6000 148.2000 ;
	    RECT 45.4000 133.2000 45.7000 150.8000 ;
	    RECT 38.2000 133.1000 38.6000 133.2000 ;
	    RECT 39.0000 133.1000 39.4000 133.2000 ;
	    RECT 38.2000 132.8000 39.4000 133.1000 ;
	    RECT 45.4000 132.8000 45.8000 133.2000 ;
         LAYER metal3 ;
	    RECT 30.2000 151.1000 30.6000 151.2000 ;
	    RECT 42.2000 151.1000 42.6000 151.2000 ;
	    RECT 45.4000 151.1000 45.8000 151.2000 ;
	    RECT 30.2000 150.8000 45.8000 151.1000 ;
	    RECT 39.0000 133.1000 39.4000 133.2000 ;
	    RECT 45.4000 133.1000 45.8000 133.2000 ;
	    RECT 39.0000 132.8000 45.8000 133.1000 ;
      END
   END DATA_A[13]
   PIN DATA_A[12]
      PORT
         LAYER metal1 ;
	    RECT 56.6000 152.4000 57.0000 153.2000 ;
	    RECT 19.8000 147.8000 20.2000 148.6000 ;
	    RECT 35.8000 147.8000 36.2000 148.6000 ;
	    RECT 55.0000 147.8000 55.4000 148.6000 ;
         LAYER metal2 ;
	    RECT 56.6000 163.8000 57.0000 164.2000 ;
	    RECT 56.6000 153.2000 56.9000 163.8000 ;
	    RECT 56.6000 152.8000 57.0000 153.2000 ;
	    RECT 56.6000 150.2000 56.9000 152.8000 ;
	    RECT 55.0000 149.8000 55.4000 150.2000 ;
	    RECT 56.6000 149.8000 57.0000 150.2000 ;
	    RECT 19.8000 148.8000 20.2000 149.2000 ;
	    RECT 35.8000 148.8000 36.2000 149.2000 ;
	    RECT 19.8000 148.2000 20.1000 148.8000 ;
	    RECT 35.8000 148.2000 36.1000 148.8000 ;
	    RECT 55.0000 148.2000 55.3000 149.8000 ;
	    RECT 19.8000 147.8000 20.2000 148.2000 ;
	    RECT 35.8000 147.8000 36.2000 148.2000 ;
	    RECT 55.0000 147.8000 55.4000 148.2000 ;
         LAYER metal3 ;
	    RECT 55.0000 150.1000 55.4000 150.2000 ;
	    RECT 56.6000 150.1000 57.0000 150.2000 ;
	    RECT 35.8000 149.8000 57.0000 150.1000 ;
	    RECT 35.8000 149.2000 36.1000 149.8000 ;
	    RECT 19.8000 149.1000 20.2000 149.2000 ;
	    RECT 35.8000 149.1000 36.2000 149.2000 ;
	    RECT 19.8000 148.8000 36.2000 149.1000 ;
      END
   END DATA_A[12]
   PIN DATA_A[11]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 86.8000 21.1000 87.2000 ;
	    RECT 83.8000 87.1000 84.2000 87.2000 ;
	    RECT 84.6000 87.1000 85.1000 87.2000 ;
	    RECT 83.8000 86.8000 85.1000 87.1000 ;
	    RECT 20.8000 86.4000 21.2000 86.8000 ;
	    RECT 84.8000 86.4000 85.2000 86.8000 ;
	    RECT 16.0000 74.2000 16.4000 74.6000 ;
	    RECT 75.6000 74.2000 76.0000 74.6000 ;
	    RECT 15.8000 73.8000 16.3000 74.2000 ;
	    RECT 75.7000 73.8000 76.2000 74.2000 ;
         LAYER metal2 ;
	    RECT 20.6000 86.8000 21.0000 87.2000 ;
	    RECT 83.8000 86.8000 84.2000 87.2000 ;
	    RECT 20.6000 82.2000 20.9000 86.8000 ;
	    RECT 15.8000 81.8000 16.2000 82.2000 ;
	    RECT 20.6000 81.8000 21.0000 82.2000 ;
	    RECT 15.8000 76.2000 16.1000 81.8000 ;
	    RECT 20.6000 78.2000 20.9000 81.8000 ;
	    RECT 83.8000 78.2000 84.1000 86.8000 ;
	    RECT 20.6000 77.8000 21.0000 78.2000 ;
	    RECT 75.8000 77.8000 76.2000 78.2000 ;
	    RECT 83.8000 77.8000 84.2000 78.2000 ;
	    RECT 15.8000 75.8000 16.2000 76.2000 ;
	    RECT 15.8000 74.2000 16.1000 75.8000 ;
	    RECT 75.8000 74.2000 76.1000 77.8000 ;
	    RECT 15.8000 73.8000 16.2000 74.2000 ;
	    RECT 75.8000 73.8000 76.2000 74.2000 ;
         LAYER metal3 ;
	    RECT 15.8000 82.1000 16.2000 82.2000 ;
	    RECT 20.6000 82.1000 21.0000 82.2000 ;
	    RECT 15.8000 81.8000 21.0000 82.1000 ;
	    RECT 20.6000 78.1000 21.0000 78.2000 ;
	    RECT 75.8000 78.1000 76.2000 78.2000 ;
	    RECT 83.8000 78.1000 84.2000 78.2000 ;
	    RECT 20.6000 77.8000 84.2000 78.1000 ;
	    RECT 5.4000 76.1000 5.8000 76.2000 ;
	    RECT 15.8000 76.1000 16.2000 76.2000 ;
	    RECT 5.4000 75.8000 16.2000 76.1000 ;
	    RECT -2.6000 74.1000 -2.2000 74.2000 ;
	    RECT 5.4000 74.1000 5.8000 74.2000 ;
	    RECT -2.6000 73.8000 5.8000 74.1000 ;
         LAYER metal4 ;
	    RECT 5.4000 75.8000 5.8000 76.2000 ;
	    RECT 5.4000 74.2000 5.7000 75.8000 ;
	    RECT 5.4000 73.8000 5.8000 74.2000 ;
      END
   END DATA_A[11]
   PIN DATA_A[10]
      PORT
         LAYER metal1 ;
	    RECT 25.6000 114.2000 26.0000 114.6000 ;
	    RECT 49.6000 114.2000 50.0000 114.6000 ;
	    RECT 25.4000 113.8000 25.9000 114.2000 ;
	    RECT 49.4000 113.8000 49.9000 114.2000 ;
	    RECT 52.8000 74.2000 53.2000 74.6000 ;
	    RECT 52.6000 73.8000 53.1000 74.2000 ;
	    RECT 5.3000 46.8000 5.8000 47.2000 ;
	    RECT 5.2000 46.4000 5.6000 46.8000 ;
         LAYER metal2 ;
	    RECT 25.4000 113.8000 25.8000 114.2000 ;
	    RECT 49.4000 114.1000 49.8000 114.2000 ;
	    RECT 50.2000 114.1000 50.6000 114.2000 ;
	    RECT 49.4000 113.8000 50.6000 114.1000 ;
	    RECT 25.4000 111.2000 25.7000 113.8000 ;
	    RECT 25.4000 110.8000 25.8000 111.2000 ;
	    RECT 52.6000 92.8000 53.0000 93.2000 ;
	    RECT 52.6000 74.2000 52.9000 92.8000 ;
	    RECT 52.6000 73.8000 53.0000 74.2000 ;
	    RECT 5.4000 50.8000 5.8000 51.2000 ;
	    RECT 5.4000 47.2000 5.7000 50.8000 ;
	    RECT 5.4000 46.8000 5.8000 47.2000 ;
         LAYER metal3 ;
	    RECT 49.4000 114.1000 49.8000 114.2000 ;
	    RECT 50.2000 114.1000 50.6000 114.2000 ;
	    RECT 49.4000 113.8000 50.6000 114.1000 ;
	    RECT 25.4000 111.1000 25.8000 111.2000 ;
	    RECT 26.2000 111.1000 26.6000 111.2000 ;
	    RECT 25.4000 110.8000 26.6000 111.1000 ;
	    RECT 49.4000 93.1000 49.8000 93.2000 ;
	    RECT 52.6000 93.1000 53.0000 93.2000 ;
	    RECT 49.4000 92.8000 53.0000 93.1000 ;
	    RECT -2.6000 51.1000 -2.2000 51.2000 ;
	    RECT 5.4000 51.1000 5.8000 51.2000 ;
	    RECT 6.2000 51.1000 6.6000 51.2000 ;
	    RECT -2.6000 50.8000 6.6000 51.1000 ;
         LAYER metal4 ;
	    RECT 49.4000 113.8000 49.8000 114.2000 ;
	    RECT 49.4000 111.2000 49.7000 113.8000 ;
	    RECT 6.2000 110.8000 6.6000 111.2000 ;
	    RECT 25.4000 111.1000 25.8000 111.2000 ;
	    RECT 26.2000 111.1000 26.6000 111.2000 ;
	    RECT 25.4000 110.8000 26.6000 111.1000 ;
	    RECT 49.4000 110.8000 49.8000 111.2000 ;
	    RECT 6.2000 51.2000 6.5000 110.8000 ;
	    RECT 49.4000 93.2000 49.7000 110.8000 ;
	    RECT 49.4000 92.8000 49.8000 93.2000 ;
	    RECT 6.2000 50.8000 6.6000 51.2000 ;
         LAYER metal5 ;
	    RECT 6.2000 111.1000 6.6000 111.2000 ;
	    RECT 25.4000 111.1000 25.8000 111.2000 ;
	    RECT 49.4000 111.1000 49.8000 111.2000 ;
	    RECT 6.2000 110.8000 49.8000 111.1000 ;
      END
   END DATA_A[10]
   PIN DATA_A[9]
      PORT
         LAYER metal1 ;
	    RECT 34.0000 94.2000 34.4000 94.6000 ;
	    RECT 94.4000 94.2000 94.8000 94.6000 ;
	    RECT 34.1000 93.8000 34.6000 94.2000 ;
	    RECT 94.2000 93.8000 94.7000 94.2000 ;
	    RECT 78.4000 74.2000 78.8000 74.6000 ;
	    RECT 77.4000 74.1000 77.8000 74.2000 ;
	    RECT 78.2000 74.1000 78.7000 74.2000 ;
	    RECT 77.4000 73.8000 78.7000 74.1000 ;
	    RECT 30.8000 54.2000 31.2000 54.6000 ;
	    RECT 30.9000 53.8000 31.4000 54.2000 ;
         LAYER metal2 ;
	    RECT 33.4000 94.1000 33.8000 94.2000 ;
	    RECT 34.2000 94.1000 34.6000 94.2000 ;
	    RECT 33.4000 93.8000 34.6000 94.1000 ;
	    RECT 94.2000 93.8000 94.6000 94.2000 ;
	    RECT 94.2000 89.2000 94.5000 93.8000 ;
	    RECT 77.4000 88.8000 77.8000 89.2000 ;
	    RECT 94.2000 88.8000 94.6000 89.2000 ;
	    RECT 77.4000 74.2000 77.7000 88.8000 ;
	    RECT 77.4000 73.8000 77.8000 74.2000 ;
	    RECT 77.4000 73.2000 77.7000 73.8000 ;
	    RECT 77.4000 72.8000 77.8000 73.2000 ;
	    RECT 31.0000 61.8000 31.4000 62.2000 ;
	    RECT 31.0000 54.2000 31.3000 61.8000 ;
	    RECT 31.0000 53.8000 31.4000 54.2000 ;
         LAYER metal3 ;
	    RECT 32.6000 94.1000 33.0000 94.2000 ;
	    RECT 33.4000 94.1000 33.8000 94.2000 ;
	    RECT 32.6000 93.8000 33.8000 94.1000 ;
	    RECT 77.4000 89.1000 77.8000 89.2000 ;
	    RECT 94.2000 89.1000 94.6000 89.2000 ;
	    RECT 77.4000 88.8000 94.6000 89.1000 ;
	    RECT 74.2000 73.1000 74.6000 73.2000 ;
	    RECT 77.4000 73.1000 77.8000 73.2000 ;
	    RECT 74.2000 72.8000 77.8000 73.1000 ;
	    RECT 4.6000 62.1000 5.0000 62.2000 ;
	    RECT 31.0000 62.1000 31.4000 62.2000 ;
	    RECT 33.4000 62.1000 33.8000 62.2000 ;
	    RECT 4.6000 61.8000 33.8000 62.1000 ;
	    RECT -2.6000 60.1000 -2.2000 60.2000 ;
	    RECT 4.6000 60.1000 5.0000 60.2000 ;
	    RECT -2.6000 59.8000 5.0000 60.1000 ;
         LAYER metal4 ;
	    RECT 32.6000 94.1000 33.0000 94.2000 ;
	    RECT 32.6000 93.8000 33.7000 94.1000 ;
	    RECT 33.4000 73.2000 33.7000 93.8000 ;
	    RECT 33.4000 72.8000 33.8000 73.2000 ;
	    RECT 73.4000 73.1000 73.8000 73.2000 ;
	    RECT 74.2000 73.1000 74.6000 73.2000 ;
	    RECT 73.4000 72.8000 74.6000 73.1000 ;
	    RECT 33.4000 62.2000 33.7000 72.8000 ;
	    RECT 4.6000 61.8000 5.0000 62.2000 ;
	    RECT 33.4000 61.8000 33.8000 62.2000 ;
	    RECT 4.6000 60.2000 4.9000 61.8000 ;
	    RECT 4.6000 59.8000 5.0000 60.2000 ;
         LAYER metal5 ;
	    RECT 33.4000 73.1000 33.8000 73.2000 ;
	    RECT 73.4000 73.1000 73.8000 73.2000 ;
	    RECT 33.4000 72.8000 73.8000 73.1000 ;
      END
   END DATA_A[9]
   PIN DATA_A[8]
      PORT
         LAYER metal1 ;
	    RECT 12.5000 106.8000 13.0000 107.2000 ;
	    RECT 41.4000 107.1000 41.8000 107.2000 ;
	    RECT 42.2000 107.1000 42.7000 107.2000 ;
	    RECT 41.4000 106.8000 42.7000 107.1000 ;
	    RECT 12.4000 106.4000 12.8000 106.8000 ;
	    RECT 42.4000 106.4000 42.8000 106.8000 ;
	    RECT 68.0000 94.2000 68.4000 94.6000 ;
	    RECT 67.8000 93.8000 68.3000 94.2000 ;
	    RECT 6.2000 87.1000 6.6000 87.2000 ;
	    RECT 7.0000 87.1000 7.5000 87.2000 ;
	    RECT 6.2000 86.8000 7.5000 87.1000 ;
	    RECT 7.2000 86.4000 7.6000 86.8000 ;
         LAYER metal2 ;
	    RECT 12.6000 106.8000 13.0000 107.2000 ;
	    RECT 41.4000 106.8000 41.8000 107.2000 ;
	    RECT 12.6000 100.2000 12.9000 106.8000 ;
	    RECT 41.4000 100.2000 41.7000 106.8000 ;
	    RECT 12.6000 99.8000 13.0000 100.2000 ;
	    RECT 41.4000 99.8000 41.8000 100.2000 ;
	    RECT 41.4000 98.2000 41.7000 99.8000 ;
	    RECT 41.4000 97.8000 41.8000 98.2000 ;
	    RECT 67.8000 97.8000 68.2000 98.2000 ;
	    RECT 67.8000 94.2000 68.1000 97.8000 ;
	    RECT 67.8000 93.8000 68.2000 94.2000 ;
	    RECT 5.4000 87.1000 5.8000 87.2000 ;
	    RECT 6.2000 87.1000 6.6000 87.2000 ;
	    RECT 5.4000 86.8000 6.6000 87.1000 ;
         LAYER metal3 ;
	    RECT 7.8000 100.1000 8.2000 100.2000 ;
	    RECT 12.6000 100.1000 13.0000 100.2000 ;
	    RECT 41.4000 100.1000 41.8000 100.2000 ;
	    RECT 7.8000 99.8000 41.8000 100.1000 ;
	    RECT 41.4000 98.1000 41.8000 98.2000 ;
	    RECT 67.8000 98.1000 68.2000 98.2000 ;
	    RECT 41.4000 97.8000 68.2000 98.1000 ;
	    RECT -2.6000 87.8000 -2.2000 88.2000 ;
	    RECT -2.6000 87.1000 -2.3000 87.8000 ;
	    RECT 5.4000 87.1000 5.8000 87.2000 ;
	    RECT 7.8000 87.1000 8.2000 87.2000 ;
	    RECT -2.6000 86.8000 8.2000 87.1000 ;
         LAYER metal4 ;
	    RECT 7.8000 99.8000 8.2000 100.2000 ;
	    RECT 7.8000 87.2000 8.1000 99.8000 ;
	    RECT 7.8000 86.8000 8.2000 87.2000 ;
      END
   END DATA_A[8]
   PIN DATA_A[7]
      PORT
         LAYER metal1 ;
	    RECT 54.4000 94.2000 54.8000 94.6000 ;
	    RECT 54.2000 93.8000 54.7000 94.2000 ;
	    RECT 36.5000 86.8000 37.0000 87.2000 ;
	    RECT 51.8000 86.8000 52.3000 87.2000 ;
	    RECT 36.4000 86.4000 36.8000 86.8000 ;
	    RECT 52.0000 86.4000 52.4000 86.8000 ;
	    RECT 6.2000 66.8000 6.7000 67.2000 ;
	    RECT 6.4000 66.4000 6.8000 66.8000 ;
         LAYER metal2 ;
	    RECT 54.2000 93.8000 54.6000 94.2000 ;
	    RECT 36.6000 86.8000 37.0000 87.2000 ;
	    RECT 51.8000 86.8000 52.2000 87.2000 ;
	    RECT 36.6000 83.2000 36.9000 86.8000 ;
	    RECT 51.8000 83.2000 52.1000 86.8000 ;
	    RECT 54.2000 83.2000 54.5000 93.8000 ;
	    RECT 36.6000 82.8000 37.0000 83.2000 ;
	    RECT 51.8000 82.8000 52.2000 83.2000 ;
	    RECT 54.2000 82.8000 54.6000 83.2000 ;
	    RECT 6.2000 69.8000 6.6000 70.2000 ;
	    RECT 6.2000 67.2000 6.5000 69.8000 ;
	    RECT 6.2000 66.8000 6.6000 67.2000 ;
         LAYER metal3 ;
	    RECT 19.0000 83.1000 19.4000 83.2000 ;
	    RECT 36.6000 83.1000 37.0000 83.2000 ;
	    RECT 51.8000 83.1000 52.2000 83.2000 ;
	    RECT 54.2000 83.1000 54.6000 83.2000 ;
	    RECT 19.0000 82.8000 54.6000 83.1000 ;
	    RECT -2.6000 70.1000 -2.2000 70.2000 ;
	    RECT 6.2000 70.1000 6.6000 70.2000 ;
	    RECT 19.0000 70.1000 19.4000 70.2000 ;
	    RECT -2.6000 69.8000 19.4000 70.1000 ;
         LAYER metal4 ;
	    RECT 19.0000 82.8000 19.4000 83.2000 ;
	    RECT 19.0000 70.2000 19.3000 82.8000 ;
	    RECT 19.0000 69.8000 19.4000 70.2000 ;
      END
   END DATA_A[7]
   PIN DATA_A[6]
      PORT
         LAYER metal1 ;
	    RECT 5.3000 146.8000 5.8000 147.2000 ;
	    RECT 47.8000 146.8000 48.3000 147.2000 ;
	    RECT 5.2000 146.4000 5.6000 146.8000 ;
	    RECT 48.0000 146.4000 48.4000 146.8000 ;
	    RECT 22.9000 126.8000 23.4000 127.2000 ;
	    RECT 51.0000 126.8000 51.5000 127.2000 ;
	    RECT 22.8000 126.4000 23.2000 126.8000 ;
	    RECT 51.2000 126.4000 51.6000 126.8000 ;
         LAYER metal2 ;
	    RECT 5.4000 147.8000 5.8000 148.2000 ;
	    RECT 5.4000 147.2000 5.7000 147.8000 ;
	    RECT 5.4000 146.8000 5.8000 147.2000 ;
	    RECT 47.8000 146.8000 48.2000 147.2000 ;
	    RECT 5.4000 143.2000 5.7000 146.8000 ;
	    RECT 5.4000 142.8000 5.8000 143.2000 ;
	    RECT 47.8000 139.2000 48.1000 146.8000 ;
	    RECT 47.8000 138.8000 48.2000 139.2000 ;
	    RECT 51.0000 138.8000 51.4000 139.2000 ;
	    RECT 51.0000 129.2000 51.3000 138.8000 ;
	    RECT 23.0000 128.8000 23.4000 129.2000 ;
	    RECT 51.0000 128.8000 51.4000 129.2000 ;
	    RECT 23.0000 127.2000 23.3000 128.8000 ;
	    RECT 51.0000 127.2000 51.3000 128.8000 ;
	    RECT 23.0000 126.8000 23.4000 127.2000 ;
	    RECT 51.0000 126.8000 51.4000 127.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 148.1000 -2.2000 148.2000 ;
	    RECT 5.4000 148.1000 5.8000 148.2000 ;
	    RECT -2.6000 147.8000 5.8000 148.1000 ;
	    RECT 5.4000 143.1000 5.8000 143.2000 ;
	    RECT 6.2000 143.1000 6.6000 143.2000 ;
	    RECT 5.4000 142.8000 6.6000 143.1000 ;
	    RECT 47.8000 139.1000 48.2000 139.2000 ;
	    RECT 51.0000 139.1000 51.4000 139.2000 ;
	    RECT 47.8000 138.8000 51.4000 139.1000 ;
	    RECT 6.2000 129.1000 6.6000 129.2000 ;
	    RECT 23.0000 129.1000 23.4000 129.2000 ;
	    RECT 51.0000 129.1000 51.4000 129.2000 ;
	    RECT 6.2000 128.8000 51.4000 129.1000 ;
         LAYER metal4 ;
	    RECT 6.2000 142.8000 6.6000 143.2000 ;
	    RECT 6.2000 129.2000 6.5000 142.8000 ;
	    RECT 6.2000 128.8000 6.6000 129.2000 ;
      END
   END DATA_A[6]
   PIN DATA_A[5]
      PORT
         LAYER metal1 ;
	    RECT 6.4000 134.2000 6.8000 134.6000 ;
	    RECT 33.6000 134.2000 34.0000 134.6000 ;
	    RECT 65.6000 134.2000 66.0000 134.6000 ;
	    RECT 73.6000 134.2000 74.0000 134.6000 ;
	    RECT 4.6000 134.1000 5.0000 134.2000 ;
	    RECT 6.2000 134.1000 6.7000 134.2000 ;
	    RECT 4.6000 133.8000 6.7000 134.1000 ;
	    RECT 33.4000 133.8000 33.9000 134.2000 ;
	    RECT 65.4000 133.8000 65.9000 134.2000 ;
	    RECT 73.4000 133.8000 73.9000 134.2000 ;
         LAYER metal2 ;
	    RECT 73.4000 135.8000 73.8000 136.2000 ;
	    RECT 4.6000 134.8000 5.0000 135.2000 ;
	    RECT 65.4000 134.8000 65.8000 135.2000 ;
	    RECT 4.6000 134.2000 4.9000 134.8000 ;
	    RECT 65.4000 134.2000 65.7000 134.8000 ;
	    RECT 73.4000 134.2000 73.7000 135.8000 ;
	    RECT 4.6000 133.8000 5.0000 134.2000 ;
	    RECT 32.6000 134.1000 33.0000 134.2000 ;
	    RECT 33.4000 134.1000 33.8000 134.2000 ;
	    RECT 32.6000 133.8000 33.8000 134.1000 ;
	    RECT 65.4000 133.8000 65.8000 134.2000 ;
	    RECT 73.4000 133.8000 73.8000 134.2000 ;
         LAYER metal3 ;
	    RECT 73.4000 136.1000 73.8000 136.2000 ;
	    RECT 65.4000 135.8000 73.8000 136.1000 ;
	    RECT 65.4000 135.2000 65.7000 135.8000 ;
	    RECT -2.6000 135.1000 -2.2000 135.2000 ;
	    RECT 4.6000 135.1000 5.0000 135.2000 ;
	    RECT -2.6000 134.8000 5.0000 135.1000 ;
	    RECT 64.6000 135.1000 65.0000 135.2000 ;
	    RECT 65.4000 135.1000 65.8000 135.2000 ;
	    RECT 64.6000 134.8000 65.8000 135.1000 ;
	    RECT 27.0000 134.1000 27.4000 134.2000 ;
	    RECT 32.6000 134.1000 33.0000 134.2000 ;
	    RECT 27.0000 133.8000 33.0000 134.1000 ;
         LAYER metal4 ;
	    RECT 4.6000 134.8000 5.0000 135.2000 ;
	    RECT 64.6000 135.1000 65.0000 135.2000 ;
	    RECT 64.6000 134.8000 65.7000 135.1000 ;
	    RECT 4.6000 134.2000 4.9000 134.8000 ;
	    RECT 65.4000 134.2000 65.7000 134.8000 ;
	    RECT 4.6000 133.8000 5.0000 134.2000 ;
	    RECT 26.2000 134.1000 26.6000 134.2000 ;
	    RECT 27.0000 134.1000 27.4000 134.2000 ;
	    RECT 26.2000 133.8000 27.4000 134.1000 ;
	    RECT 65.4000 133.8000 65.8000 134.2000 ;
         LAYER metal5 ;
	    RECT 4.6000 134.1000 5.0000 134.2000 ;
	    RECT 26.2000 134.1000 26.6000 134.2000 ;
	    RECT 65.4000 134.1000 65.8000 134.2000 ;
	    RECT 4.6000 133.8000 65.8000 134.1000 ;
      END
   END DATA_A[5]
   PIN DATA_A[4]
      PORT
         LAYER metal1 ;
	    RECT 25.3000 146.8000 25.8000 147.2000 ;
	    RECT 62.2000 146.8000 62.7000 147.2000 ;
	    RECT 25.2000 146.4000 25.6000 146.8000 ;
	    RECT 62.4000 146.4000 62.8000 146.8000 ;
	    RECT 25.4000 126.8000 25.9000 127.2000 ;
	    RECT 64.6000 126.8000 65.1000 127.2000 ;
	    RECT 25.6000 126.4000 26.0000 126.8000 ;
	    RECT 64.8000 126.4000 65.2000 126.8000 ;
         LAYER metal2 ;
	    RECT 63.0000 163.8000 63.4000 164.2000 ;
	    RECT 63.0000 161.2000 63.3000 163.8000 ;
	    RECT 63.0000 160.8000 63.4000 161.2000 ;
	    RECT 25.4000 146.8000 25.8000 147.2000 ;
	    RECT 62.2000 146.8000 62.6000 147.2000 ;
	    RECT 25.4000 144.2000 25.7000 146.8000 ;
	    RECT 62.2000 144.2000 62.5000 146.8000 ;
	    RECT 25.4000 143.8000 25.8000 144.2000 ;
	    RECT 62.2000 143.8000 62.6000 144.2000 ;
	    RECT 25.4000 133.1000 25.7000 143.8000 ;
	    RECT 25.4000 132.8000 26.5000 133.1000 ;
	    RECT 25.4000 127.1000 25.8000 127.2000 ;
	    RECT 26.2000 127.1000 26.5000 132.8000 ;
	    RECT 25.4000 126.8000 26.5000 127.1000 ;
	    RECT 64.6000 127.8000 65.0000 128.2000 ;
	    RECT 64.6000 127.2000 64.9000 127.8000 ;
	    RECT 64.6000 126.8000 65.0000 127.2000 ;
         LAYER metal3 ;
	    RECT 62.2000 161.1000 62.6000 161.2000 ;
	    RECT 63.0000 161.1000 63.4000 161.2000 ;
	    RECT 62.2000 160.8000 63.4000 161.1000 ;
	    RECT 25.4000 144.1000 25.8000 144.2000 ;
	    RECT 62.2000 144.1000 62.6000 144.2000 ;
	    RECT 63.0000 144.1000 63.4000 144.2000 ;
	    RECT 25.4000 143.8000 63.4000 144.1000 ;
	    RECT 63.0000 128.1000 63.4000 128.2000 ;
	    RECT 64.6000 128.1000 65.0000 128.2000 ;
	    RECT 63.0000 127.8000 65.0000 128.1000 ;
         LAYER metal4 ;
	    RECT 62.2000 161.1000 62.6000 161.2000 ;
	    RECT 62.2000 160.8000 63.3000 161.1000 ;
	    RECT 63.0000 144.2000 63.3000 160.8000 ;
	    RECT 63.0000 143.8000 63.4000 144.2000 ;
	    RECT 63.0000 128.2000 63.3000 143.8000 ;
	    RECT 63.0000 127.8000 63.4000 128.2000 ;
      END
   END DATA_A[4]
   PIN DATA_A[3]
      PORT
         LAYER metal1 ;
	    RECT 7.0000 92.4000 7.4000 93.2000 ;
	    RECT 43.0000 92.4000 43.4000 93.2000 ;
	    RECT 32.6000 72.4000 33.0000 73.2000 ;
	    RECT 45.4000 72.4000 45.8000 73.2000 ;
         LAYER metal2 ;
	    RECT 7.0000 92.8000 7.4000 93.2000 ;
	    RECT 43.0000 92.8000 43.4000 93.2000 ;
	    RECT 7.0000 81.2000 7.3000 92.8000 ;
	    RECT 7.0000 80.8000 7.4000 81.2000 ;
	    RECT 7.0000 80.2000 7.3000 80.8000 ;
	    RECT 7.0000 79.8000 7.4000 80.2000 ;
	    RECT 32.6000 79.8000 33.0000 80.2000 ;
	    RECT 32.6000 76.2000 32.9000 79.8000 ;
	    RECT 43.0000 76.2000 43.3000 92.8000 ;
	    RECT 32.6000 75.8000 33.0000 76.2000 ;
	    RECT 43.0000 75.8000 43.4000 76.2000 ;
	    RECT 45.4000 75.8000 45.8000 76.2000 ;
	    RECT 32.6000 73.2000 32.9000 75.8000 ;
	    RECT 45.4000 73.2000 45.7000 75.8000 ;
	    RECT 32.6000 72.8000 33.0000 73.2000 ;
	    RECT 45.4000 72.8000 45.8000 73.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 86.1000 -2.2000 86.2000 ;
	    RECT 1.4000 86.1000 1.8000 86.2000 ;
	    RECT -2.6000 85.8000 1.8000 86.1000 ;
	    RECT 1.4000 81.1000 1.8000 81.2000 ;
	    RECT 7.0000 81.1000 7.4000 81.2000 ;
	    RECT 1.4000 80.8000 7.4000 81.1000 ;
	    RECT 7.0000 80.1000 7.4000 80.2000 ;
	    RECT 32.6000 80.1000 33.0000 80.2000 ;
	    RECT 7.0000 79.8000 33.0000 80.1000 ;
	    RECT 32.6000 76.1000 33.0000 76.2000 ;
	    RECT 43.0000 76.1000 43.4000 76.2000 ;
	    RECT 45.4000 76.1000 45.8000 76.2000 ;
	    RECT 32.6000 75.8000 45.8000 76.1000 ;
         LAYER metal4 ;
	    RECT 1.4000 85.8000 1.8000 86.2000 ;
	    RECT 1.4000 81.2000 1.7000 85.8000 ;
	    RECT 1.4000 80.8000 1.8000 81.2000 ;
      END
   END DATA_A[3]
   PIN DATA_A[2]
      PORT
         LAYER metal1 ;
	    RECT 52.6000 106.8000 53.1000 107.2000 ;
	    RECT 52.8000 106.4000 53.2000 106.8000 ;
	    RECT 14.4000 94.2000 14.8000 94.6000 ;
	    RECT 14.2000 93.8000 14.7000 94.2000 ;
	    RECT 57.4000 87.1000 57.8000 87.2000 ;
	    RECT 58.2000 87.1000 58.7000 87.2000 ;
	    RECT 57.4000 86.8000 58.7000 87.1000 ;
	    RECT 58.4000 86.4000 58.8000 86.8000 ;
	    RECT 4.4000 74.2000 4.8000 74.6000 ;
	    RECT 4.5000 73.8000 5.0000 74.2000 ;
         LAYER metal2 ;
	    RECT 52.6000 106.8000 53.0000 107.2000 ;
	    RECT 52.6000 105.2000 52.9000 106.8000 ;
	    RECT 52.6000 104.8000 53.0000 105.2000 ;
	    RECT 14.2000 93.8000 14.6000 94.2000 ;
	    RECT 14.2000 91.2000 14.5000 93.8000 ;
	    RECT 14.2000 90.8000 14.6000 91.2000 ;
	    RECT 57.4000 87.1000 57.8000 87.2000 ;
	    RECT 58.2000 87.1000 58.6000 87.2000 ;
	    RECT 57.4000 86.8000 58.6000 87.1000 ;
	    RECT 4.6000 75.8000 5.0000 76.2000 ;
	    RECT 4.6000 74.2000 4.9000 75.8000 ;
	    RECT 4.6000 73.8000 5.0000 74.2000 ;
         LAYER metal3 ;
	    RECT 52.6000 105.1000 53.0000 105.2000 ;
	    RECT 54.2000 105.1000 54.6000 105.2000 ;
	    RECT 52.6000 104.8000 54.6000 105.1000 ;
	    RECT 0.6000 91.1000 1.0000 91.2000 ;
	    RECT 14.2000 91.1000 14.6000 91.2000 ;
	    RECT 54.2000 91.1000 54.6000 91.2000 ;
	    RECT 0.6000 90.8000 54.6000 91.1000 ;
	    RECT 54.2000 87.1000 54.6000 87.2000 ;
	    RECT 58.2000 87.1000 58.6000 87.2000 ;
	    RECT 54.2000 86.8000 58.6000 87.1000 ;
	    RECT -2.6000 76.1000 -2.2000 76.2000 ;
	    RECT 0.6000 76.1000 1.0000 76.2000 ;
	    RECT 4.6000 76.1000 5.0000 76.2000 ;
	    RECT -2.6000 75.8000 5.0000 76.1000 ;
         LAYER metal4 ;
	    RECT 54.2000 104.8000 54.6000 105.2000 ;
	    RECT 54.2000 91.2000 54.5000 104.8000 ;
	    RECT 0.6000 90.8000 1.0000 91.2000 ;
	    RECT 54.2000 90.8000 54.6000 91.2000 ;
	    RECT 0.6000 76.2000 0.9000 90.8000 ;
	    RECT 54.2000 87.2000 54.5000 90.8000 ;
	    RECT 54.2000 86.8000 54.6000 87.2000 ;
	    RECT 0.6000 75.8000 1.0000 76.2000 ;
      END
   END DATA_A[2]
   PIN DATA_A[1]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 106.8000 21.1000 107.2000 ;
	    RECT 20.8000 106.4000 21.2000 106.8000 ;
	    RECT 77.6000 94.2000 78.0000 94.6000 ;
	    RECT 77.4000 93.8000 77.9000 94.2000 ;
	    RECT 27.8000 66.8000 28.3000 67.2000 ;
	    RECT 71.7000 66.8000 72.2000 67.2000 ;
	    RECT 28.0000 66.4000 28.4000 66.8000 ;
	    RECT 71.6000 66.4000 72.0000 66.8000 ;
         LAYER metal2 ;
	    RECT 20.6000 107.1000 21.0000 107.2000 ;
	    RECT 21.4000 107.1000 21.8000 107.2000 ;
	    RECT 20.6000 106.8000 21.8000 107.1000 ;
	    RECT 77.4000 93.8000 77.8000 94.2000 ;
	    RECT 77.4000 92.2000 77.7000 93.8000 ;
	    RECT 71.0000 91.8000 71.4000 92.2000 ;
	    RECT 77.4000 91.8000 77.8000 92.2000 ;
	    RECT 27.8000 71.8000 28.2000 72.2000 ;
	    RECT 27.8000 68.2000 28.1000 71.8000 ;
	    RECT 27.8000 67.8000 28.2000 68.2000 ;
	    RECT 27.8000 67.2000 28.1000 67.8000 ;
	    RECT 71.0000 67.2000 71.3000 91.8000 ;
	    RECT 27.8000 66.8000 28.2000 67.2000 ;
	    RECT 71.0000 67.1000 71.4000 67.2000 ;
	    RECT 71.8000 67.1000 72.2000 67.2000 ;
	    RECT 71.0000 66.8000 72.2000 67.1000 ;
         LAYER metal3 ;
	    RECT -2.6000 108.1000 -2.2000 108.2000 ;
	    RECT -2.6000 107.8000 20.9000 108.1000 ;
	    RECT 20.6000 107.2000 20.9000 107.8000 ;
	    RECT 20.6000 107.1000 21.0000 107.2000 ;
	    RECT 21.4000 107.1000 21.8000 107.2000 ;
	    RECT 20.6000 106.8000 21.8000 107.1000 ;
	    RECT 71.0000 92.1000 71.4000 92.2000 ;
	    RECT 77.4000 92.1000 77.8000 92.2000 ;
	    RECT 71.0000 91.8000 77.8000 92.1000 ;
	    RECT 20.6000 72.1000 21.0000 72.2000 ;
	    RECT 27.8000 72.1000 28.2000 72.2000 ;
	    RECT 20.6000 71.8000 28.2000 72.1000 ;
	    RECT 27.8000 68.1000 28.2000 68.2000 ;
	    RECT 27.8000 67.8000 55.3000 68.1000 ;
	    RECT 55.0000 67.1000 55.3000 67.8000 ;
	    RECT 71.0000 67.1000 71.4000 67.2000 ;
	    RECT 55.0000 66.8000 71.4000 67.1000 ;
         LAYER metal4 ;
	    RECT 20.6000 106.8000 21.0000 107.2000 ;
	    RECT 20.6000 72.2000 20.9000 106.8000 ;
	    RECT 20.6000 71.8000 21.0000 72.2000 ;
      END
   END DATA_A[1]
   PIN DATA_A[0]
      PORT
         LAYER metal1 ;
	    RECT 44.6000 126.8000 45.1000 127.2000 ;
	    RECT 44.8000 126.4000 45.2000 126.8000 ;
	    RECT 1.6000 114.2000 2.0000 114.6000 ;
	    RECT 16.4000 114.2000 16.8000 114.6000 ;
	    RECT 43.2000 114.2000 43.6000 114.6000 ;
	    RECT 0.6000 114.1000 1.0000 114.2000 ;
	    RECT 1.4000 114.1000 1.9000 114.2000 ;
	    RECT 0.6000 113.8000 1.9000 114.1000 ;
	    RECT 16.5000 113.8000 17.0000 114.2000 ;
	    RECT 43.0000 113.8000 43.5000 114.2000 ;
         LAYER metal2 ;
	    RECT 44.6000 126.8000 45.0000 127.2000 ;
	    RECT 44.6000 116.2000 44.9000 126.8000 ;
	    RECT 43.0000 115.8000 43.4000 116.2000 ;
	    RECT 44.6000 115.8000 45.0000 116.2000 ;
	    RECT 0.6000 114.8000 1.0000 115.2000 ;
	    RECT 16.6000 114.8000 17.0000 115.2000 ;
	    RECT 0.6000 114.2000 0.9000 114.8000 ;
	    RECT 16.6000 114.2000 16.9000 114.8000 ;
	    RECT 43.0000 114.2000 43.3000 115.8000 ;
	    RECT 0.6000 113.8000 1.0000 114.2000 ;
	    RECT 16.6000 113.8000 17.0000 114.2000 ;
	    RECT 43.0000 113.8000 43.4000 114.2000 ;
         LAYER metal3 ;
	    RECT 43.0000 116.1000 43.4000 116.2000 ;
	    RECT 44.6000 116.1000 45.0000 116.2000 ;
	    RECT 31.8000 115.8000 45.0000 116.1000 ;
	    RECT -2.6000 115.1000 -2.2000 115.2000 ;
	    RECT 0.6000 115.1000 1.0000 115.2000 ;
	    RECT 16.6000 115.1000 17.0000 115.2000 ;
	    RECT 31.8000 115.1000 32.1000 115.8000 ;
	    RECT -2.6000 114.8000 32.1000 115.1000 ;
      END
   END DATA_A[0]
   PIN DATA_B[31]
      PORT
         LAYER metal1 ;
	    RECT 128.6000 52.4000 129.0000 53.2000 ;
	    RECT 166.2000 52.4000 166.6000 53.2000 ;
	    RECT 48.6000 47.8000 49.0000 48.6000 ;
	    RECT 79.8000 47.8000 80.2000 48.6000 ;
         LAYER metal2 ;
	    RECT 166.2000 60.8000 166.6000 61.2000 ;
	    RECT 166.2000 53.2000 166.5000 60.8000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 128.6000 53.1000 129.0000 53.2000 ;
	    RECT 127.8000 52.8000 129.0000 53.1000 ;
	    RECT 166.2000 52.8000 166.6000 53.2000 ;
	    RECT 48.6000 50.8000 49.0000 51.2000 ;
	    RECT 79.8000 50.8000 80.2000 51.2000 ;
	    RECT 48.6000 48.2000 48.9000 50.8000 ;
	    RECT 79.8000 48.2000 80.1000 50.8000 ;
	    RECT 128.6000 50.2000 128.9000 52.8000 ;
	    RECT 166.2000 50.2000 166.5000 52.8000 ;
	    RECT 128.6000 49.8000 129.0000 50.2000 ;
	    RECT 166.2000 49.8000 166.6000 50.2000 ;
	    RECT 48.6000 47.8000 49.0000 48.2000 ;
	    RECT 79.8000 47.8000 80.2000 48.2000 ;
         LAYER metal3 ;
	    RECT 166.2000 61.1000 166.6000 61.2000 ;
	    RECT 175.8000 61.1000 176.2000 61.2000 ;
	    RECT 166.2000 60.8000 176.2000 61.1000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 128.6000 53.1000 129.0000 53.2000 ;
	    RECT 127.8000 52.8000 129.0000 53.1000 ;
	    RECT 48.6000 51.1000 49.0000 51.2000 ;
	    RECT 79.8000 51.1000 80.2000 51.2000 ;
	    RECT 110.2000 51.1000 110.6000 51.2000 ;
	    RECT 48.6000 50.8000 110.6000 51.1000 ;
	    RECT 128.6000 50.1000 129.0000 50.2000 ;
	    RECT 166.2000 50.1000 166.6000 50.2000 ;
	    RECT 128.6000 49.8000 166.6000 50.1000 ;
         LAYER metal4 ;
	    RECT 110.2000 52.8000 110.6000 53.2000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 128.6000 53.1000 129.0000 53.2000 ;
	    RECT 127.8000 52.8000 129.0000 53.1000 ;
	    RECT 110.2000 51.2000 110.5000 52.8000 ;
	    RECT 110.2000 50.8000 110.6000 51.2000 ;
         LAYER metal5 ;
	    RECT 110.2000 53.1000 110.6000 53.2000 ;
	    RECT 127.8000 53.1000 128.2000 53.2000 ;
	    RECT 110.2000 52.8000 128.2000 53.1000 ;
      END
   END DATA_B[31]
   PIN DATA_B[30]
      PORT
         LAYER metal1 ;
	    RECT 4.6000 4.4000 5.0000 5.2000 ;
	    RECT 68.6000 4.4000 69.0000 5.2000 ;
	    RECT 95.0000 4.4000 95.4000 5.2000 ;
	    RECT 137.4000 4.1000 137.8000 4.2000 ;
	    RECT 138.2000 4.1000 138.6000 5.2000 ;
	    RECT 137.4000 3.8000 138.6000 4.1000 ;
         LAYER metal2 ;
	    RECT 4.6000 4.8000 5.0000 5.2000 ;
	    RECT 68.6000 4.8000 69.0000 5.2000 ;
	    RECT 95.0000 4.8000 95.4000 5.2000 ;
	    RECT 4.6000 1.2000 4.9000 4.8000 ;
	    RECT 68.6000 2.2000 68.9000 4.8000 ;
	    RECT 95.0000 2.2000 95.3000 4.8000 ;
	    RECT 137.4000 3.8000 137.8000 4.2000 ;
	    RECT 137.4000 3.2000 137.7000 3.8000 ;
	    RECT 137.4000 2.8000 137.8000 3.2000 ;
	    RECT 68.6000 1.8000 69.0000 2.2000 ;
	    RECT 95.0000 1.8000 95.4000 2.2000 ;
	    RECT 4.6000 0.8000 5.0000 1.2000 ;
	    RECT 4.6000 -1.8000 4.9000 0.8000 ;
	    RECT 4.6000 -2.2000 5.0000 -1.8000 ;
         LAYER metal3 ;
	    RECT 131.0000 3.1000 131.4000 3.2000 ;
	    RECT 137.4000 3.1000 137.8000 3.2000 ;
	    RECT 131.0000 2.8000 137.8000 3.1000 ;
	    RECT 46.2000 2.1000 46.6000 2.2000 ;
	    RECT 68.6000 2.1000 69.0000 2.2000 ;
	    RECT 95.0000 2.1000 95.4000 2.2000 ;
	    RECT 95.8000 2.1000 96.2000 2.2000 ;
	    RECT 46.2000 1.8000 96.2000 2.1000 ;
	    RECT 4.6000 1.1000 5.0000 1.2000 ;
	    RECT 5.4000 1.1000 5.8000 1.2000 ;
	    RECT 4.6000 0.8000 5.8000 1.1000 ;
         LAYER metal4 ;
	    RECT 131.0000 2.8000 131.4000 3.2000 ;
	    RECT 131.0000 2.2000 131.3000 2.8000 ;
	    RECT 46.2000 1.8000 46.6000 2.2000 ;
	    RECT 95.0000 2.1000 95.4000 2.2000 ;
	    RECT 95.8000 2.1000 96.2000 2.2000 ;
	    RECT 95.0000 1.8000 96.2000 2.1000 ;
	    RECT 131.0000 1.8000 131.4000 2.2000 ;
	    RECT 46.2000 1.2000 46.5000 1.8000 ;
	    RECT 4.6000 1.1000 5.0000 1.2000 ;
	    RECT 5.4000 1.1000 5.8000 1.2000 ;
	    RECT 4.6000 0.8000 5.8000 1.1000 ;
	    RECT 46.2000 0.8000 46.6000 1.2000 ;
         LAYER metal5 ;
	    RECT 95.0000 2.1000 95.4000 2.2000 ;
	    RECT 131.0000 2.1000 131.4000 2.2000 ;
	    RECT 95.0000 1.8000 131.4000 2.1000 ;
	    RECT 4.6000 1.1000 5.0000 1.2000 ;
	    RECT 46.2000 1.1000 46.6000 1.2000 ;
	    RECT 4.6000 0.8000 46.6000 1.1000 ;
      END
   END DATA_B[30]
   PIN DATA_B[29]
      PORT
         LAYER metal1 ;
	    RECT 45.4000 7.8000 45.8000 8.6000 ;
	    RECT 81.4000 7.8000 81.8000 8.6000 ;
	    RECT 106.2000 7.8000 106.6000 8.6000 ;
	    RECT 134.2000 7.8000 134.6000 8.6000 ;
         LAYER metal2 ;
	    RECT 45.4000 7.8000 45.8000 8.2000 ;
	    RECT 81.4000 7.8000 81.8000 8.2000 ;
	    RECT 105.4000 8.1000 105.8000 8.2000 ;
	    RECT 106.2000 8.1000 106.6000 8.2000 ;
	    RECT 105.4000 7.8000 106.6000 8.1000 ;
	    RECT 134.2000 7.8000 134.6000 8.2000 ;
	    RECT 45.4000 5.2000 45.7000 7.8000 ;
	    RECT 81.4000 7.2000 81.7000 7.8000 ;
	    RECT 134.2000 7.2000 134.5000 7.8000 ;
	    RECT 81.4000 6.8000 81.8000 7.2000 ;
	    RECT 134.2000 6.8000 134.6000 7.2000 ;
	    RECT 45.4000 4.8000 45.8000 5.2000 ;
	    RECT 107.8000 1.8000 108.2000 2.2000 ;
	    RECT 107.8000 -1.8000 108.1000 1.8000 ;
	    RECT 107.8000 -2.2000 108.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 105.4000 8.1000 105.8000 8.2000 ;
	    RECT 106.2000 8.1000 106.6000 8.2000 ;
	    RECT 105.4000 7.8000 106.6000 8.1000 ;
	    RECT 80.6000 7.1000 81.0000 7.2000 ;
	    RECT 81.4000 7.1000 81.8000 7.2000 ;
	    RECT 80.6000 6.8000 81.8000 7.1000 ;
	    RECT 133.4000 7.1000 133.8000 7.2000 ;
	    RECT 134.2000 7.1000 134.6000 7.2000 ;
	    RECT 133.4000 6.8000 134.6000 7.1000 ;
	    RECT 45.4000 5.1000 45.8000 5.2000 ;
	    RECT 47.0000 5.1000 47.4000 5.2000 ;
	    RECT 45.4000 4.8000 47.4000 5.1000 ;
	    RECT 106.2000 2.1000 106.6000 2.2000 ;
	    RECT 107.8000 2.1000 108.2000 2.2000 ;
	    RECT 106.2000 1.8000 108.2000 2.1000 ;
         LAYER metal4 ;
	    RECT 106.2000 7.8000 106.6000 8.2000 ;
	    RECT 106.2000 7.2000 106.5000 7.8000 ;
	    RECT 47.0000 6.8000 47.4000 7.2000 ;
	    RECT 80.6000 7.1000 81.0000 7.2000 ;
	    RECT 81.4000 7.1000 81.8000 7.2000 ;
	    RECT 80.6000 6.8000 81.8000 7.1000 ;
	    RECT 106.2000 6.8000 106.6000 7.2000 ;
	    RECT 133.4000 7.1000 133.8000 7.2000 ;
	    RECT 133.4000 6.8000 134.5000 7.1000 ;
	    RECT 47.0000 5.2000 47.3000 6.8000 ;
	    RECT 106.2000 6.2000 106.5000 6.8000 ;
	    RECT 134.2000 6.2000 134.5000 6.8000 ;
	    RECT 106.2000 5.8000 106.6000 6.2000 ;
	    RECT 134.2000 5.8000 134.6000 6.2000 ;
	    RECT 47.0000 4.8000 47.4000 5.2000 ;
	    RECT 106.2000 2.2000 106.5000 5.8000 ;
	    RECT 106.2000 1.8000 106.6000 2.2000 ;
         LAYER metal5 ;
	    RECT 47.0000 7.1000 47.4000 7.2000 ;
	    RECT 81.4000 7.1000 81.8000 7.2000 ;
	    RECT 106.2000 7.1000 106.6000 7.2000 ;
	    RECT 47.0000 6.8000 106.6000 7.1000 ;
	    RECT 106.2000 6.1000 106.6000 6.2000 ;
	    RECT 134.2000 6.1000 134.6000 6.2000 ;
	    RECT 106.2000 5.8000 134.6000 6.1000 ;
      END
   END DATA_B[29]
   PIN DATA_B[28]
      PORT
         LAYER metal1 ;
	    RECT 41.4000 27.8000 41.8000 28.6000 ;
	    RECT 87.8000 27.8000 88.2000 28.6000 ;
	    RECT 25.4000 7.8000 25.8000 8.6000 ;
	    RECT 85.4000 7.8000 85.8000 8.6000 ;
         LAYER metal2 ;
	    RECT 41.4000 27.8000 41.8000 28.2000 ;
	    RECT 87.8000 27.8000 88.2000 28.2000 ;
	    RECT 41.4000 21.2000 41.7000 27.8000 ;
	    RECT 25.4000 20.8000 25.8000 21.2000 ;
	    RECT 41.4000 20.8000 41.8000 21.2000 ;
	    RECT 25.4000 8.2000 25.7000 20.8000 ;
	    RECT 41.4000 19.2000 41.7000 20.8000 ;
	    RECT 87.8000 19.2000 88.1000 27.8000 ;
	    RECT 41.4000 18.8000 41.8000 19.2000 ;
	    RECT 87.8000 18.8000 88.2000 19.2000 ;
	    RECT 85.4000 8.8000 85.8000 9.2000 ;
	    RECT 85.4000 8.2000 85.7000 8.8000 ;
	    RECT 25.4000 7.8000 25.8000 8.2000 ;
	    RECT 85.4000 8.1000 85.8000 8.2000 ;
	    RECT 85.4000 7.8000 86.5000 8.1000 ;
	    RECT 86.2000 -1.8000 86.5000 7.8000 ;
	    RECT 86.2000 -2.2000 86.6000 -1.8000 ;
         LAYER metal3 ;
	    RECT 25.4000 21.1000 25.8000 21.2000 ;
	    RECT 41.4000 21.1000 41.8000 21.2000 ;
	    RECT 25.4000 20.8000 41.8000 21.1000 ;
	    RECT 41.4000 19.1000 41.8000 19.2000 ;
	    RECT 85.4000 19.1000 85.8000 19.2000 ;
	    RECT 87.8000 19.1000 88.2000 19.2000 ;
	    RECT 41.4000 18.8000 88.2000 19.1000 ;
	    RECT 85.4000 8.8000 85.8000 9.2000 ;
	    RECT 85.4000 8.2000 85.7000 8.8000 ;
	    RECT 85.4000 7.8000 85.8000 8.2000 ;
         LAYER metal4 ;
	    RECT 85.4000 18.8000 85.8000 19.2000 ;
	    RECT 85.4000 8.2000 85.7000 18.8000 ;
	    RECT 85.4000 7.8000 85.8000 8.2000 ;
      END
   END DATA_B[28]
   PIN DATA_B[27]
      PORT
         LAYER metal1 ;
	    RECT 47.8000 4.4000 48.2000 5.2000 ;
	    RECT 56.6000 4.4000 57.0000 5.2000 ;
	    RECT 123.8000 4.4000 124.2000 5.2000 ;
	    RECT 147.0000 4.4000 147.4000 5.2000 ;
         LAYER metal2 ;
	    RECT 47.8000 4.8000 48.2000 5.2000 ;
	    RECT 56.6000 4.8000 57.0000 5.2000 ;
	    RECT 123.8000 4.8000 124.2000 5.2000 ;
	    RECT 147.0000 4.8000 147.4000 5.2000 ;
	    RECT 47.8000 4.2000 48.1000 4.8000 ;
	    RECT 56.6000 4.2000 56.9000 4.8000 ;
	    RECT 123.8000 4.2000 124.1000 4.8000 ;
	    RECT 147.0000 4.2000 147.3000 4.8000 ;
	    RECT 47.8000 3.8000 48.2000 4.2000 ;
	    RECT 56.6000 3.8000 57.0000 4.2000 ;
	    RECT 123.8000 3.8000 124.2000 4.2000 ;
	    RECT 126.2000 3.8000 126.6000 4.2000 ;
	    RECT 147.0000 3.8000 147.4000 4.2000 ;
	    RECT 126.2000 -1.8000 126.5000 3.8000 ;
	    RECT 126.2000 -2.2000 126.6000 -1.8000 ;
         LAYER metal3 ;
	    RECT 47.8000 4.8000 56.9000 5.1000 ;
	    RECT 47.8000 4.2000 48.1000 4.8000 ;
	    RECT 56.6000 4.2000 56.9000 4.8000 ;
	    RECT 47.8000 3.8000 48.2000 4.2000 ;
	    RECT 56.6000 4.1000 57.0000 4.2000 ;
	    RECT 123.8000 4.1000 124.2000 4.2000 ;
	    RECT 126.2000 4.1000 126.6000 4.2000 ;
	    RECT 147.0000 4.1000 147.4000 4.2000 ;
	    RECT 56.6000 3.8000 147.4000 4.1000 ;
      END
   END DATA_B[27]
   PIN DATA_B[26]
      PORT
         LAYER metal1 ;
	    RECT 119.0000 52.4000 119.4000 53.2000 ;
	    RECT 151.0000 52.4000 151.4000 53.2000 ;
	    RECT 93.4000 47.8000 93.8000 48.6000 ;
	    RECT 95.0000 47.8000 95.4000 48.6000 ;
         LAYER metal2 ;
	    RECT 151.0000 57.8000 151.4000 58.2000 ;
	    RECT 151.0000 57.2000 151.3000 57.8000 ;
	    RECT 119.0000 56.8000 119.4000 57.2000 ;
	    RECT 151.0000 56.8000 151.4000 57.2000 ;
	    RECT 119.0000 53.2000 119.3000 56.8000 ;
	    RECT 151.0000 53.2000 151.3000 56.8000 ;
	    RECT 95.0000 52.8000 95.4000 53.2000 ;
	    RECT 119.0000 52.8000 119.4000 53.2000 ;
	    RECT 151.0000 52.8000 151.4000 53.2000 ;
	    RECT 95.0000 48.2000 95.3000 52.8000 ;
	    RECT 93.4000 48.1000 93.8000 48.2000 ;
	    RECT 94.2000 48.1000 94.6000 48.2000 ;
	    RECT 93.4000 47.8000 94.6000 48.1000 ;
	    RECT 95.0000 47.8000 95.4000 48.2000 ;
         LAYER metal3 ;
	    RECT 151.0000 58.1000 151.4000 58.2000 ;
	    RECT 173.4000 58.1000 173.8000 58.2000 ;
	    RECT 151.0000 57.8000 173.8000 58.1000 ;
	    RECT 119.0000 57.1000 119.4000 57.2000 ;
	    RECT 151.0000 57.1000 151.4000 57.2000 ;
	    RECT 119.0000 56.8000 151.4000 57.1000 ;
	    RECT 173.4000 55.1000 173.8000 55.2000 ;
	    RECT 175.8000 55.1000 176.2000 55.2000 ;
	    RECT 173.4000 54.8000 176.2000 55.1000 ;
	    RECT 95.0000 53.1000 95.4000 53.2000 ;
	    RECT 119.0000 53.1000 119.4000 53.2000 ;
	    RECT 95.0000 52.8000 119.4000 53.1000 ;
	    RECT 94.2000 48.1000 94.6000 48.2000 ;
	    RECT 95.0000 48.1000 95.4000 48.2000 ;
	    RECT 94.2000 47.8000 95.4000 48.1000 ;
         LAYER metal4 ;
	    RECT 173.4000 57.8000 173.8000 58.2000 ;
	    RECT 173.4000 55.2000 173.7000 57.8000 ;
	    RECT 173.4000 54.8000 173.8000 55.2000 ;
      END
   END DATA_B[26]
   PIN DATA_B[25]
      PORT
         LAYER metal1 ;
	    RECT 39.0000 4.4000 39.4000 5.2000 ;
	    RECT 55.8000 4.4000 56.2000 5.2000 ;
	    RECT 114.2000 4.4000 114.6000 5.2000 ;
	    RECT 140.6000 4.4000 141.0000 5.2000 ;
         LAYER metal2 ;
	    RECT 39.0000 5.8000 39.4000 6.2000 ;
	    RECT 55.8000 5.8000 56.2000 6.2000 ;
	    RECT 114.2000 6.1000 114.6000 6.2000 ;
	    RECT 114.2000 5.8000 115.3000 6.1000 ;
	    RECT 39.0000 5.2000 39.3000 5.8000 ;
	    RECT 55.8000 5.2000 56.1000 5.8000 ;
	    RECT 114.2000 5.2000 114.5000 5.8000 ;
	    RECT 39.0000 4.8000 39.4000 5.2000 ;
	    RECT 55.8000 4.8000 56.2000 5.2000 ;
	    RECT 114.2000 4.8000 114.6000 5.2000 ;
	    RECT 115.0000 -1.8000 115.3000 5.8000 ;
	    RECT 140.6000 5.8000 141.0000 6.2000 ;
	    RECT 140.6000 5.2000 140.9000 5.8000 ;
	    RECT 140.6000 4.8000 141.0000 5.2000 ;
	    RECT 115.0000 -2.2000 115.4000 -1.8000 ;
         LAYER metal3 ;
	    RECT 39.0000 6.1000 39.4000 6.2000 ;
	    RECT 55.8000 6.1000 56.2000 6.2000 ;
	    RECT 66.2000 6.1000 66.6000 6.2000 ;
	    RECT 39.0000 5.8000 66.6000 6.1000 ;
	    RECT 104.6000 6.1000 105.0000 6.2000 ;
	    RECT 114.2000 6.1000 114.6000 6.2000 ;
	    RECT 121.4000 6.1000 121.8000 6.2000 ;
	    RECT 104.6000 5.8000 121.8000 6.1000 ;
	    RECT 139.8000 6.1000 140.2000 6.2000 ;
	    RECT 140.6000 6.1000 141.0000 6.2000 ;
	    RECT 139.8000 5.8000 141.0000 6.1000 ;
         LAYER metal4 ;
	    RECT 66.2000 6.1000 66.6000 6.2000 ;
	    RECT 67.0000 6.1000 67.4000 6.2000 ;
	    RECT 66.2000 5.8000 67.4000 6.1000 ;
	    RECT 103.8000 6.1000 104.2000 6.2000 ;
	    RECT 104.6000 6.1000 105.0000 6.2000 ;
	    RECT 103.8000 5.8000 105.0000 6.1000 ;
	    RECT 121.4000 5.8000 121.8000 6.2000 ;
	    RECT 139.8000 6.1000 140.2000 6.2000 ;
	    RECT 139.8000 5.8000 140.9000 6.1000 ;
	    RECT 121.4000 5.2000 121.7000 5.8000 ;
	    RECT 140.6000 5.2000 140.9000 5.8000 ;
	    RECT 121.4000 4.8000 121.8000 5.2000 ;
	    RECT 140.6000 4.8000 141.0000 5.2000 ;
         LAYER metal5 ;
	    RECT 67.0000 6.1000 67.4000 6.2000 ;
	    RECT 103.8000 6.1000 104.2000 6.2000 ;
	    RECT 67.0000 5.8000 104.2000 6.1000 ;
	    RECT 121.4000 5.1000 121.8000 5.2000 ;
	    RECT 140.6000 5.1000 141.0000 5.2000 ;
	    RECT 121.4000 4.8000 141.0000 5.1000 ;
      END
   END DATA_B[25]
   PIN DATA_B[24]
      PORT
         LAYER metal1 ;
	    RECT 43.0000 45.1000 43.4000 45.2000 ;
	    RECT 43.8000 45.1000 44.2000 45.2000 ;
	    RECT 43.0000 44.8000 44.2000 45.1000 ;
	    RECT 43.0000 44.4000 43.4000 44.8000 ;
	    RECT 81.4000 44.4000 81.8000 45.2000 ;
	    RECT 106.2000 44.4000 106.6000 45.2000 ;
	    RECT 161.4000 44.4000 161.8000 45.2000 ;
         LAYER metal2 ;
	    RECT 43.8000 45.8000 44.2000 46.2000 ;
	    RECT 81.4000 45.8000 81.8000 46.2000 ;
	    RECT 43.8000 45.2000 44.1000 45.8000 ;
	    RECT 81.4000 45.2000 81.7000 45.8000 ;
	    RECT 43.8000 44.8000 44.2000 45.2000 ;
	    RECT 81.4000 44.8000 81.8000 45.2000 ;
	    RECT 105.4000 45.1000 105.8000 45.2000 ;
	    RECT 106.2000 45.1000 106.6000 45.2000 ;
	    RECT 105.4000 44.8000 106.6000 45.1000 ;
	    RECT 160.6000 45.1000 161.0000 45.2000 ;
	    RECT 161.4000 45.1000 161.8000 45.2000 ;
	    RECT 160.6000 44.8000 161.8000 45.1000 ;
         LAYER metal3 ;
	    RECT 173.4000 49.1000 173.8000 49.2000 ;
	    RECT 175.8000 49.1000 176.2000 49.2000 ;
	    RECT 173.4000 48.8000 176.2000 49.1000 ;
	    RECT 43.8000 46.1000 44.2000 46.2000 ;
	    RECT 81.4000 46.1000 81.8000 46.2000 ;
	    RECT 83.0000 46.1000 83.4000 46.2000 ;
	    RECT 43.8000 45.8000 83.4000 46.1000 ;
	    RECT 96.6000 45.1000 97.0000 45.2000 ;
	    RECT 105.4000 45.1000 105.8000 45.2000 ;
	    RECT 107.0000 45.1000 107.4000 45.2000 ;
	    RECT 96.6000 44.8000 107.4000 45.1000 ;
	    RECT 160.6000 45.1000 161.0000 45.2000 ;
	    RECT 161.4000 45.1000 161.8000 45.2000 ;
	    RECT 160.6000 44.8000 161.8000 45.1000 ;
         LAYER metal4 ;
	    RECT 173.4000 48.8000 173.8000 49.2000 ;
	    RECT 83.0000 45.8000 83.4000 46.2000 ;
	    RECT 83.0000 45.2000 83.3000 45.8000 ;
	    RECT 173.4000 45.2000 173.7000 48.8000 ;
	    RECT 83.0000 44.8000 83.4000 45.2000 ;
	    RECT 95.8000 45.1000 96.2000 45.2000 ;
	    RECT 96.6000 45.1000 97.0000 45.2000 ;
	    RECT 95.8000 44.8000 97.0000 45.1000 ;
	    RECT 107.0000 45.1000 107.4000 45.2000 ;
	    RECT 107.8000 45.1000 108.2000 45.2000 ;
	    RECT 107.0000 44.8000 108.2000 45.1000 ;
	    RECT 161.4000 45.1000 161.8000 45.2000 ;
	    RECT 162.2000 45.1000 162.6000 45.2000 ;
	    RECT 161.4000 44.8000 162.6000 45.1000 ;
	    RECT 173.4000 44.8000 173.8000 45.2000 ;
         LAYER metal5 ;
	    RECT 83.0000 45.1000 83.4000 45.2000 ;
	    RECT 95.8000 45.1000 96.2000 45.2000 ;
	    RECT 83.0000 44.8000 96.2000 45.1000 ;
	    RECT 107.8000 45.1000 108.2000 45.2000 ;
	    RECT 162.2000 45.1000 162.6000 45.2000 ;
	    RECT 173.4000 45.1000 173.8000 45.2000 ;
	    RECT 107.8000 44.8000 173.8000 45.1000 ;
      END
   END DATA_B[24]
   PIN DATA_B[23]
      PORT
         LAYER metal1 ;
	    RECT 132.6000 52.4000 133.0000 53.2000 ;
	    RECT 156.6000 52.4000 157.0000 53.2000 ;
	    RECT 47.0000 47.8000 47.4000 48.6000 ;
	    RECT 49.4000 47.8000 49.8000 48.6000 ;
	    RECT 47.0000 47.2000 47.3000 47.8000 ;
	    RECT 47.0000 46.8000 47.4000 47.2000 ;
         LAYER metal2 ;
	    RECT 156.6000 58.8000 157.0000 59.2000 ;
	    RECT 156.6000 53.2000 156.9000 58.8000 ;
	    RECT 132.6000 52.8000 133.0000 53.2000 ;
	    RECT 156.6000 52.8000 157.0000 53.2000 ;
	    RECT 132.6000 49.2000 132.9000 52.8000 ;
	    RECT 156.6000 49.2000 156.9000 52.8000 ;
	    RECT 132.6000 48.8000 133.0000 49.2000 ;
	    RECT 156.6000 48.8000 157.0000 49.2000 ;
	    RECT 47.0000 47.8000 47.4000 48.2000 ;
	    RECT 49.4000 48.1000 49.8000 48.2000 ;
	    RECT 50.2000 48.1000 50.6000 48.2000 ;
	    RECT 49.4000 47.8000 50.6000 48.1000 ;
	    RECT 47.0000 47.2000 47.3000 47.8000 ;
	    RECT 47.0000 46.8000 47.4000 47.2000 ;
         LAYER metal3 ;
	    RECT 156.6000 59.1000 157.0000 59.2000 ;
	    RECT 175.8000 59.1000 176.2000 59.2000 ;
	    RECT 156.6000 58.8000 176.2000 59.1000 ;
	    RECT 132.6000 49.1000 133.0000 49.2000 ;
	    RECT 156.6000 49.1000 157.0000 49.2000 ;
	    RECT 50.2000 48.8000 157.0000 49.1000 ;
	    RECT 50.2000 48.2000 50.5000 48.8000 ;
	    RECT 47.0000 48.1000 47.4000 48.2000 ;
	    RECT 50.2000 48.1000 50.6000 48.2000 ;
	    RECT 47.0000 47.8000 50.6000 48.1000 ;
      END
   END DATA_B[23]
   PIN DATA_B[22]
      PORT
         LAYER metal1 ;
	    RECT 103.8000 32.4000 104.2000 33.2000 ;
	    RECT 40.6000 27.8000 41.0000 28.6000 ;
	    RECT 92.6000 27.8000 93.0000 28.6000 ;
	    RECT 100.6000 12.4000 101.0000 13.2000 ;
         LAYER metal2 ;
	    RECT 103.8000 32.8000 104.2000 33.2000 ;
	    RECT 103.8000 30.2000 104.1000 32.8000 ;
	    RECT 92.6000 29.8000 93.0000 30.2000 ;
	    RECT 103.8000 29.8000 104.2000 30.2000 ;
	    RECT 92.6000 28.2000 92.9000 29.8000 ;
	    RECT 40.6000 27.8000 41.0000 28.2000 ;
	    RECT 92.6000 27.8000 93.0000 28.2000 ;
	    RECT 40.6000 27.2000 40.9000 27.8000 ;
	    RECT 40.6000 26.8000 41.0000 27.2000 ;
	    RECT 103.8000 18.2000 104.1000 29.8000 ;
	    RECT 100.6000 17.8000 101.0000 18.2000 ;
	    RECT 103.8000 17.8000 104.2000 18.2000 ;
	    RECT 100.6000 13.2000 100.9000 17.8000 ;
	    RECT 100.6000 13.1000 101.0000 13.2000 ;
	    RECT 100.6000 12.8000 101.7000 13.1000 ;
	    RECT 101.4000 -1.9000 101.7000 12.8000 ;
	    RECT 102.2000 -1.9000 102.6000 -1.8000 ;
	    RECT 101.4000 -2.2000 102.6000 -1.9000 ;
         LAYER metal3 ;
	    RECT 92.6000 30.1000 93.0000 30.2000 ;
	    RECT 103.8000 30.1000 104.2000 30.2000 ;
	    RECT 51.0000 29.8000 104.2000 30.1000 ;
	    RECT 51.0000 29.1000 51.3000 29.8000 ;
	    RECT 41.4000 28.8000 51.3000 29.1000 ;
	    RECT 41.4000 28.1000 41.7000 28.8000 ;
	    RECT 40.6000 27.8000 41.7000 28.1000 ;
	    RECT 40.6000 27.2000 40.9000 27.8000 ;
	    RECT 40.6000 26.8000 41.0000 27.2000 ;
	    RECT 100.6000 18.1000 101.0000 18.2000 ;
	    RECT 103.8000 18.1000 104.2000 18.2000 ;
	    RECT 100.6000 17.8000 104.2000 18.1000 ;
      END
   END DATA_B[22]
   PIN DATA_B[21]
      PORT
         LAYER metal1 ;
	    RECT 31.8000 7.8000 32.2000 8.6000 ;
	    RECT 74.2000 7.8000 74.6000 8.6000 ;
	    RECT 107.0000 7.8000 107.4000 8.6000 ;
	    RECT 128.6000 7.8000 129.0000 8.6000 ;
         LAYER metal2 ;
	    RECT 128.6000 8.8000 129.0000 9.2000 ;
	    RECT 128.6000 8.2000 128.9000 8.8000 ;
	    RECT 31.8000 8.1000 32.2000 8.2000 ;
	    RECT 32.6000 8.1000 33.0000 8.2000 ;
	    RECT 31.8000 7.8000 33.0000 8.1000 ;
	    RECT 74.2000 7.8000 74.6000 8.2000 ;
	    RECT 107.0000 8.1000 107.4000 8.2000 ;
	    RECT 107.8000 8.1000 108.2000 8.2000 ;
	    RECT 107.0000 7.8000 108.2000 8.1000 ;
	    RECT 113.4000 7.8000 113.8000 8.2000 ;
	    RECT 128.6000 7.8000 129.0000 8.2000 ;
	    RECT 74.2000 7.2000 74.5000 7.8000 ;
	    RECT 74.2000 6.8000 74.6000 7.2000 ;
	    RECT 113.4000 -1.8000 113.7000 7.8000 ;
	    RECT 113.4000 -2.2000 113.8000 -1.8000 ;
         LAYER metal3 ;
	    RECT 128.6000 8.8000 129.0000 9.2000 ;
	    RECT 32.6000 8.1000 33.0000 8.2000 ;
	    RECT 107.0000 8.1000 107.4000 8.2000 ;
	    RECT 107.8000 8.1000 108.2000 8.2000 ;
	    RECT 113.4000 8.1000 113.8000 8.2000 ;
	    RECT 128.6000 8.1000 128.9000 8.8000 ;
	    RECT 31.8000 7.8000 53.7000 8.1000 ;
	    RECT 107.0000 7.8000 128.9000 8.1000 ;
	    RECT 53.4000 7.1000 53.7000 7.8000 ;
	    RECT 74.2000 7.1000 74.6000 7.2000 ;
	    RECT 79.8000 7.1000 80.2000 7.2000 ;
	    RECT 53.4000 6.8000 80.2000 7.1000 ;
         LAYER metal4 ;
	    RECT 79.8000 7.8000 80.2000 8.2000 ;
	    RECT 107.0000 7.8000 107.4000 8.2000 ;
	    RECT 79.8000 7.2000 80.1000 7.8000 ;
	    RECT 107.0000 7.2000 107.3000 7.8000 ;
	    RECT 79.8000 6.8000 80.2000 7.2000 ;
	    RECT 107.0000 6.8000 107.4000 7.2000 ;
         LAYER metal5 ;
	    RECT 79.8000 8.1000 80.2000 8.2000 ;
	    RECT 79.8000 7.8000 107.3000 8.1000 ;
	    RECT 107.0000 7.2000 107.3000 7.8000 ;
	    RECT 107.0000 6.8000 107.4000 7.2000 ;
      END
   END DATA_B[21]
   PIN DATA_B[20]
      PORT
         LAYER metal1 ;
	    RECT 43.8000 7.8000 44.2000 8.6000 ;
	    RECT 51.0000 7.8000 51.4000 8.6000 ;
	    RECT 92.6000 7.8000 93.0000 8.6000 ;
	    RECT 130.2000 7.8000 130.6000 8.6000 ;
         LAYER metal2 ;
	    RECT 43.8000 7.8000 44.2000 8.2000 ;
	    RECT 51.0000 7.8000 51.4000 8.2000 ;
	    RECT 92.6000 8.1000 93.0000 8.2000 ;
	    RECT 91.8000 7.8000 93.0000 8.1000 ;
	    RECT 130.2000 7.8000 130.6000 8.2000 ;
	    RECT 43.8000 3.2000 44.1000 7.8000 ;
	    RECT 51.0000 3.2000 51.3000 7.8000 ;
	    RECT 91.8000 3.2000 92.1000 7.8000 ;
	    RECT 130.2000 3.2000 130.5000 7.8000 ;
	    RECT 43.8000 2.8000 44.2000 3.2000 ;
	    RECT 51.0000 2.8000 51.4000 3.2000 ;
	    RECT 91.8000 2.8000 92.2000 3.2000 ;
	    RECT 130.2000 2.8000 130.6000 3.2000 ;
	    RECT 91.8000 1.2000 92.1000 2.8000 ;
	    RECT 91.8000 0.8000 92.2000 1.2000 ;
	    RECT 91.8000 -1.8000 92.1000 0.8000 ;
	    RECT 91.8000 -2.2000 92.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 43.8000 3.1000 44.2000 3.2000 ;
	    RECT 51.0000 3.1000 51.4000 3.2000 ;
	    RECT 61.4000 3.1000 61.8000 3.2000 ;
	    RECT 43.8000 2.8000 61.8000 3.1000 ;
	    RECT 91.8000 3.1000 92.2000 3.2000 ;
	    RECT 130.2000 3.1000 130.6000 3.2000 ;
	    RECT 91.8000 2.8000 130.6000 3.1000 ;
	    RECT 91.0000 1.1000 91.4000 1.2000 ;
	    RECT 91.8000 1.1000 92.2000 1.2000 ;
	    RECT 91.0000 0.8000 92.2000 1.1000 ;
         LAYER metal4 ;
	    RECT 61.4000 2.8000 61.8000 3.2000 ;
	    RECT 61.4000 2.2000 61.7000 2.8000 ;
	    RECT 61.4000 1.8000 61.8000 2.2000 ;
	    RECT 91.8000 1.8000 92.2000 2.2000 ;
	    RECT 91.0000 1.1000 91.4000 1.2000 ;
	    RECT 91.8000 1.1000 92.1000 1.8000 ;
	    RECT 91.0000 0.8000 92.1000 1.1000 ;
         LAYER metal5 ;
	    RECT 61.4000 2.1000 61.8000 2.2000 ;
	    RECT 91.8000 2.1000 92.2000 2.2000 ;
	    RECT 61.4000 1.8000 92.2000 2.1000 ;
      END
   END DATA_B[20]
   PIN DATA_B[19]
      PORT
         LAYER metal1 ;
	    RECT 67.8000 7.8000 68.2000 8.6000 ;
	    RECT 78.2000 7.8000 78.6000 8.6000 ;
	    RECT 127.8000 7.8000 128.2000 8.6000 ;
	    RECT 143.0000 7.8000 143.4000 8.6000 ;
         LAYER metal2 ;
	    RECT 67.8000 7.8000 68.2000 8.2000 ;
	    RECT 78.2000 7.8000 78.6000 8.2000 ;
	    RECT 127.8000 7.8000 128.2000 8.2000 ;
	    RECT 143.0000 7.8000 143.4000 8.2000 ;
	    RECT 67.8000 6.2000 68.1000 7.8000 ;
	    RECT 78.2000 6.2000 78.5000 7.8000 ;
	    RECT 67.8000 5.8000 68.2000 6.2000 ;
	    RECT 78.2000 5.8000 78.6000 6.2000 ;
	    RECT 127.8000 5.2000 128.1000 7.8000 ;
	    RECT 143.0000 5.2000 143.3000 7.8000 ;
	    RECT 127.8000 4.8000 128.2000 5.2000 ;
	    RECT 143.0000 4.8000 143.4000 5.2000 ;
	    RECT 127.8000 -1.8000 128.1000 4.8000 ;
	    RECT 127.8000 -2.2000 128.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 67.8000 6.1000 68.2000 6.2000 ;
	    RECT 78.2000 6.1000 78.6000 6.2000 ;
	    RECT 67.8000 5.8000 78.6000 6.1000 ;
	    RECT 78.2000 5.1000 78.5000 5.8000 ;
	    RECT 127.8000 5.1000 128.2000 5.2000 ;
	    RECT 143.0000 5.1000 143.4000 5.2000 ;
	    RECT 78.2000 4.8000 143.4000 5.1000 ;
      END
   END DATA_B[19]
   PIN DATA_B[18]
      PORT
         LAYER metal1 ;
	    RECT 127.8000 33.8000 128.2000 34.2000 ;
	    RECT 127.8000 33.2000 128.1000 33.8000 ;
	    RECT 50.2000 32.4000 50.6000 33.2000 ;
	    RECT 83.0000 32.4000 83.4000 33.2000 ;
	    RECT 127.8000 32.4000 128.2000 33.2000 ;
	    RECT 0.6000 27.8000 1.0000 28.6000 ;
         LAYER metal2 ;
	    RECT 127.8000 33.8000 128.2000 34.2000 ;
	    RECT 127.8000 33.2000 128.1000 33.8000 ;
	    RECT 50.2000 32.8000 50.6000 33.2000 ;
	    RECT 83.0000 33.1000 83.4000 33.2000 ;
	    RECT 83.8000 33.1000 84.2000 33.2000 ;
	    RECT 83.0000 32.8000 84.2000 33.1000 ;
	    RECT 127.8000 32.8000 128.2000 33.2000 ;
	    RECT 50.2000 32.2000 50.5000 32.8000 ;
	    RECT 50.2000 31.8000 50.6000 32.2000 ;
	    RECT 0.6000 29.8000 1.0000 30.2000 ;
	    RECT 0.6000 28.2000 0.9000 29.8000 ;
	    RECT 0.6000 27.8000 1.0000 28.2000 ;
         LAYER metal3 ;
	    RECT 83.0000 33.1000 83.4000 33.2000 ;
	    RECT 83.8000 33.1000 84.2000 33.2000 ;
	    RECT 83.0000 32.8000 84.2000 33.1000 ;
	    RECT 126.2000 33.1000 126.6000 33.2000 ;
	    RECT 127.8000 33.1000 128.2000 33.2000 ;
	    RECT 126.2000 32.8000 128.2000 33.1000 ;
	    RECT 50.2000 32.1000 50.6000 32.2000 ;
	    RECT 51.0000 32.1000 51.4000 32.2000 ;
	    RECT 50.2000 31.8000 51.4000 32.1000 ;
	    RECT -2.6000 30.1000 -2.2000 30.2000 ;
	    RECT 0.6000 30.1000 1.0000 30.2000 ;
	    RECT 50.2000 30.1000 50.6000 30.2000 ;
	    RECT -2.6000 29.8000 50.6000 30.1000 ;
         LAYER metal4 ;
	    RECT 83.0000 32.8000 83.4000 33.2000 ;
	    RECT 126.2000 32.8000 126.6000 33.2000 ;
	    RECT 83.0000 32.2000 83.3000 32.8000 ;
	    RECT 126.2000 32.2000 126.5000 32.8000 ;
	    RECT 50.2000 32.1000 50.6000 32.2000 ;
	    RECT 51.0000 32.1000 51.4000 32.2000 ;
	    RECT 50.2000 31.8000 51.4000 32.1000 ;
	    RECT 83.0000 31.8000 83.4000 32.2000 ;
	    RECT 126.2000 31.8000 126.6000 32.2000 ;
	    RECT 50.2000 30.2000 50.5000 31.8000 ;
	    RECT 50.2000 29.8000 50.6000 30.2000 ;
         LAYER metal5 ;
	    RECT 50.2000 32.1000 50.6000 32.2000 ;
	    RECT 83.0000 32.1000 83.4000 32.2000 ;
	    RECT 126.2000 32.1000 126.6000 32.2000 ;
	    RECT 50.2000 31.8000 126.6000 32.1000 ;
      END
   END DATA_B[18]
   PIN DATA_B[17]
      PORT
         LAYER metal1 ;
	    RECT 132.6000 32.4000 133.0000 33.2000 ;
	    RECT 103.0000 27.8000 103.4000 28.6000 ;
	    RECT 16.6000 7.8000 17.0000 8.6000 ;
	    RECT 65.4000 7.8000 65.8000 8.6000 ;
         LAYER metal2 ;
	    RECT 131.8000 33.1000 132.2000 33.2000 ;
	    RECT 132.6000 33.1000 133.0000 33.2000 ;
	    RECT 131.8000 32.8000 133.0000 33.1000 ;
	    RECT 103.0000 27.8000 103.4000 28.2000 ;
	    RECT 103.0000 21.2000 103.3000 27.8000 ;
	    RECT 103.0000 20.8000 103.4000 21.2000 ;
	    RECT 16.6000 8.8000 17.0000 9.2000 ;
	    RECT 65.4000 8.8000 65.8000 9.2000 ;
	    RECT 16.6000 8.2000 16.9000 8.8000 ;
	    RECT 65.4000 8.2000 65.7000 8.8000 ;
	    RECT 16.6000 7.8000 17.0000 8.2000 ;
	    RECT 65.4000 7.8000 65.8000 8.2000 ;
	    RECT 106.2000 0.8000 106.6000 1.2000 ;
	    RECT 106.2000 -1.8000 106.5000 0.8000 ;
	    RECT 106.2000 -2.2000 106.6000 -1.8000 ;
         LAYER metal3 ;
	    RECT 131.8000 33.1000 132.2000 33.2000 ;
	    RECT 132.6000 33.1000 133.0000 33.2000 ;
	    RECT 131.8000 32.8000 133.0000 33.1000 ;
	    RECT 79.8000 21.1000 80.2000 21.2000 ;
	    RECT 103.0000 21.1000 103.4000 21.2000 ;
	    RECT 105.4000 21.1000 105.8000 21.2000 ;
	    RECT 79.8000 20.8000 105.8000 21.1000 ;
	    RECT 16.6000 9.1000 17.0000 9.2000 ;
	    RECT 65.4000 9.1000 65.8000 9.2000 ;
	    RECT 79.8000 9.1000 80.2000 9.2000 ;
	    RECT 16.6000 8.8000 80.2000 9.1000 ;
	    RECT 105.4000 1.1000 105.8000 1.2000 ;
	    RECT 106.2000 1.1000 106.6000 1.2000 ;
	    RECT 105.4000 0.8000 106.6000 1.1000 ;
         LAYER metal4 ;
	    RECT 132.6000 32.8000 133.0000 33.2000 ;
	    RECT 132.6000 24.2000 132.9000 32.8000 ;
	    RECT 105.4000 23.8000 105.8000 24.2000 ;
	    RECT 132.6000 23.8000 133.0000 24.2000 ;
	    RECT 105.4000 21.2000 105.7000 23.8000 ;
	    RECT 79.8000 20.8000 80.2000 21.2000 ;
	    RECT 105.4000 20.8000 105.8000 21.2000 ;
	    RECT 79.8000 9.2000 80.1000 20.8000 ;
	    RECT 79.8000 8.8000 80.2000 9.2000 ;
	    RECT 105.4000 1.2000 105.7000 20.8000 ;
	    RECT 105.4000 0.8000 105.8000 1.2000 ;
         LAYER metal5 ;
	    RECT 105.4000 24.1000 105.8000 24.2000 ;
	    RECT 132.6000 24.1000 133.0000 24.2000 ;
	    RECT 105.4000 23.8000 133.0000 24.1000 ;
      END
   END DATA_B[17]
   PIN DATA_B[16]
      PORT
         LAYER metal1 ;
	    RECT 38.2000 33.8000 38.6000 34.2000 ;
	    RECT 38.2000 33.2000 38.5000 33.8000 ;
	    RECT 38.2000 32.4000 38.6000 33.2000 ;
	    RECT 87.0000 32.4000 87.4000 33.2000 ;
	    RECT 167.8000 32.4000 168.2000 33.2000 ;
	    RECT 45.4000 27.8000 45.8000 28.6000 ;
         LAYER metal2 ;
	    RECT 38.2000 33.8000 38.6000 34.2000 ;
	    RECT 167.8000 33.8000 168.2000 34.2000 ;
	    RECT 38.2000 33.2000 38.5000 33.8000 ;
	    RECT 167.8000 33.2000 168.1000 33.8000 ;
	    RECT 38.2000 32.8000 38.6000 33.2000 ;
	    RECT 45.4000 32.8000 45.8000 33.2000 ;
	    RECT 86.2000 33.1000 86.6000 33.2000 ;
	    RECT 87.0000 33.1000 87.4000 33.2000 ;
	    RECT 86.2000 32.8000 87.4000 33.1000 ;
	    RECT 167.8000 32.8000 168.2000 33.2000 ;
	    RECT 45.4000 28.2000 45.7000 32.8000 ;
	    RECT 45.4000 27.8000 45.8000 28.2000 ;
         LAYER metal3 ;
	    RECT 167.8000 33.8000 168.2000 34.2000 ;
	    RECT 38.2000 33.1000 38.6000 33.2000 ;
	    RECT 45.4000 33.1000 45.8000 33.2000 ;
	    RECT 53.4000 33.1000 53.8000 33.2000 ;
	    RECT 38.2000 32.8000 53.8000 33.1000 ;
	    RECT 86.2000 33.1000 86.6000 33.2000 ;
	    RECT 87.0000 33.1000 87.4000 33.2000 ;
	    RECT 86.2000 32.8000 87.4000 33.1000 ;
	    RECT 147.8000 33.1000 148.2000 33.2000 ;
	    RECT 167.8000 33.1000 168.1000 33.8000 ;
	    RECT 175.8000 33.1000 176.2000 33.2000 ;
	    RECT 147.8000 32.8000 176.2000 33.1000 ;
         LAYER metal4 ;
	    RECT 53.4000 33.1000 53.8000 33.2000 ;
	    RECT 54.2000 33.1000 54.6000 33.2000 ;
	    RECT 53.4000 32.8000 54.6000 33.1000 ;
	    RECT 86.2000 33.1000 86.6000 33.2000 ;
	    RECT 87.0000 33.1000 87.4000 33.2000 ;
	    RECT 86.2000 32.8000 87.4000 33.1000 ;
	    RECT 147.0000 33.1000 147.4000 33.2000 ;
	    RECT 147.8000 33.1000 148.2000 33.2000 ;
	    RECT 147.0000 32.8000 148.2000 33.1000 ;
         LAYER metal5 ;
	    RECT 54.2000 33.1000 54.6000 33.2000 ;
	    RECT 86.2000 33.1000 86.6000 33.2000 ;
	    RECT 147.0000 33.1000 147.4000 33.2000 ;
	    RECT 54.2000 32.8000 147.4000 33.1000 ;
      END
   END DATA_B[16]
   PIN DATA_B[15]
      PORT
         LAYER metal1 ;
	    RECT 37.3000 46.8000 37.8000 47.2000 ;
	    RECT 75.7000 46.8000 76.2000 47.2000 ;
	    RECT 133.3000 46.8000 133.8000 47.2000 ;
	    RECT 170.1000 46.8000 170.6000 47.2000 ;
	    RECT 37.2000 46.4000 37.6000 46.8000 ;
	    RECT 75.6000 46.4000 76.0000 46.8000 ;
	    RECT 133.2000 46.4000 133.6000 46.8000 ;
	    RECT 170.0000 46.4000 170.4000 46.8000 ;
         LAYER metal2 ;
	    RECT 37.4000 51.8000 37.8000 52.2000 ;
	    RECT 75.8000 51.8000 76.2000 52.2000 ;
	    RECT 133.4000 51.8000 133.8000 52.2000 ;
	    RECT 170.2000 51.8000 170.6000 52.2000 ;
	    RECT 37.4000 47.2000 37.7000 51.8000 ;
	    RECT 75.8000 47.2000 76.1000 51.8000 ;
	    RECT 133.4000 47.2000 133.7000 51.8000 ;
	    RECT 170.2000 47.2000 170.5000 51.8000 ;
	    RECT 37.4000 46.8000 37.8000 47.2000 ;
	    RECT 75.8000 46.8000 76.2000 47.2000 ;
	    RECT 133.4000 46.8000 133.8000 47.2000 ;
	    RECT 170.2000 46.8000 170.6000 47.2000 ;
         LAYER metal3 ;
	    RECT 175.8000 53.1000 176.2000 53.2000 ;
	    RECT 170.2000 52.8000 176.2000 53.1000 ;
	    RECT 170.2000 52.2000 170.5000 52.8000 ;
	    RECT 37.4000 52.1000 37.8000 52.2000 ;
	    RECT 75.8000 52.1000 76.2000 52.2000 ;
	    RECT 133.4000 52.1000 133.8000 52.2000 ;
	    RECT 170.2000 52.1000 170.6000 52.2000 ;
	    RECT 37.4000 51.8000 170.6000 52.1000 ;
      END
   END DATA_B[15]
   PIN DATA_B[14]
      PORT
         LAYER metal1 ;
	    RECT 77.4000 12.4000 77.8000 13.2000 ;
	    RECT 137.4000 12.4000 137.8000 13.2000 ;
	    RECT 11.8000 7.8000 12.2000 8.6000 ;
	    RECT 95.8000 7.8000 96.2000 8.6000 ;
         LAYER metal2 ;
	    RECT 77.4000 12.8000 77.8000 13.2000 ;
	    RECT 137.4000 12.8000 137.8000 13.2000 ;
	    RECT 77.4000 10.2000 77.7000 12.8000 ;
	    RECT 137.4000 10.2000 137.7000 12.8000 ;
	    RECT 11.8000 9.8000 12.2000 10.2000 ;
	    RECT 14.2000 9.8000 14.6000 10.2000 ;
	    RECT 77.4000 9.8000 77.8000 10.2000 ;
	    RECT 137.4000 9.8000 137.8000 10.2000 ;
	    RECT 11.8000 8.2000 12.1000 9.8000 ;
	    RECT 11.8000 7.8000 12.2000 8.2000 ;
	    RECT 13.4000 -1.9000 13.8000 -1.8000 ;
	    RECT 14.2000 -1.9000 14.5000 9.8000 ;
	    RECT 95.8000 8.1000 96.2000 8.2000 ;
	    RECT 96.6000 8.1000 97.0000 8.2000 ;
	    RECT 95.8000 7.8000 97.0000 8.1000 ;
	    RECT 13.4000 -2.2000 14.5000 -1.9000 ;
         LAYER metal3 ;
	    RECT 11.8000 10.1000 12.2000 10.2000 ;
	    RECT 14.2000 10.1000 14.6000 10.2000 ;
	    RECT 77.4000 10.1000 77.8000 10.2000 ;
	    RECT 95.8000 10.1000 96.2000 10.2000 ;
	    RECT 11.8000 9.8000 96.2000 10.1000 ;
	    RECT 113.4000 10.1000 113.8000 10.2000 ;
	    RECT 137.4000 10.1000 137.8000 10.2000 ;
	    RECT 113.4000 9.8000 137.8000 10.1000 ;
	    RECT 95.8000 8.1000 96.2000 8.2000 ;
	    RECT 96.6000 8.1000 97.0000 8.2000 ;
	    RECT 95.8000 7.8000 97.0000 8.1000 ;
         LAYER metal4 ;
	    RECT 95.8000 9.8000 96.2000 10.2000 ;
	    RECT 113.4000 9.8000 113.8000 10.2000 ;
	    RECT 95.8000 9.2000 96.1000 9.8000 ;
	    RECT 113.4000 9.2000 113.7000 9.8000 ;
	    RECT 95.8000 8.8000 96.2000 9.2000 ;
	    RECT 113.4000 8.8000 113.8000 9.2000 ;
	    RECT 95.8000 8.2000 96.1000 8.8000 ;
	    RECT 95.8000 7.8000 96.2000 8.2000 ;
         LAYER metal5 ;
	    RECT 95.8000 9.1000 96.2000 9.2000 ;
	    RECT 113.4000 9.1000 113.8000 9.2000 ;
	    RECT 95.8000 8.8000 113.8000 9.1000 ;
      END
   END DATA_B[14]
   PIN DATA_B[13]
      PORT
         LAYER metal1 ;
	    RECT 39.6000 14.2000 40.0000 14.6000 ;
	    RECT 89.2000 14.2000 89.6000 14.6000 ;
	    RECT 120.4000 14.2000 120.8000 14.6000 ;
	    RECT 39.7000 14.1000 40.2000 14.2000 ;
	    RECT 40.6000 14.1000 41.0000 14.2000 ;
	    RECT 39.7000 13.8000 41.0000 14.1000 ;
	    RECT 89.3000 13.8000 89.8000 14.2000 ;
	    RECT 120.5000 13.8000 121.0000 14.2000 ;
	    RECT 155.8000 6.8000 156.3000 7.2000 ;
	    RECT 156.0000 6.4000 156.4000 6.8000 ;
         LAYER metal2 ;
	    RECT 39.8000 14.1000 40.2000 14.2000 ;
	    RECT 40.6000 14.1000 41.0000 14.2000 ;
	    RECT 39.8000 13.8000 41.0000 14.1000 ;
	    RECT 89.4000 13.8000 89.8000 14.2000 ;
	    RECT 120.6000 13.8000 121.0000 14.2000 ;
	    RECT 89.4000 13.2000 89.7000 13.8000 ;
	    RECT 120.6000 13.2000 120.9000 13.8000 ;
	    RECT 89.4000 12.8000 89.8000 13.2000 ;
	    RECT 120.6000 12.8000 121.0000 13.2000 ;
	    RECT 155.8000 6.8000 156.2000 7.2000 ;
	    RECT 155.8000 2.2000 156.1000 6.8000 ;
	    RECT 155.8000 1.8000 156.2000 2.2000 ;
	    RECT 155.8000 -1.8000 156.1000 1.8000 ;
	    RECT 155.8000 -2.2000 156.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 39.8000 14.1000 40.2000 14.2000 ;
	    RECT 40.6000 14.1000 41.0000 14.2000 ;
	    RECT 39.8000 13.8000 41.0000 14.1000 ;
	    RECT 88.6000 13.1000 89.0000 13.2000 ;
	    RECT 89.4000 13.1000 89.8000 13.2000 ;
	    RECT 88.6000 12.8000 89.8000 13.1000 ;
	    RECT 119.8000 13.1000 120.2000 13.2000 ;
	    RECT 120.6000 13.1000 121.0000 13.2000 ;
	    RECT 119.8000 12.8000 121.0000 13.1000 ;
	    RECT 120.6000 2.1000 121.0000 2.2000 ;
	    RECT 155.8000 2.1000 156.2000 2.2000 ;
	    RECT 120.6000 1.8000 156.2000 2.1000 ;
         LAYER metal4 ;
	    RECT 40.6000 13.8000 41.0000 14.2000 ;
	    RECT 40.6000 12.2000 40.9000 13.8000 ;
	    RECT 88.6000 13.1000 89.0000 13.2000 ;
	    RECT 119.8000 13.1000 120.2000 13.2000 ;
	    RECT 88.6000 12.8000 89.7000 13.1000 ;
	    RECT 119.8000 12.8000 120.9000 13.1000 ;
	    RECT 89.4000 12.2000 89.7000 12.8000 ;
	    RECT 120.6000 12.2000 120.9000 12.8000 ;
	    RECT 40.6000 11.8000 41.0000 12.2000 ;
	    RECT 89.4000 11.8000 89.8000 12.2000 ;
	    RECT 120.6000 11.8000 121.0000 12.2000 ;
	    RECT 120.6000 2.2000 120.9000 11.8000 ;
	    RECT 120.6000 1.8000 121.0000 2.2000 ;
         LAYER metal5 ;
	    RECT 40.6000 12.1000 41.0000 12.2000 ;
	    RECT 89.4000 12.1000 89.8000 12.2000 ;
	    RECT 120.6000 12.1000 121.0000 12.2000 ;
	    RECT 40.6000 11.8000 121.0000 12.1000 ;
      END
   END DATA_B[13]
   PIN DATA_B[12]
      PORT
         LAYER metal1 ;
	    RECT 50.2000 26.8000 50.7000 27.2000 ;
	    RECT 119.8000 26.8000 120.3000 27.2000 ;
	    RECT 50.4000 26.4000 50.8000 26.8000 ;
	    RECT 120.0000 26.4000 120.4000 26.8000 ;
	    RECT 105.6000 14.2000 106.0000 14.6000 ;
	    RECT 105.4000 13.8000 105.9000 14.2000 ;
	    RECT 13.4000 6.8000 13.9000 7.2000 ;
	    RECT 13.6000 6.4000 14.0000 6.8000 ;
         LAYER metal2 ;
	    RECT 50.2000 26.8000 50.6000 27.2000 ;
	    RECT 119.8000 26.8000 120.2000 27.2000 ;
	    RECT 50.2000 26.2000 50.5000 26.8000 ;
	    RECT 50.2000 25.8000 50.6000 26.2000 ;
	    RECT 119.8000 24.2000 120.1000 26.8000 ;
	    RECT 105.4000 23.8000 105.8000 24.2000 ;
	    RECT 119.8000 23.8000 120.2000 24.2000 ;
	    RECT 105.4000 14.2000 105.7000 23.8000 ;
	    RECT 105.4000 13.8000 105.8000 14.2000 ;
	    RECT 13.4000 6.8000 13.8000 7.2000 ;
	    RECT 13.4000 1.2000 13.7000 6.8000 ;
	    RECT 13.4000 0.8000 13.8000 1.2000 ;
	    RECT 15.8000 0.8000 16.2000 1.2000 ;
	    RECT 15.8000 -1.8000 16.1000 0.8000 ;
	    RECT 15.8000 -2.2000 16.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 50.2000 26.8000 50.6000 27.2000 ;
	    RECT 50.2000 26.2000 50.5000 26.8000 ;
	    RECT 50.2000 25.8000 50.6000 26.2000 ;
	    RECT 50.2000 24.1000 50.6000 24.2000 ;
	    RECT 105.4000 24.1000 105.8000 24.2000 ;
	    RECT 119.8000 24.1000 120.2000 24.2000 ;
	    RECT 50.2000 23.8000 120.2000 24.1000 ;
	    RECT 13.4000 1.1000 13.8000 1.2000 ;
	    RECT 15.8000 1.1000 16.2000 1.2000 ;
	    RECT 50.2000 1.1000 50.6000 1.2000 ;
	    RECT 13.4000 0.8000 50.6000 1.1000 ;
         LAYER metal4 ;
	    RECT 50.2000 26.8000 50.6000 27.2000 ;
	    RECT 50.2000 24.2000 50.5000 26.8000 ;
	    RECT 50.2000 23.8000 50.6000 24.2000 ;
	    RECT 50.2000 1.2000 50.5000 23.8000 ;
	    RECT 50.2000 0.8000 50.6000 1.2000 ;
      END
   END DATA_B[12]
   PIN DATA_B[11]
      PORT
         LAYER metal1 ;
	    RECT 48.6000 13.8000 49.0000 14.2000 ;
	    RECT 48.6000 13.2000 48.9000 13.8000 ;
	    RECT 48.6000 12.4000 49.0000 13.2000 ;
	    RECT 62.2000 12.4000 62.6000 13.2000 ;
	    RECT 146.2000 12.4000 146.6000 13.2000 ;
	    RECT 168.6000 12.4000 169.0000 13.2000 ;
         LAYER metal2 ;
	    RECT 168.6000 14.8000 169.0000 15.2000 ;
	    RECT 48.6000 13.8000 49.0000 14.2000 ;
	    RECT 62.2000 13.8000 62.6000 14.2000 ;
	    RECT 48.6000 13.2000 48.9000 13.8000 ;
	    RECT 62.2000 13.2000 62.5000 13.8000 ;
	    RECT 168.6000 13.2000 168.9000 14.8000 ;
	    RECT 48.6000 12.8000 49.0000 13.2000 ;
	    RECT 61.4000 13.1000 61.8000 13.2000 ;
	    RECT 62.2000 13.1000 62.6000 13.2000 ;
	    RECT 61.4000 12.8000 62.6000 13.1000 ;
	    RECT 145.4000 13.1000 145.8000 13.2000 ;
	    RECT 146.2000 13.1000 146.6000 13.2000 ;
	    RECT 145.4000 12.8000 146.6000 13.1000 ;
	    RECT 167.8000 13.1000 168.2000 13.2000 ;
	    RECT 168.6000 13.1000 169.0000 13.2000 ;
	    RECT 167.8000 12.8000 169.0000 13.1000 ;
         LAYER metal3 ;
	    RECT 168.6000 15.1000 169.0000 15.2000 ;
	    RECT 175.8000 15.1000 176.2000 15.2000 ;
	    RECT 168.6000 14.8000 176.2000 15.1000 ;
	    RECT 62.2000 14.1000 62.6000 14.2000 ;
	    RECT 62.2000 13.8000 134.5000 14.1000 ;
	    RECT 48.6000 13.1000 49.0000 13.2000 ;
	    RECT 61.4000 13.1000 61.8000 13.2000 ;
	    RECT 48.6000 12.8000 61.8000 13.1000 ;
	    RECT 134.2000 13.1000 134.5000 13.8000 ;
	    RECT 145.4000 13.1000 145.8000 13.2000 ;
	    RECT 167.8000 13.1000 168.2000 13.2000 ;
	    RECT 134.2000 12.8000 168.2000 13.1000 ;
      END
   END DATA_B[11]
   PIN DATA_B[10]
      PORT
         LAYER metal1 ;
	    RECT 139.2000 54.2000 139.6000 54.6000 ;
	    RECT 138.2000 54.1000 138.6000 54.2000 ;
	    RECT 139.0000 54.1000 139.5000 54.2000 ;
	    RECT 138.2000 53.8000 139.5000 54.1000 ;
	    RECT 22.1000 46.8000 22.6000 47.2000 ;
	    RECT 88.5000 46.8000 89.0000 47.2000 ;
	    RECT 120.5000 46.8000 121.0000 47.2000 ;
	    RECT 22.0000 46.4000 22.4000 46.8000 ;
	    RECT 88.4000 46.4000 88.8000 46.8000 ;
	    RECT 120.4000 46.4000 120.8000 46.8000 ;
         LAYER metal2 ;
	    RECT 138.2000 54.1000 138.6000 54.2000 ;
	    RECT 137.4000 53.8000 138.6000 54.1000 ;
	    RECT 120.6000 47.8000 121.0000 48.2000 ;
	    RECT 120.6000 47.2000 120.9000 47.8000 ;
	    RECT 137.4000 47.2000 137.7000 53.8000 ;
	    RECT 22.2000 46.8000 22.6000 47.2000 ;
	    RECT 88.6000 46.8000 89.0000 47.2000 ;
	    RECT 120.6000 47.1000 121.0000 47.2000 ;
	    RECT 121.4000 47.1000 121.8000 47.2000 ;
	    RECT 120.6000 46.8000 121.8000 47.1000 ;
	    RECT 137.4000 46.8000 137.8000 47.2000 ;
	    RECT 22.2000 46.2000 22.5000 46.8000 ;
	    RECT 88.6000 46.2000 88.9000 46.8000 ;
	    RECT 22.2000 45.8000 22.6000 46.2000 ;
	    RECT 88.6000 45.8000 89.0000 46.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 49.1000 -2.2000 49.2000 ;
	    RECT 1.4000 49.1000 1.8000 49.2000 ;
	    RECT -2.6000 48.8000 1.8000 49.1000 ;
	    RECT 95.8000 48.1000 96.2000 48.2000 ;
	    RECT 120.6000 48.1000 121.0000 48.2000 ;
	    RECT 95.8000 47.8000 121.0000 48.1000 ;
	    RECT 22.2000 46.8000 22.6000 47.2000 ;
	    RECT 121.4000 47.1000 121.8000 47.2000 ;
	    RECT 137.4000 47.1000 137.8000 47.2000 ;
	    RECT 121.4000 46.8000 137.8000 47.1000 ;
	    RECT 22.2000 46.2000 22.5000 46.8000 ;
	    RECT 22.2000 45.8000 22.6000 46.2000 ;
	    RECT 84.6000 46.1000 85.0000 46.2000 ;
	    RECT 88.6000 46.1000 89.0000 46.2000 ;
	    RECT 95.8000 46.1000 96.2000 46.2000 ;
	    RECT 84.6000 45.8000 96.2000 46.1000 ;
         LAYER metal4 ;
	    RECT 1.4000 48.8000 1.8000 49.2000 ;
	    RECT 1.4000 46.2000 1.7000 48.8000 ;
	    RECT 95.8000 47.8000 96.2000 48.2000 ;
	    RECT 22.2000 46.8000 22.6000 47.2000 ;
	    RECT 22.2000 46.2000 22.5000 46.8000 ;
	    RECT 95.8000 46.2000 96.1000 47.8000 ;
	    RECT 1.4000 45.8000 1.8000 46.2000 ;
	    RECT 22.2000 45.8000 22.6000 46.2000 ;
	    RECT 83.8000 46.1000 84.2000 46.2000 ;
	    RECT 84.6000 46.1000 85.0000 46.2000 ;
	    RECT 83.8000 45.8000 85.0000 46.1000 ;
	    RECT 95.8000 45.8000 96.2000 46.2000 ;
         LAYER metal5 ;
	    RECT 1.4000 46.1000 1.8000 46.2000 ;
	    RECT 22.2000 46.1000 22.6000 46.2000 ;
	    RECT 83.8000 46.1000 84.2000 46.2000 ;
	    RECT 1.4000 45.8000 84.2000 46.1000 ;
      END
   END DATA_B[10]
   PIN DATA_B[9]
      PORT
         LAYER metal1 ;
	    RECT 59.8000 12.4000 60.2000 13.2000 ;
	    RECT 156.6000 12.4000 157.0000 13.2000 ;
	    RECT 49.4000 7.8000 49.8000 8.6000 ;
	    RECT 119.0000 7.8000 119.4000 8.6000 ;
         LAYER metal2 ;
	    RECT 59.8000 12.8000 60.2000 13.2000 ;
	    RECT 156.6000 12.8000 157.0000 13.2000 ;
	    RECT 59.8000 12.2000 60.1000 12.8000 ;
	    RECT 156.6000 12.2000 156.9000 12.8000 ;
	    RECT 49.4000 11.8000 49.8000 12.2000 ;
	    RECT 59.8000 11.8000 60.2000 12.2000 ;
	    RECT 119.0000 11.8000 119.4000 12.2000 ;
	    RECT 156.6000 11.8000 157.0000 12.2000 ;
	    RECT 49.4000 8.2000 49.7000 11.8000 ;
	    RECT 119.0000 8.2000 119.3000 11.8000 ;
	    RECT 49.4000 7.8000 49.8000 8.2000 ;
	    RECT 119.0000 7.8000 119.4000 8.2000 ;
	    RECT 119.0000 -1.9000 119.3000 7.8000 ;
	    RECT 119.8000 -1.9000 120.2000 -1.8000 ;
	    RECT 119.0000 -2.2000 120.2000 -1.9000 ;
         LAYER metal3 ;
	    RECT 49.4000 12.1000 49.8000 12.2000 ;
	    RECT 59.8000 12.1000 60.2000 12.2000 ;
	    RECT 70.2000 12.1000 70.6000 12.2000 ;
	    RECT 49.4000 11.8000 70.6000 12.1000 ;
	    RECT 107.0000 12.1000 107.4000 12.2000 ;
	    RECT 119.0000 12.1000 119.4000 12.2000 ;
	    RECT 123.0000 12.1000 123.4000 12.2000 ;
	    RECT 107.0000 11.8000 123.4000 12.1000 ;
	    RECT 151.0000 12.1000 151.4000 12.2000 ;
	    RECT 156.6000 12.1000 157.0000 12.2000 ;
	    RECT 151.0000 11.8000 157.0000 12.1000 ;
         LAYER metal4 ;
	    RECT 70.2000 11.8000 70.6000 12.2000 ;
	    RECT 107.0000 11.8000 107.4000 12.2000 ;
	    RECT 123.0000 12.1000 123.4000 12.2000 ;
	    RECT 123.8000 12.1000 124.2000 12.2000 ;
	    RECT 123.0000 11.8000 124.2000 12.1000 ;
	    RECT 150.2000 12.1000 150.6000 12.2000 ;
	    RECT 151.0000 12.1000 151.4000 12.2000 ;
	    RECT 150.2000 11.8000 151.4000 12.1000 ;
	    RECT 70.2000 11.2000 70.5000 11.8000 ;
	    RECT 107.0000 11.2000 107.3000 11.8000 ;
	    RECT 70.2000 10.8000 70.6000 11.2000 ;
	    RECT 107.0000 10.8000 107.4000 11.2000 ;
         LAYER metal5 ;
	    RECT 123.8000 12.1000 124.2000 12.2000 ;
	    RECT 150.2000 12.1000 150.6000 12.2000 ;
	    RECT 123.8000 11.8000 150.6000 12.1000 ;
	    RECT 70.2000 11.1000 70.6000 11.2000 ;
	    RECT 107.0000 11.1000 107.4000 11.2000 ;
	    RECT 70.2000 10.8000 107.4000 11.1000 ;
      END
   END DATA_B[9]
   PIN DATA_B[8]
      PORT
         LAYER metal1 ;
	    RECT 158.2000 52.4000 158.6000 53.2000 ;
	    RECT 111.0000 47.8000 111.4000 48.6000 ;
	    RECT 43.0000 32.4000 43.4000 33.2000 ;
	    RECT 79.8000 32.4000 80.2000 33.2000 ;
         LAYER metal2 ;
	    RECT 157.4000 53.1000 157.8000 53.2000 ;
	    RECT 158.2000 53.1000 158.6000 53.2000 ;
	    RECT 157.4000 52.8000 158.6000 53.1000 ;
	    RECT 111.0000 47.8000 111.4000 48.2000 ;
	    RECT 111.0000 43.2000 111.3000 47.8000 ;
	    RECT 111.0000 42.8000 111.4000 43.2000 ;
	    RECT 111.0000 42.2000 111.3000 42.8000 ;
	    RECT 43.0000 41.8000 43.4000 42.2000 ;
	    RECT 79.8000 41.8000 80.2000 42.2000 ;
	    RECT 111.0000 41.8000 111.4000 42.2000 ;
	    RECT 43.0000 33.2000 43.3000 41.8000 ;
	    RECT 79.8000 33.2000 80.1000 41.8000 ;
	    RECT 43.0000 32.8000 43.4000 33.2000 ;
	    RECT 79.8000 32.8000 80.2000 33.2000 ;
         LAYER metal3 ;
	    RECT 158.2000 57.1000 158.6000 57.2000 ;
	    RECT 175.8000 57.1000 176.2000 57.2000 ;
	    RECT 158.2000 56.8000 176.2000 57.1000 ;
	    RECT 157.4000 53.1000 157.8000 53.2000 ;
	    RECT 158.2000 53.1000 158.6000 53.2000 ;
	    RECT 157.4000 52.8000 158.6000 53.1000 ;
	    RECT 111.0000 43.1000 111.4000 43.2000 ;
	    RECT 158.2000 43.1000 158.6000 43.2000 ;
	    RECT 111.0000 42.8000 158.6000 43.1000 ;
	    RECT 43.0000 42.1000 43.4000 42.2000 ;
	    RECT 79.8000 42.1000 80.2000 42.2000 ;
	    RECT 111.0000 42.1000 111.4000 42.2000 ;
	    RECT 43.0000 41.8000 111.4000 42.1000 ;
         LAYER metal4 ;
	    RECT 158.2000 56.8000 158.6000 57.2000 ;
	    RECT 158.2000 53.2000 158.5000 56.8000 ;
	    RECT 158.2000 52.8000 158.6000 53.2000 ;
	    RECT 158.2000 43.2000 158.5000 52.8000 ;
	    RECT 158.2000 42.8000 158.6000 43.2000 ;
      END
   END DATA_B[8]
   PIN DATA_B[7]
      PORT
         LAYER metal1 ;
	    RECT 62.2000 46.8000 62.7000 47.2000 ;
	    RECT 135.8000 46.8000 136.3000 47.2000 ;
	    RECT 153.4000 47.1000 153.8000 47.2000 ;
	    RECT 154.2000 47.1000 154.7000 47.2000 ;
	    RECT 153.4000 46.8000 154.7000 47.1000 ;
	    RECT 62.4000 46.4000 62.8000 46.8000 ;
	    RECT 136.0000 46.4000 136.4000 46.8000 ;
	    RECT 154.4000 46.4000 154.8000 46.8000 ;
	    RECT 26.8000 34.2000 27.2000 34.6000 ;
	    RECT 26.9000 34.1000 27.4000 34.2000 ;
	    RECT 27.8000 34.1000 28.2000 34.2000 ;
	    RECT 26.9000 33.8000 28.2000 34.1000 ;
         LAYER metal2 ;
	    RECT 62.2000 46.8000 62.6000 47.2000 ;
	    RECT 135.8000 46.8000 136.2000 47.2000 ;
	    RECT 153.4000 46.8000 153.8000 47.2000 ;
	    RECT 62.2000 39.2000 62.5000 46.8000 ;
	    RECT 135.8000 39.2000 136.1000 46.8000 ;
	    RECT 153.4000 46.2000 153.7000 46.8000 ;
	    RECT 153.4000 45.8000 153.8000 46.2000 ;
	    RECT 153.4000 39.2000 153.7000 45.8000 ;
	    RECT 27.8000 38.8000 28.2000 39.2000 ;
	    RECT 62.2000 38.8000 62.6000 39.2000 ;
	    RECT 135.8000 38.8000 136.2000 39.2000 ;
	    RECT 153.4000 38.8000 153.8000 39.2000 ;
	    RECT 27.8000 34.2000 28.1000 38.8000 ;
	    RECT 27.8000 33.8000 28.2000 34.2000 ;
         LAYER metal3 ;
	    RECT 155.0000 51.1000 155.4000 51.2000 ;
	    RECT 175.8000 51.1000 176.2000 51.2000 ;
	    RECT 155.0000 50.8000 176.2000 51.1000 ;
	    RECT 153.4000 46.1000 153.8000 46.2000 ;
	    RECT 155.0000 46.1000 155.4000 46.2000 ;
	    RECT 153.4000 45.8000 155.4000 46.1000 ;
	    RECT 27.8000 39.1000 28.2000 39.2000 ;
	    RECT 62.2000 39.1000 62.6000 39.2000 ;
	    RECT 135.8000 39.1000 136.2000 39.2000 ;
	    RECT 153.4000 39.1000 153.8000 39.2000 ;
	    RECT 27.8000 38.8000 153.8000 39.1000 ;
         LAYER metal4 ;
	    RECT 155.0000 50.8000 155.4000 51.2000 ;
	    RECT 155.0000 46.2000 155.3000 50.8000 ;
	    RECT 155.0000 45.8000 155.4000 46.2000 ;
      END
   END DATA_B[7]
   PIN DATA_B[6]
      PORT
         LAYER metal1 ;
	    RECT 26.9000 26.8000 27.4000 27.2000 ;
	    RECT 85.4000 26.8000 85.9000 27.2000 ;
	    RECT 26.8000 26.4000 27.2000 26.8000 ;
	    RECT 85.6000 26.4000 86.0000 26.8000 ;
	    RECT 95.6000 14.2000 96.0000 14.6000 ;
	    RECT 151.6000 14.2000 152.0000 14.6000 ;
	    RECT 95.7000 13.8000 96.2000 14.2000 ;
	    RECT 151.7000 13.8000 152.2000 14.2000 ;
         LAYER metal2 ;
	    RECT 27.0000 27.1000 27.4000 27.2000 ;
	    RECT 27.8000 27.1000 28.2000 27.2000 ;
	    RECT 27.0000 26.8000 28.2000 27.1000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 85.4000 26.8000 86.5000 27.1000 ;
	    RECT 86.2000 20.2000 86.5000 26.8000 ;
	    RECT 86.2000 19.8000 86.6000 20.2000 ;
	    RECT 95.8000 19.8000 96.2000 20.2000 ;
	    RECT 95.8000 14.2000 96.1000 19.8000 ;
	    RECT 151.8000 18.8000 152.2000 19.2000 ;
	    RECT 151.8000 14.2000 152.1000 18.8000 ;
	    RECT 95.8000 13.8000 96.2000 14.2000 ;
	    RECT 151.8000 13.8000 152.2000 14.2000 ;
	    RECT 98.2000 0.8000 98.6000 1.2000 ;
	    RECT 98.2000 -1.8000 98.5000 0.8000 ;
	    RECT 98.2000 -2.2000 98.6000 -1.8000 ;
         LAYER metal3 ;
	    RECT 27.0000 27.1000 27.4000 27.2000 ;
	    RECT 27.8000 27.1000 28.2000 27.2000 ;
	    RECT 27.0000 26.8000 28.2000 27.1000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 86.2000 27.1000 86.6000 27.2000 ;
	    RECT 85.4000 26.8000 86.6000 27.1000 ;
	    RECT 86.2000 20.1000 86.6000 20.2000 ;
	    RECT 95.8000 20.1000 96.2000 20.2000 ;
	    RECT 97.4000 20.1000 97.8000 20.2000 ;
	    RECT 86.2000 19.8000 132.1000 20.1000 ;
	    RECT 131.8000 19.1000 132.1000 19.8000 ;
	    RECT 151.8000 19.1000 152.2000 19.2000 ;
	    RECT 131.8000 18.8000 152.2000 19.1000 ;
	    RECT 97.4000 1.1000 97.8000 1.2000 ;
	    RECT 98.2000 1.1000 98.6000 1.2000 ;
	    RECT 97.4000 0.8000 98.6000 1.1000 ;
         LAYER metal4 ;
	    RECT 27.0000 27.1000 27.4000 27.2000 ;
	    RECT 27.8000 27.1000 28.2000 27.2000 ;
	    RECT 27.0000 26.8000 28.2000 27.1000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 86.2000 27.1000 86.6000 27.2000 ;
	    RECT 85.4000 26.8000 86.6000 27.1000 ;
	    RECT 97.4000 19.8000 97.8000 20.2000 ;
	    RECT 97.4000 1.2000 97.7000 19.8000 ;
	    RECT 97.4000 0.8000 97.8000 1.2000 ;
         LAYER metal5 ;
	    RECT 27.8000 27.1000 28.2000 27.2000 ;
	    RECT 85.4000 27.1000 85.8000 27.2000 ;
	    RECT 27.8000 26.8000 85.8000 27.1000 ;
      END
   END DATA_B[6]
   PIN DATA_B[5]
      PORT
         LAYER metal1 ;
	    RECT 42.8000 14.2000 43.2000 14.6000 ;
	    RECT 79.2000 14.2000 79.6000 14.6000 ;
	    RECT 132.4000 14.2000 132.8000 14.6000 ;
	    RECT 42.9000 14.1000 43.4000 14.2000 ;
	    RECT 43.8000 14.1000 44.2000 14.2000 ;
	    RECT 42.9000 13.8000 44.2000 14.1000 ;
	    RECT 79.0000 13.8000 79.5000 14.2000 ;
	    RECT 132.5000 13.8000 133.0000 14.2000 ;
	    RECT 152.6000 6.8000 153.1000 7.2000 ;
	    RECT 152.8000 6.4000 153.2000 6.8000 ;
         LAYER metal2 ;
	    RECT 43.0000 14.1000 43.4000 14.2000 ;
	    RECT 43.8000 14.1000 44.2000 14.2000 ;
	    RECT 43.0000 13.8000 44.2000 14.1000 ;
	    RECT 79.0000 13.8000 79.4000 14.2000 ;
	    RECT 132.6000 13.8000 133.0000 14.2000 ;
	    RECT 79.0000 13.2000 79.3000 13.8000 ;
	    RECT 132.6000 13.2000 132.9000 13.8000 ;
	    RECT 79.0000 12.8000 79.4000 13.2000 ;
	    RECT 132.6000 12.8000 133.0000 13.2000 ;
	    RECT 132.6000 8.2000 132.9000 12.8000 ;
	    RECT 132.6000 7.8000 133.0000 8.2000 ;
	    RECT 152.6000 7.8000 153.0000 8.2000 ;
	    RECT 152.6000 7.2000 152.9000 7.8000 ;
	    RECT 152.6000 6.8000 153.0000 7.2000 ;
	    RECT 152.6000 -1.8000 152.9000 6.8000 ;
	    RECT 152.6000 -2.2000 153.0000 -1.8000 ;
         LAYER metal3 ;
	    RECT 43.0000 14.1000 43.4000 14.2000 ;
	    RECT 43.8000 14.1000 44.2000 14.2000 ;
	    RECT 43.0000 13.8000 44.2000 14.1000 ;
	    RECT 76.6000 13.1000 77.0000 13.2000 ;
	    RECT 79.0000 13.1000 79.4000 13.2000 ;
	    RECT 76.6000 12.8000 79.4000 13.1000 ;
	    RECT 131.8000 13.1000 132.2000 13.2000 ;
	    RECT 132.6000 13.1000 133.0000 13.2000 ;
	    RECT 131.8000 12.8000 133.0000 13.1000 ;
	    RECT 132.6000 8.1000 133.0000 8.2000 ;
	    RECT 152.6000 8.1000 153.0000 8.2000 ;
	    RECT 132.6000 7.8000 153.0000 8.1000 ;
         LAYER metal4 ;
	    RECT 43.8000 13.8000 44.2000 14.2000 ;
	    RECT 43.8000 13.2000 44.1000 13.8000 ;
	    RECT 43.8000 12.8000 44.2000 13.2000 ;
	    RECT 75.8000 13.1000 76.2000 13.2000 ;
	    RECT 76.6000 13.1000 77.0000 13.2000 ;
	    RECT 75.8000 12.8000 77.0000 13.1000 ;
	    RECT 131.8000 13.1000 132.2000 13.2000 ;
	    RECT 132.6000 13.1000 133.0000 13.2000 ;
	    RECT 131.8000 12.8000 133.0000 13.1000 ;
         LAYER metal5 ;
	    RECT 43.8000 13.1000 44.2000 13.2000 ;
	    RECT 75.8000 13.1000 76.2000 13.2000 ;
	    RECT 132.6000 13.1000 133.0000 13.2000 ;
	    RECT 43.8000 12.8000 133.0000 13.1000 ;
      END
   END DATA_B[5]
   PIN DATA_B[4]
      PORT
         LAYER metal1 ;
	    RECT 38.1000 27.1000 38.6000 27.2000 ;
	    RECT 39.0000 27.1000 39.4000 27.2000 ;
	    RECT 38.1000 26.8000 39.4000 27.1000 ;
	    RECT 128.6000 26.8000 129.1000 27.2000 ;
	    RECT 38.0000 26.4000 38.4000 26.8000 ;
	    RECT 128.8000 26.4000 129.2000 26.8000 ;
	    RECT 54.0000 14.2000 54.4000 14.6000 ;
	    RECT 117.2000 14.2000 117.6000 14.6000 ;
	    RECT 54.1000 13.8000 54.6000 14.2000 ;
	    RECT 117.3000 13.8000 117.8000 14.2000 ;
         LAYER metal2 ;
	    RECT 39.0000 26.8000 39.4000 27.2000 ;
	    RECT 128.6000 26.8000 129.0000 27.2000 ;
	    RECT 39.0000 16.2000 39.3000 26.8000 ;
	    RECT 128.6000 22.2000 128.9000 26.8000 ;
	    RECT 128.6000 21.8000 129.0000 22.2000 ;
	    RECT 39.0000 15.8000 39.4000 16.2000 ;
	    RECT 54.2000 15.8000 54.6000 16.2000 ;
	    RECT 54.2000 14.2000 54.5000 15.8000 ;
	    RECT 117.4000 14.8000 117.8000 15.2000 ;
	    RECT 117.4000 14.2000 117.7000 14.8000 ;
	    RECT 54.2000 13.8000 54.6000 14.2000 ;
	    RECT 117.4000 13.8000 117.8000 14.2000 ;
	    RECT 117.4000 1.2000 117.7000 13.8000 ;
	    RECT 117.4000 0.8000 117.8000 1.2000 ;
	    RECT 121.4000 0.8000 121.8000 1.2000 ;
	    RECT 121.4000 -1.9000 121.7000 0.8000 ;
	    RECT 122.2000 -1.9000 122.6000 -1.8000 ;
	    RECT 121.4000 -2.2000 122.6000 -1.9000 ;
         LAYER metal3 ;
	    RECT 117.4000 22.1000 117.8000 22.2000 ;
	    RECT 128.6000 22.1000 129.0000 22.2000 ;
	    RECT 117.4000 21.8000 129.0000 22.1000 ;
	    RECT 39.0000 16.1000 39.4000 16.2000 ;
	    RECT 54.2000 16.1000 54.6000 16.2000 ;
	    RECT 70.2000 16.1000 70.6000 16.2000 ;
	    RECT 39.0000 15.8000 70.6000 16.1000 ;
	    RECT 116.6000 15.1000 117.0000 15.2000 ;
	    RECT 117.4000 15.1000 117.8000 15.2000 ;
	    RECT 116.6000 14.8000 117.8000 15.1000 ;
	    RECT 117.4000 1.1000 117.8000 1.2000 ;
	    RECT 121.4000 1.1000 121.8000 1.2000 ;
	    RECT 117.4000 0.8000 121.8000 1.1000 ;
         LAYER metal4 ;
	    RECT 117.4000 21.8000 117.8000 22.2000 ;
	    RECT 70.2000 15.8000 70.6000 16.2000 ;
	    RECT 70.2000 15.2000 70.5000 15.8000 ;
	    RECT 117.4000 15.2000 117.7000 21.8000 ;
	    RECT 70.2000 14.8000 70.6000 15.2000 ;
	    RECT 116.6000 15.1000 117.0000 15.2000 ;
	    RECT 117.4000 15.1000 117.8000 15.2000 ;
	    RECT 116.6000 14.8000 117.8000 15.1000 ;
         LAYER metal5 ;
	    RECT 70.2000 15.1000 70.6000 15.2000 ;
	    RECT 117.4000 15.1000 117.8000 15.2000 ;
	    RECT 70.2000 14.8000 117.8000 15.1000 ;
      END
   END DATA_B[4]
   PIN DATA_B[3]
      PORT
         LAYER metal1 ;
	    RECT 71.0000 26.8000 71.5000 27.2000 ;
	    RECT 140.6000 26.8000 141.1000 27.2000 ;
	    RECT 71.2000 26.4000 71.6000 26.8000 ;
	    RECT 140.8000 26.4000 141.2000 26.8000 ;
	    RECT 36.4000 14.2000 36.8000 14.6000 ;
	    RECT 135.6000 14.2000 136.0000 14.6000 ;
	    RECT 36.5000 14.1000 37.0000 14.2000 ;
	    RECT 37.4000 14.1000 37.8000 14.2000 ;
	    RECT 36.5000 13.8000 37.8000 14.1000 ;
	    RECT 135.7000 13.8000 136.2000 14.2000 ;
         LAYER metal2 ;
	    RECT 71.0000 26.8000 71.4000 27.2000 ;
	    RECT 139.8000 27.1000 140.2000 27.2000 ;
	    RECT 140.6000 27.1000 141.0000 27.2000 ;
	    RECT 139.8000 26.8000 141.0000 27.1000 ;
	    RECT 71.0000 18.2000 71.3000 26.8000 ;
	    RECT 37.4000 17.8000 37.8000 18.2000 ;
	    RECT 71.0000 17.8000 71.4000 18.2000 ;
	    RECT 37.4000 14.2000 37.7000 17.8000 ;
	    RECT 37.4000 13.8000 37.8000 14.2000 ;
	    RECT 135.0000 14.1000 135.4000 14.2000 ;
	    RECT 135.8000 14.1000 136.2000 14.2000 ;
	    RECT 135.0000 13.8000 136.2000 14.1000 ;
	    RECT 132.6000 0.8000 133.0000 1.2000 ;
	    RECT 132.6000 -1.8000 132.9000 0.8000 ;
	    RECT 132.6000 -2.2000 133.0000 -1.8000 ;
         LAYER metal3 ;
	    RECT 135.8000 27.1000 136.2000 27.2000 ;
	    RECT 139.8000 27.1000 140.2000 27.2000 ;
	    RECT 135.8000 26.8000 140.2000 27.1000 ;
	    RECT 37.4000 18.1000 37.8000 18.2000 ;
	    RECT 71.0000 18.1000 71.4000 18.2000 ;
	    RECT 94.2000 18.1000 94.6000 18.2000 ;
	    RECT 37.4000 17.8000 94.6000 18.1000 ;
	    RECT 135.0000 14.1000 135.4000 14.2000 ;
	    RECT 135.8000 14.1000 136.2000 14.2000 ;
	    RECT 135.0000 13.8000 136.2000 14.1000 ;
	    RECT 132.6000 1.1000 133.0000 1.2000 ;
	    RECT 135.0000 1.1000 135.4000 1.2000 ;
	    RECT 132.6000 0.8000 135.4000 1.1000 ;
         LAYER metal4 ;
	    RECT 135.8000 26.8000 136.2000 27.2000 ;
	    RECT 94.2000 17.8000 94.6000 18.2000 ;
	    RECT 94.2000 14.2000 94.5000 17.8000 ;
	    RECT 135.8000 14.2000 136.1000 26.8000 ;
	    RECT 94.2000 13.8000 94.6000 14.2000 ;
	    RECT 135.0000 14.1000 135.4000 14.2000 ;
	    RECT 135.8000 14.1000 136.2000 14.2000 ;
	    RECT 135.0000 13.8000 136.2000 14.1000 ;
	    RECT 135.0000 1.2000 135.3000 13.8000 ;
	    RECT 135.0000 0.8000 135.4000 1.2000 ;
         LAYER metal5 ;
	    RECT 94.2000 14.1000 94.6000 14.2000 ;
	    RECT 135.0000 14.1000 135.4000 14.2000 ;
	    RECT 94.2000 13.8000 135.4000 14.1000 ;
      END
   END DATA_B[3]
   PIN DATA_B[2]
      PORT
         LAYER metal1 ;
	    RECT 53.4000 47.8000 53.8000 48.6000 ;
	    RECT 138.2000 47.8000 138.6000 48.6000 ;
	    RECT 103.0000 32.4000 103.4000 33.2000 ;
	    RECT 7.0000 27.8000 7.4000 28.6000 ;
         LAYER metal2 ;
	    RECT 53.4000 48.1000 53.8000 48.2000 ;
	    RECT 53.4000 47.8000 54.5000 48.1000 ;
	    RECT 54.2000 37.2000 54.5000 47.8000 ;
	    RECT 138.2000 47.8000 138.6000 48.2000 ;
	    RECT 138.2000 38.2000 138.5000 47.8000 ;
	    RECT 138.2000 37.8000 138.6000 38.2000 ;
	    RECT 54.2000 36.8000 54.6000 37.2000 ;
	    RECT 103.0000 36.8000 103.4000 37.2000 ;
	    RECT 103.0000 33.2000 103.3000 36.8000 ;
	    RECT 103.0000 32.8000 103.4000 33.2000 ;
	    RECT 7.0000 28.8000 7.4000 29.2000 ;
	    RECT 7.0000 28.2000 7.3000 28.8000 ;
	    RECT 7.0000 27.8000 7.4000 28.2000 ;
         LAYER metal3 ;
	    RECT 138.2000 38.1000 138.6000 38.2000 ;
	    RECT 125.4000 37.8000 138.6000 38.1000 ;
	    RECT 7.0000 37.1000 7.4000 37.2000 ;
	    RECT 54.2000 37.1000 54.6000 37.2000 ;
	    RECT 103.0000 37.1000 103.4000 37.2000 ;
	    RECT 125.4000 37.1000 125.7000 37.8000 ;
	    RECT 7.0000 36.8000 125.7000 37.1000 ;
	    RECT 7.0000 29.1000 7.4000 29.2000 ;
	    RECT 7.8000 29.1000 8.2000 29.2000 ;
	    RECT -2.6000 28.8000 8.2000 29.1000 ;
	    RECT -2.6000 28.2000 -2.3000 28.8000 ;
	    RECT -2.6000 27.8000 -2.2000 28.2000 ;
         LAYER metal4 ;
	    RECT 7.0000 36.8000 7.4000 37.2000 ;
	    RECT 7.0000 29.1000 7.3000 36.8000 ;
	    RECT 7.8000 29.1000 8.2000 29.2000 ;
	    RECT 7.0000 28.8000 8.2000 29.1000 ;
      END
   END DATA_B[2]
   PIN DATA_B[1]
      PORT
         LAYER metal1 ;
	    RECT 114.4000 34.2000 114.8000 34.6000 ;
	    RECT 130.4000 34.2000 130.8000 34.6000 ;
	    RECT 113.4000 34.1000 113.8000 34.2000 ;
	    RECT 114.2000 34.1000 114.7000 34.2000 ;
	    RECT 113.4000 33.8000 114.7000 34.1000 ;
	    RECT 130.2000 33.8000 130.7000 34.2000 ;
	    RECT 7.6000 14.2000 8.0000 14.6000 ;
	    RECT 71.2000 14.2000 71.6000 14.6000 ;
	    RECT 7.7000 13.8000 8.2000 14.2000 ;
	    RECT 71.0000 13.8000 71.5000 14.2000 ;
         LAYER metal2 ;
	    RECT 113.4000 33.8000 113.8000 34.2000 ;
	    RECT 130.2000 33.8000 130.6000 34.2000 ;
	    RECT 113.4000 23.2000 113.7000 33.8000 ;
	    RECT 130.2000 29.1000 130.5000 33.8000 ;
	    RECT 129.4000 28.8000 130.5000 29.1000 ;
	    RECT 129.4000 23.2000 129.7000 28.8000 ;
	    RECT 113.4000 22.8000 113.8000 23.2000 ;
	    RECT 129.4000 22.8000 129.8000 23.2000 ;
	    RECT 7.8000 19.8000 8.2000 20.2000 ;
	    RECT 7.8000 14.2000 8.1000 19.8000 ;
	    RECT 71.0000 15.8000 71.4000 16.2000 ;
	    RECT 71.0000 14.2000 71.3000 15.8000 ;
	    RECT 7.8000 13.8000 8.2000 14.2000 ;
	    RECT 71.0000 13.8000 71.4000 14.2000 ;
         LAYER metal3 ;
	    RECT 71.8000 23.1000 72.2000 23.2000 ;
	    RECT 113.4000 23.1000 113.8000 23.2000 ;
	    RECT 129.4000 23.1000 129.8000 23.2000 ;
	    RECT 71.8000 22.8000 129.8000 23.1000 ;
	    RECT 0.6000 20.1000 1.0000 20.2000 ;
	    RECT 7.8000 20.1000 8.2000 20.2000 ;
	    RECT 15.8000 20.1000 16.2000 20.2000 ;
	    RECT 0.6000 19.8000 16.2000 20.1000 ;
	    RECT -2.6000 18.1000 -2.2000 18.2000 ;
	    RECT 0.6000 18.1000 1.0000 18.2000 ;
	    RECT -2.6000 17.8000 1.0000 18.1000 ;
	    RECT 71.0000 16.1000 71.4000 16.2000 ;
	    RECT 71.8000 16.1000 72.2000 16.2000 ;
	    RECT 71.0000 15.8000 72.2000 16.1000 ;
         LAYER metal4 ;
	    RECT 71.8000 22.8000 72.2000 23.2000 ;
	    RECT 0.6000 19.8000 1.0000 20.2000 ;
	    RECT 15.8000 19.8000 16.2000 20.2000 ;
	    RECT 0.6000 18.2000 0.9000 19.8000 ;
	    RECT 0.6000 17.8000 1.0000 18.2000 ;
	    RECT 15.8000 16.2000 16.1000 19.8000 ;
	    RECT 71.8000 16.2000 72.1000 22.8000 ;
	    RECT 15.8000 15.8000 16.2000 16.2000 ;
	    RECT 71.0000 16.1000 71.4000 16.2000 ;
	    RECT 71.8000 16.1000 72.2000 16.2000 ;
	    RECT 71.0000 15.8000 72.2000 16.1000 ;
         LAYER metal5 ;
	    RECT 15.8000 16.1000 16.2000 16.2000 ;
	    RECT 71.0000 16.1000 71.4000 16.2000 ;
	    RECT 15.8000 15.8000 71.4000 16.1000 ;
      END
   END DATA_B[1]
   PIN DATA_B[0]
      PORT
         LAYER metal1 ;
	    RECT 33.2000 34.2000 33.6000 34.6000 ;
	    RECT 44.8000 34.2000 45.2000 34.6000 ;
	    RECT 92.0000 34.2000 92.4000 34.6000 ;
	    RECT 33.3000 33.8000 33.8000 34.2000 ;
	    RECT 44.6000 33.8000 45.1000 34.2000 ;
	    RECT 91.8000 33.8000 92.3000 34.2000 ;
	    RECT 169.4000 26.8000 169.9000 27.2000 ;
	    RECT 169.6000 26.4000 170.0000 26.8000 ;
         LAYER metal2 ;
	    RECT 33.4000 33.8000 33.8000 34.2000 ;
	    RECT 44.6000 33.8000 45.0000 34.2000 ;
	    RECT 91.8000 33.8000 92.2000 34.2000 ;
	    RECT 33.4000 32.2000 33.7000 33.8000 ;
	    RECT 44.6000 32.2000 44.9000 33.8000 ;
	    RECT 91.8000 32.2000 92.1000 33.8000 ;
	    RECT 33.4000 31.8000 33.8000 32.2000 ;
	    RECT 44.6000 31.8000 45.0000 32.2000 ;
	    RECT 91.8000 31.8000 92.2000 32.2000 ;
	    RECT 91.8000 31.2000 92.1000 31.8000 ;
	    RECT 91.8000 30.8000 92.2000 31.2000 ;
	    RECT 169.4000 30.8000 169.8000 31.2000 ;
	    RECT 169.4000 27.2000 169.7000 30.8000 ;
	    RECT 169.4000 26.8000 169.8000 27.2000 ;
         LAYER metal3 ;
	    RECT 33.4000 32.1000 33.8000 32.2000 ;
	    RECT 44.6000 32.1000 45.0000 32.2000 ;
	    RECT 33.4000 31.8000 45.0000 32.1000 ;
	    RECT 91.8000 32.1000 92.2000 32.2000 ;
	    RECT 91.8000 31.8000 131.3000 32.1000 ;
	    RECT 44.6000 31.1000 44.9000 31.8000 ;
	    RECT 91.8000 31.1000 92.2000 31.2000 ;
	    RECT 44.6000 30.8000 92.2000 31.1000 ;
	    RECT 131.0000 31.1000 131.3000 31.8000 ;
	    RECT 169.4000 31.1000 169.8000 31.2000 ;
	    RECT 131.0000 30.8000 169.8000 31.1000 ;
	    RECT 169.4000 27.1000 169.8000 27.2000 ;
	    RECT 175.8000 27.1000 176.2000 27.2000 ;
	    RECT 169.4000 26.8000 176.2000 27.1000 ;
      END
   END DATA_B[0]
   PIN DATA_OUT[3]
      PORT
         LAYER metal1 ;
	    RECT 169.4000 66.2000 169.8000 69.9000 ;
	    RECT 169.5000 65.1000 169.8000 66.2000 ;
	    RECT 169.4000 61.1000 169.8000 65.1000 ;
         LAYER metal2 ;
	    RECT 169.4000 69.8000 169.8000 70.2000 ;
	    RECT 169.4000 69.2000 169.7000 69.8000 ;
	    RECT 169.4000 68.8000 169.8000 69.2000 ;
         LAYER metal3 ;
	    RECT 169.4000 70.1000 169.8000 70.2000 ;
	    RECT 175.8000 70.1000 176.2000 70.2000 ;
	    RECT 169.4000 69.8000 176.2000 70.1000 ;
      END
   END DATA_OUT[3]
   PIN DATA_OUT[2]
      PORT
         LAYER metal1 ;
	    RECT 170.2000 86.2000 170.6000 89.9000 ;
	    RECT 170.3000 85.1000 170.6000 86.2000 ;
	    RECT 170.2000 81.1000 170.6000 85.1000 ;
         LAYER metal2 ;
	    RECT 170.2000 84.8000 170.6000 85.2000 ;
	    RECT 170.2000 84.2000 170.5000 84.8000 ;
	    RECT 170.2000 83.8000 170.6000 84.2000 ;
         LAYER metal3 ;
	    RECT 170.2000 85.1000 170.6000 85.2000 ;
	    RECT 175.8000 85.1000 176.2000 85.2000 ;
	    RECT 170.2000 84.8000 176.2000 85.1000 ;
      END
   END DATA_OUT[2]
   PIN DATA_OUT[1]
      PORT
         LAYER metal1 ;
	    RECT 171.8000 59.1000 172.2000 59.9000 ;
	    RECT 173.4000 59.1000 173.8000 59.2000 ;
	    RECT 171.8000 58.8000 173.8000 59.1000 ;
	    RECT 171.8000 55.9000 172.2000 58.8000 ;
	    RECT 171.9000 54.8000 172.2000 55.9000 ;
	    RECT 171.8000 51.1000 172.2000 54.8000 ;
         LAYER metal2 ;
	    RECT 173.4000 62.8000 173.8000 63.2000 ;
	    RECT 173.4000 59.2000 173.7000 62.8000 ;
	    RECT 173.4000 58.8000 173.8000 59.2000 ;
         LAYER metal3 ;
	    RECT 173.4000 63.1000 173.8000 63.2000 ;
	    RECT 175.8000 63.1000 176.2000 63.2000 ;
	    RECT 173.4000 62.8000 176.2000 63.1000 ;
      END
   END DATA_OUT[1]
   PIN DATA_OUT[0]
      PORT
         LAYER metal1 ;
	    RECT 171.8000 68.1000 172.2000 69.9000 ;
	    RECT 172.6000 68.1000 173.0000 68.2000 ;
	    RECT 171.8000 67.8000 173.0000 68.1000 ;
	    RECT 171.8000 66.2000 172.2000 67.8000 ;
	    RECT 171.9000 65.1000 172.2000 66.2000 ;
	    RECT 171.8000 61.1000 172.2000 65.1000 ;
         LAYER metal2 ;
	    RECT 172.6000 68.1000 173.0000 68.2000 ;
	    RECT 173.4000 68.1000 173.8000 68.2000 ;
	    RECT 172.6000 67.8000 173.8000 68.1000 ;
         LAYER metal3 ;
	    RECT 173.4000 68.1000 173.8000 68.2000 ;
	    RECT 175.8000 68.1000 176.2000 68.2000 ;
	    RECT 173.4000 67.8000 176.2000 68.1000 ;
      END
   END DATA_OUT[0]
   PIN RESET_L
      PORT
         LAYER metal1 ;
	    RECT 123.8000 125.8000 124.2000 126.6000 ;
	    RECT 140.6000 94.4000 141.0000 95.2000 ;
	    RECT 115.8000 85.8000 116.2000 86.6000 ;
	    RECT 111.8000 74.4000 112.2000 75.2000 ;
	    RECT 139.8000 74.4000 140.2000 75.2000 ;
         LAYER metal2 ;
	    RECT 123.0000 163.8000 123.4000 164.2000 ;
	    RECT 123.0000 161.2000 123.3000 163.8000 ;
	    RECT 123.0000 160.8000 123.4000 161.2000 ;
	    RECT 123.0000 126.1000 123.4000 126.2000 ;
	    RECT 123.8000 126.1000 124.2000 126.2000 ;
	    RECT 123.0000 125.8000 124.2000 126.1000 ;
	    RECT 139.8000 95.1000 140.2000 95.2000 ;
	    RECT 140.6000 95.1000 141.0000 95.2000 ;
	    RECT 139.8000 94.8000 141.0000 95.1000 ;
	    RECT 115.8000 85.8000 116.2000 86.2000 ;
	    RECT 115.8000 85.2000 116.1000 85.8000 ;
	    RECT 111.8000 84.8000 112.2000 85.2000 ;
	    RECT 115.8000 84.8000 116.2000 85.2000 ;
	    RECT 111.8000 77.2000 112.1000 84.8000 ;
	    RECT 111.8000 76.8000 112.2000 77.2000 ;
	    RECT 139.8000 76.8000 140.2000 77.2000 ;
	    RECT 111.8000 75.2000 112.1000 76.8000 ;
	    RECT 139.8000 75.2000 140.1000 76.8000 ;
	    RECT 111.8000 74.8000 112.2000 75.2000 ;
	    RECT 139.8000 74.8000 140.2000 75.2000 ;
         LAYER metal3 ;
	    RECT 123.0000 161.1000 123.4000 161.2000 ;
	    RECT 123.8000 161.1000 124.2000 161.2000 ;
	    RECT 123.0000 160.8000 124.2000 161.1000 ;
	    RECT 123.0000 126.1000 123.4000 126.2000 ;
	    RECT 123.8000 126.1000 124.2000 126.2000 ;
	    RECT 123.0000 125.8000 124.2000 126.1000 ;
	    RECT 139.8000 95.1000 140.2000 95.2000 ;
	    RECT 140.6000 95.1000 141.0000 95.2000 ;
	    RECT 139.8000 94.8000 141.0000 95.1000 ;
	    RECT 111.8000 85.1000 112.2000 85.2000 ;
	    RECT 115.8000 85.1000 116.2000 85.2000 ;
	    RECT 111.8000 84.8000 116.2000 85.1000 ;
	    RECT 139.8000 77.8000 140.2000 78.2000 ;
	    RECT 139.8000 77.2000 140.1000 77.8000 ;
	    RECT 111.8000 77.1000 112.2000 77.2000 ;
	    RECT 123.8000 77.1000 124.2000 77.2000 ;
	    RECT 139.8000 77.1000 140.2000 77.2000 ;
	    RECT 111.8000 76.8000 140.2000 77.1000 ;
         LAYER metal4 ;
	    RECT 123.8000 160.8000 124.2000 161.2000 ;
	    RECT 123.8000 126.2000 124.1000 160.8000 ;
	    RECT 123.8000 125.8000 124.2000 126.2000 ;
	    RECT 123.8000 77.2000 124.1000 125.8000 ;
	    RECT 140.6000 95.1000 141.0000 95.2000 ;
	    RECT 139.8000 94.8000 141.0000 95.1000 ;
	    RECT 139.8000 78.2000 140.1000 94.8000 ;
	    RECT 139.8000 77.8000 140.2000 78.2000 ;
	    RECT 123.8000 76.8000 124.2000 77.2000 ;
      END
   END RESET_L
   PIN SEL_A[11]
      PORT
         LAYER metal1 ;
	    RECT 18.2000 154.4000 18.6000 155.2000 ;
	    RECT 23.0000 135.1000 23.4000 135.2000 ;
	    RECT 23.8000 135.1000 24.2000 135.2000 ;
	    RECT 23.0000 134.8000 24.2000 135.1000 ;
	    RECT 23.8000 134.4000 24.2000 134.8000 ;
	    RECT 18.2000 114.4000 18.6000 115.2000 ;
	    RECT 19.0000 105.8000 19.4000 106.6000 ;
	    RECT 23.8000 94.4000 24.2000 95.2000 ;
         LAYER metal2 ;
	    RECT 19.8000 163.8000 20.2000 164.2000 ;
	    RECT 18.2000 155.1000 18.6000 155.2000 ;
	    RECT 19.0000 155.1000 19.4000 155.2000 ;
	    RECT 19.8000 155.1000 20.1000 163.8000 ;
	    RECT 18.2000 154.8000 20.1000 155.1000 ;
	    RECT 23.0000 134.8000 23.4000 135.2000 ;
	    RECT 23.0000 131.2000 23.3000 134.8000 ;
	    RECT 18.2000 130.8000 18.6000 131.2000 ;
	    RECT 23.0000 130.8000 23.4000 131.2000 ;
	    RECT 18.2000 115.2000 18.5000 130.8000 ;
	    RECT 18.2000 114.8000 18.6000 115.2000 ;
	    RECT 18.2000 103.1000 18.5000 114.8000 ;
	    RECT 19.0000 105.8000 19.4000 106.2000 ;
	    RECT 19.0000 103.2000 19.3000 105.8000 ;
	    RECT 19.0000 103.1000 19.4000 103.2000 ;
	    RECT 18.2000 102.8000 19.4000 103.1000 ;
	    RECT 23.8000 102.8000 24.2000 103.2000 ;
	    RECT 23.8000 95.2000 24.1000 102.8000 ;
	    RECT 23.8000 94.8000 24.2000 95.2000 ;
         LAYER metal3 ;
	    RECT 19.0000 154.8000 19.4000 155.2000 ;
	    RECT 19.0000 154.2000 19.3000 154.8000 ;
	    RECT 19.0000 153.8000 19.4000 154.2000 ;
	    RECT 18.2000 131.1000 18.6000 131.2000 ;
	    RECT 19.0000 131.1000 19.4000 131.2000 ;
	    RECT 23.0000 131.1000 23.4000 131.2000 ;
	    RECT 18.2000 130.8000 23.4000 131.1000 ;
	    RECT 19.0000 103.1000 19.4000 103.2000 ;
	    RECT 23.8000 103.1000 24.2000 103.2000 ;
	    RECT 19.0000 102.8000 24.2000 103.1000 ;
         LAYER metal4 ;
	    RECT 19.0000 153.8000 19.4000 154.2000 ;
	    RECT 19.0000 131.2000 19.3000 153.8000 ;
	    RECT 19.0000 130.8000 19.4000 131.2000 ;
      END
   END SEL_A[11]
   PIN SEL_A[10]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 133.4000 21.0000 134.2000 ;
	    RECT 30.2000 133.4000 30.6000 134.2000 ;
	    RECT 35.8000 133.4000 36.2000 134.2000 ;
	    RECT 7.8000 126.8000 8.2000 127.6000 ;
	    RECT 7.8000 126.2000 8.1000 126.8000 ;
	    RECT 7.8000 125.8000 8.2000 126.2000 ;
	    RECT 27.8000 115.4000 28.2000 116.2000 ;
	    RECT 10.2000 104.8000 10.6000 105.6000 ;
	    RECT 29.4000 95.4000 29.8000 96.2000 ;
	    RECT 38.2000 86.8000 38.6000 87.6000 ;
	    RECT 26.2000 84.8000 26.6000 85.6000 ;
         LAYER metal2 ;
	    RECT 20.6000 133.8000 21.0000 134.2000 ;
	    RECT 30.2000 133.8000 30.6000 134.2000 ;
	    RECT 35.8000 133.8000 36.2000 134.2000 ;
	    RECT 20.6000 133.2000 20.9000 133.8000 ;
	    RECT 30.2000 133.2000 30.5000 133.8000 ;
	    RECT 35.8000 133.2000 36.1000 133.8000 ;
	    RECT 20.6000 132.8000 21.0000 133.2000 ;
	    RECT 27.8000 132.8000 28.2000 133.2000 ;
	    RECT 30.2000 132.8000 30.6000 133.2000 ;
	    RECT 35.8000 132.8000 36.2000 133.2000 ;
	    RECT 20.6000 127.2000 20.9000 132.8000 ;
	    RECT 7.8000 126.8000 8.2000 127.2000 ;
	    RECT 20.6000 126.8000 21.0000 127.2000 ;
	    RECT 7.8000 126.2000 8.1000 126.8000 ;
	    RECT 7.8000 125.8000 8.2000 126.2000 ;
	    RECT 7.8000 110.2000 8.1000 125.8000 ;
	    RECT 27.8000 116.2000 28.1000 132.8000 ;
	    RECT 27.8000 115.8000 28.2000 116.2000 ;
	    RECT 7.8000 109.8000 8.2000 110.2000 ;
	    RECT 10.2000 109.8000 10.6000 110.2000 ;
	    RECT 10.2000 105.2000 10.5000 109.8000 ;
	    RECT 27.8000 109.2000 28.1000 115.8000 ;
	    RECT 27.8000 108.8000 28.2000 109.2000 ;
	    RECT 10.2000 104.8000 10.6000 105.2000 ;
	    RECT 29.4000 97.8000 29.8000 98.2000 ;
	    RECT 29.4000 96.2000 29.7000 97.8000 ;
	    RECT 29.4000 95.8000 29.8000 96.2000 ;
	    RECT 26.2000 86.8000 26.6000 87.2000 ;
	    RECT 37.4000 87.1000 37.8000 87.2000 ;
	    RECT 38.2000 87.1000 38.6000 87.2000 ;
	    RECT 37.4000 86.8000 38.6000 87.1000 ;
	    RECT 26.2000 85.2000 26.5000 86.8000 ;
	    RECT 26.2000 84.8000 26.6000 85.2000 ;
         LAYER metal3 ;
	    RECT 20.6000 133.1000 21.0000 133.2000 ;
	    RECT 27.8000 133.1000 28.2000 133.2000 ;
	    RECT 30.2000 133.1000 30.6000 133.2000 ;
	    RECT 35.8000 133.1000 36.2000 133.2000 ;
	    RECT 20.6000 132.8000 36.2000 133.1000 ;
	    RECT -2.6000 128.1000 -2.2000 128.2000 ;
	    RECT -2.6000 127.8000 -1.5000 128.1000 ;
	    RECT -1.8000 127.1000 -1.5000 127.8000 ;
	    RECT 7.8000 127.1000 8.2000 127.2000 ;
	    RECT 20.6000 127.1000 21.0000 127.2000 ;
	    RECT -1.8000 126.8000 21.0000 127.1000 ;
	    RECT 7.8000 110.1000 8.2000 110.2000 ;
	    RECT 10.2000 110.1000 10.6000 110.2000 ;
	    RECT 7.8000 109.8000 10.6000 110.1000 ;
	    RECT 27.8000 108.8000 28.2000 109.2000 ;
	    RECT 27.8000 108.2000 28.1000 108.8000 ;
	    RECT 27.8000 107.8000 28.2000 108.2000 ;
	    RECT 27.8000 98.1000 28.2000 98.2000 ;
	    RECT 29.4000 98.1000 29.8000 98.2000 ;
	    RECT 27.8000 97.8000 29.8000 98.1000 ;
	    RECT 26.2000 87.1000 26.6000 87.2000 ;
	    RECT 27.8000 87.1000 28.2000 87.2000 ;
	    RECT 37.4000 87.1000 37.8000 87.2000 ;
	    RECT 26.2000 86.8000 37.8000 87.1000 ;
         LAYER metal4 ;
	    RECT 27.8000 107.8000 28.2000 108.2000 ;
	    RECT 27.8000 98.2000 28.1000 107.8000 ;
	    RECT 27.8000 97.8000 28.2000 98.2000 ;
	    RECT 27.8000 87.2000 28.1000 97.8000 ;
	    RECT 27.8000 86.8000 28.2000 87.2000 ;
      END
   END SEL_A[10]
   PIN SEL_A[9]
      PORT
         LAYER metal1 ;
	    RECT 20.6000 124.8000 21.0000 125.6000 ;
	    RECT 33.4000 124.8000 33.8000 125.6000 ;
	    RECT 34.2000 115.4000 34.6000 116.2000 ;
	    RECT 27.0000 106.8000 27.4000 107.6000 ;
	    RECT 40.6000 84.8000 41.0000 85.6000 ;
         LAYER metal2 ;
	    RECT 0.6000 124.8000 1.0000 125.2000 ;
	    RECT 20.6000 125.1000 21.0000 125.2000 ;
	    RECT 21.4000 125.1000 21.8000 125.2000 ;
	    RECT 20.6000 124.8000 21.8000 125.1000 ;
	    RECT 33.4000 124.8000 33.8000 125.2000 ;
	    RECT 0.6000 123.2000 0.9000 124.8000 ;
	    RECT 20.6000 123.2000 20.9000 124.8000 ;
	    RECT 0.6000 122.8000 1.0000 123.2000 ;
	    RECT 20.6000 122.8000 21.0000 123.2000 ;
	    RECT 33.4000 119.2000 33.7000 124.8000 ;
	    RECT 33.4000 118.8000 33.8000 119.2000 ;
	    RECT 34.2000 115.8000 34.6000 116.2000 ;
	    RECT 34.2000 111.2000 34.5000 115.8000 ;
	    RECT 27.0000 110.8000 27.4000 111.2000 ;
	    RECT 34.2000 110.8000 34.6000 111.2000 ;
	    RECT 27.0000 107.2000 27.3000 110.8000 ;
	    RECT 27.0000 106.8000 27.4000 107.2000 ;
	    RECT 40.6000 95.8000 41.0000 96.2000 ;
	    RECT 40.6000 85.2000 40.9000 95.8000 ;
	    RECT 40.6000 84.8000 41.0000 85.2000 ;
         LAYER metal3 ;
	    RECT -2.6000 125.1000 -2.2000 125.2000 ;
	    RECT 0.6000 125.1000 1.0000 125.2000 ;
	    RECT -2.6000 124.8000 1.0000 125.1000 ;
	    RECT 21.4000 125.1000 21.8000 125.2000 ;
	    RECT 33.4000 125.1000 33.8000 125.2000 ;
	    RECT 21.4000 124.8000 33.8000 125.1000 ;
	    RECT 0.6000 123.1000 1.0000 123.2000 ;
	    RECT 20.6000 123.1000 21.0000 123.2000 ;
	    RECT 0.6000 122.8000 21.0000 123.1000 ;
	    RECT 33.4000 119.1000 33.8000 119.2000 ;
	    RECT 34.2000 119.1000 34.6000 119.2000 ;
	    RECT 33.4000 118.8000 34.6000 119.1000 ;
	    RECT 27.0000 111.1000 27.4000 111.2000 ;
	    RECT 33.4000 111.1000 33.8000 111.2000 ;
	    RECT 34.2000 111.1000 34.6000 111.2000 ;
	    RECT 27.0000 110.8000 34.6000 111.1000 ;
	    RECT 33.4000 96.1000 33.8000 96.2000 ;
	    RECT 40.6000 96.1000 41.0000 96.2000 ;
	    RECT 33.4000 95.8000 41.0000 96.1000 ;
         LAYER metal4 ;
	    RECT 34.2000 119.1000 34.6000 119.2000 ;
	    RECT 33.4000 118.8000 34.6000 119.1000 ;
	    RECT 33.4000 111.2000 33.7000 118.8000 ;
	    RECT 33.4000 110.8000 33.8000 111.2000 ;
	    RECT 33.4000 96.2000 33.7000 110.8000 ;
	    RECT 33.4000 95.8000 33.8000 96.2000 ;
      END
   END SEL_A[9]
   PIN SEL_A[8]
      PORT
         LAYER metal1 ;
	    RECT 41.4000 145.8000 41.8000 146.6000 ;
	    RECT 58.2000 125.8000 58.6000 126.6000 ;
	    RECT 63.8000 85.8000 64.2000 86.6000 ;
	    RECT 56.6000 74.4000 57.0000 75.2000 ;
	    RECT 65.4000 74.4000 65.8000 75.2000 ;
         LAYER metal2 ;
	    RECT 41.4000 163.8000 41.8000 164.2000 ;
	    RECT 41.4000 146.2000 41.7000 163.8000 ;
	    RECT 41.4000 146.1000 41.8000 146.2000 ;
	    RECT 41.4000 145.8000 42.5000 146.1000 ;
	    RECT 42.2000 122.2000 42.5000 145.8000 ;
	    RECT 58.2000 125.8000 58.6000 126.2000 ;
	    RECT 58.2000 122.2000 58.5000 125.8000 ;
	    RECT 42.2000 121.8000 42.6000 122.2000 ;
	    RECT 58.2000 121.8000 58.6000 122.2000 ;
	    RECT 63.8000 85.8000 64.2000 86.2000 ;
	    RECT 63.8000 83.2000 64.1000 85.8000 ;
	    RECT 63.8000 82.8000 64.2000 83.2000 ;
	    RECT 65.4000 82.8000 65.8000 83.2000 ;
	    RECT 65.4000 75.2000 65.7000 82.8000 ;
	    RECT 56.6000 75.1000 57.0000 75.2000 ;
	    RECT 57.4000 75.1000 57.8000 75.2000 ;
	    RECT 56.6000 74.8000 57.8000 75.1000 ;
	    RECT 65.4000 75.1000 65.8000 75.2000 ;
	    RECT 66.2000 75.1000 66.6000 75.2000 ;
	    RECT 65.4000 74.8000 66.6000 75.1000 ;
         LAYER metal3 ;
	    RECT 42.2000 122.1000 42.6000 122.2000 ;
	    RECT 58.2000 122.1000 58.6000 122.2000 ;
	    RECT 59.0000 122.1000 59.4000 122.2000 ;
	    RECT 42.2000 121.8000 59.4000 122.1000 ;
	    RECT 59.0000 83.1000 59.4000 83.2000 ;
	    RECT 63.8000 83.1000 64.2000 83.2000 ;
	    RECT 65.4000 83.1000 65.8000 83.2000 ;
	    RECT 59.0000 82.8000 65.8000 83.1000 ;
	    RECT 57.4000 75.1000 57.8000 75.2000 ;
	    RECT 66.2000 75.1000 66.6000 75.2000 ;
	    RECT 57.4000 74.8000 66.6000 75.1000 ;
         LAYER metal4 ;
	    RECT 59.0000 121.8000 59.4000 122.2000 ;
	    RECT 59.0000 83.2000 59.3000 121.8000 ;
	    RECT 59.0000 82.8000 59.4000 83.2000 ;
      END
   END SEL_A[8]
   PIN SEL_A[7]
      PORT
         LAYER metal1 ;
	    RECT 59.8000 133.4000 60.2000 134.2000 ;
	    RECT 63.8000 133.4000 64.2000 134.2000 ;
	    RECT 69.4000 133.4000 69.8000 134.2000 ;
	    RECT 71.8000 106.8000 72.2000 107.6000 ;
	    RECT 72.6000 95.4000 73.0000 96.2000 ;
	    RECT 59.8000 76.1000 60.2000 76.2000 ;
	    RECT 60.6000 76.1000 61.0000 76.2000 ;
	    RECT 59.8000 75.8000 61.0000 76.1000 ;
	    RECT 59.8000 75.4000 60.2000 75.8000 ;
	    RECT 73.4000 75.4000 73.8000 76.2000 ;
	    RECT 80.6000 75.4000 81.0000 76.2000 ;
	    RECT 59.8000 67.1000 60.2000 67.6000 ;
	    RECT 60.6000 67.1000 61.0000 67.2000 ;
	    RECT 59.8000 66.8000 61.0000 67.1000 ;
         LAYER metal2 ;
	    RECT 69.4000 163.8000 69.8000 164.2000 ;
	    RECT 69.4000 161.2000 69.7000 163.8000 ;
	    RECT 69.4000 160.8000 69.8000 161.2000 ;
	    RECT 59.8000 134.1000 60.2000 134.2000 ;
	    RECT 60.6000 134.1000 61.0000 134.2000 ;
	    RECT 59.8000 133.8000 61.0000 134.1000 ;
	    RECT 63.8000 134.1000 64.2000 134.2000 ;
	    RECT 64.6000 134.1000 65.0000 134.2000 ;
	    RECT 63.8000 133.8000 65.0000 134.1000 ;
	    RECT 69.4000 133.8000 69.8000 134.2000 ;
	    RECT 69.4000 125.1000 69.7000 133.8000 ;
	    RECT 69.4000 124.8000 70.5000 125.1000 ;
	    RECT 70.2000 118.2000 70.5000 124.8000 ;
	    RECT 70.2000 117.8000 70.6000 118.2000 ;
	    RECT 71.8000 117.8000 72.2000 118.2000 ;
	    RECT 71.8000 107.2000 72.1000 117.8000 ;
	    RECT 71.8000 106.8000 72.2000 107.2000 ;
	    RECT 71.8000 99.1000 72.1000 106.8000 ;
	    RECT 71.8000 98.8000 72.9000 99.1000 ;
	    RECT 72.6000 96.2000 72.9000 98.8000 ;
	    RECT 72.6000 95.8000 73.0000 96.2000 ;
	    RECT 72.6000 91.2000 72.9000 95.8000 ;
	    RECT 72.6000 90.8000 73.0000 91.2000 ;
	    RECT 80.6000 90.8000 81.0000 91.2000 ;
	    RECT 80.6000 76.2000 80.9000 90.8000 ;
	    RECT 60.6000 76.1000 61.0000 76.2000 ;
	    RECT 61.4000 76.1000 61.8000 76.2000 ;
	    RECT 60.6000 75.8000 61.8000 76.1000 ;
	    RECT 73.4000 76.1000 73.8000 76.2000 ;
	    RECT 74.2000 76.1000 74.6000 76.2000 ;
	    RECT 73.4000 75.8000 74.6000 76.1000 ;
	    RECT 80.6000 75.8000 81.0000 76.2000 ;
	    RECT 60.6000 67.2000 60.9000 75.8000 ;
	    RECT 60.6000 66.8000 61.0000 67.2000 ;
         LAYER metal3 ;
	    RECT 69.4000 160.8000 69.8000 161.2000 ;
	    RECT 69.4000 160.2000 69.7000 160.8000 ;
	    RECT 69.4000 159.8000 69.8000 160.2000 ;
	    RECT 60.6000 134.1000 61.0000 134.2000 ;
	    RECT 64.6000 134.1000 65.0000 134.2000 ;
	    RECT 69.4000 134.1000 69.8000 134.2000 ;
	    RECT 60.6000 133.8000 69.8000 134.1000 ;
	    RECT 70.2000 118.1000 70.6000 118.2000 ;
	    RECT 71.8000 118.1000 72.2000 118.2000 ;
	    RECT 70.2000 117.8000 72.2000 118.1000 ;
	    RECT 72.6000 91.1000 73.0000 91.2000 ;
	    RECT 80.6000 91.1000 81.0000 91.2000 ;
	    RECT 72.6000 90.8000 81.0000 91.1000 ;
	    RECT 61.4000 76.1000 61.8000 76.2000 ;
	    RECT 74.2000 76.1000 74.6000 76.2000 ;
	    RECT 80.6000 76.1000 81.0000 76.2000 ;
	    RECT 61.4000 75.8000 81.0000 76.1000 ;
         LAYER metal4 ;
	    RECT 69.4000 159.8000 69.8000 160.2000 ;
	    RECT 69.4000 134.2000 69.7000 159.8000 ;
	    RECT 69.4000 133.8000 69.8000 134.2000 ;
      END
   END SEL_A[7]
   PIN SEL_A[6]
      PORT
         LAYER metal1 ;
	    RECT 63.0000 124.8000 63.4000 125.6000 ;
	    RECT 67.8000 115.4000 68.2000 116.2000 ;
	    RECT 71.0000 115.4000 71.4000 116.2000 ;
	    RECT 73.4000 107.1000 73.8000 107.2000 ;
	    RECT 74.2000 107.1000 74.6000 107.6000 ;
	    RECT 73.4000 106.8000 74.6000 107.1000 ;
	    RECT 64.6000 75.4000 65.0000 76.2000 ;
         LAYER metal2 ;
	    RECT 67.0000 163.8000 67.4000 164.2000 ;
	    RECT 67.0000 158.2000 67.3000 163.8000 ;
	    RECT 67.0000 157.8000 67.4000 158.2000 ;
	    RECT 63.0000 124.8000 63.4000 125.2000 ;
	    RECT 63.0000 116.2000 63.3000 124.8000 ;
	    RECT 63.0000 115.8000 63.4000 116.2000 ;
	    RECT 67.8000 116.1000 68.2000 116.2000 ;
	    RECT 68.6000 116.1000 69.0000 116.2000 ;
	    RECT 67.8000 115.8000 69.0000 116.1000 ;
	    RECT 71.0000 115.8000 71.4000 116.2000 ;
	    RECT 73.4000 115.8000 73.8000 116.2000 ;
	    RECT 71.0000 115.2000 71.3000 115.8000 ;
	    RECT 71.0000 114.8000 71.4000 115.2000 ;
	    RECT 73.4000 107.2000 73.7000 115.8000 ;
	    RECT 73.4000 106.8000 73.8000 107.2000 ;
	    RECT 64.6000 76.8000 65.0000 77.2000 ;
	    RECT 64.6000 76.2000 64.9000 76.8000 ;
	    RECT 64.6000 75.8000 65.0000 76.2000 ;
         LAYER metal3 ;
	    RECT 67.0000 158.1000 67.4000 158.2000 ;
	    RECT 67.8000 158.1000 68.2000 158.2000 ;
	    RECT 67.0000 157.8000 68.2000 158.1000 ;
	    RECT 63.0000 116.1000 63.4000 116.2000 ;
	    RECT 65.4000 116.1000 65.8000 116.2000 ;
	    RECT 67.0000 116.1000 67.4000 116.2000 ;
	    RECT 68.6000 116.1000 69.0000 116.2000 ;
	    RECT 73.4000 116.1000 73.8000 116.2000 ;
	    RECT 63.0000 115.8000 73.8000 116.1000 ;
	    RECT 71.0000 115.2000 71.3000 115.8000 ;
	    RECT 71.0000 114.8000 71.4000 115.2000 ;
	    RECT 64.6000 77.1000 65.0000 77.2000 ;
	    RECT 65.4000 77.1000 65.8000 77.2000 ;
	    RECT 64.6000 76.8000 65.8000 77.1000 ;
         LAYER metal4 ;
	    RECT 67.8000 158.1000 68.2000 158.2000 ;
	    RECT 67.0000 157.8000 68.2000 158.1000 ;
	    RECT 67.0000 116.2000 67.3000 157.8000 ;
	    RECT 65.4000 115.8000 65.8000 116.2000 ;
	    RECT 67.0000 115.8000 67.4000 116.2000 ;
	    RECT 65.4000 77.2000 65.7000 115.8000 ;
	    RECT 65.4000 76.8000 65.8000 77.2000 ;
      END
   END SEL_A[6]
   PIN SEL_A[5]
      PORT
         LAYER metal1 ;
	    RECT 11.8000 145.8000 12.2000 146.6000 ;
	    RECT 0.6000 134.4000 1.0000 135.2000 ;
	    RECT 0.6000 94.4000 1.0000 95.2000 ;
	    RECT 6.2000 74.4000 6.6000 75.2000 ;
	    RECT 8.6000 74.4000 9.0000 75.2000 ;
         LAYER metal2 ;
	    RECT 11.8000 145.8000 12.2000 146.2000 ;
	    RECT 11.8000 145.2000 12.1000 145.8000 ;
	    RECT 0.6000 144.8000 1.0000 145.2000 ;
	    RECT 11.8000 144.8000 12.2000 145.2000 ;
	    RECT 0.6000 135.2000 0.9000 144.8000 ;
	    RECT 0.6000 134.8000 1.0000 135.2000 ;
	    RECT 0.6000 126.1000 0.9000 134.8000 ;
	    RECT 1.4000 126.1000 1.8000 126.2000 ;
	    RECT 0.6000 125.8000 1.8000 126.1000 ;
	    RECT 0.6000 97.8000 1.0000 98.2000 ;
	    RECT 0.6000 95.2000 0.9000 97.8000 ;
	    RECT 0.6000 94.8000 1.0000 95.2000 ;
	    RECT 5.4000 75.1000 5.8000 75.2000 ;
	    RECT 6.2000 75.1000 6.6000 75.2000 ;
	    RECT 5.4000 74.8000 6.6000 75.1000 ;
	    RECT 7.8000 75.1000 8.2000 75.2000 ;
	    RECT 8.6000 75.1000 9.0000 75.2000 ;
	    RECT 7.8000 74.8000 9.0000 75.1000 ;
         LAYER metal3 ;
	    RECT 0.6000 145.1000 1.0000 145.2000 ;
	    RECT 11.8000 145.1000 12.2000 145.2000 ;
	    RECT 0.6000 144.8000 12.2000 145.1000 ;
	    RECT 0.6000 126.1000 1.0000 126.2000 ;
	    RECT 1.4000 126.1000 1.8000 126.2000 ;
	    RECT 0.6000 125.8000 1.8000 126.1000 ;
	    RECT 0.6000 98.8000 1.0000 99.2000 ;
	    RECT 0.6000 98.2000 0.9000 98.8000 ;
	    RECT 0.6000 97.8000 1.0000 98.2000 ;
	    RECT -2.6000 95.1000 -2.2000 95.2000 ;
	    RECT 0.6000 95.1000 1.0000 95.2000 ;
	    RECT 4.6000 95.1000 5.0000 95.2000 ;
	    RECT -2.6000 94.8000 5.0000 95.1000 ;
	    RECT 4.6000 75.1000 5.0000 75.2000 ;
	    RECT 5.4000 75.1000 5.8000 75.2000 ;
	    RECT 7.8000 75.1000 8.2000 75.2000 ;
	    RECT 4.6000 74.8000 8.2000 75.1000 ;
         LAYER metal4 ;
	    RECT 0.6000 125.8000 1.0000 126.2000 ;
	    RECT 0.6000 99.2000 0.9000 125.8000 ;
	    RECT 0.6000 98.8000 1.0000 99.2000 ;
	    RECT 4.6000 94.8000 5.0000 95.2000 ;
	    RECT 4.6000 75.2000 4.9000 94.8000 ;
	    RECT 4.6000 74.8000 5.0000 75.2000 ;
      END
   END SEL_A[5]
   PIN SEL_A[4]
      PORT
         LAYER metal1 ;
	    RECT 3.0000 133.4000 3.4000 134.2000 ;
	    RECT 15.8000 133.4000 16.2000 134.2000 ;
	    RECT 21.4000 133.4000 21.8000 134.2000 ;
	    RECT 2.2000 126.8000 2.6000 127.6000 ;
	    RECT 11.0000 85.1000 11.4000 85.2000 ;
	    RECT 11.8000 85.1000 12.2000 85.6000 ;
	    RECT 11.0000 84.8000 12.2000 85.1000 ;
	    RECT 18.2000 64.8000 18.6000 65.6000 ;
	    RECT 26.2000 55.4000 26.6000 56.2000 ;
	    RECT 11.0000 46.8000 11.4000 47.6000 ;
	    RECT 0.6000 44.8000 1.0000 45.6000 ;
         LAYER metal2 ;
	    RECT 3.0000 134.1000 3.4000 134.2000 ;
	    RECT 2.2000 133.8000 3.4000 134.1000 ;
	    RECT 15.8000 133.8000 16.2000 134.2000 ;
	    RECT 21.4000 133.8000 21.8000 134.2000 ;
	    RECT 2.2000 132.2000 2.5000 133.8000 ;
	    RECT 15.8000 132.2000 16.1000 133.8000 ;
	    RECT 21.4000 132.2000 21.7000 133.8000 ;
	    RECT 2.2000 131.8000 2.6000 132.2000 ;
	    RECT 15.8000 131.8000 16.2000 132.2000 ;
	    RECT 21.4000 131.8000 21.8000 132.2000 ;
	    RECT 2.2000 127.2000 2.5000 131.8000 ;
	    RECT 2.2000 126.8000 2.6000 127.2000 ;
	    RECT 2.2000 120.2000 2.5000 126.8000 ;
	    RECT 2.2000 119.8000 2.6000 120.2000 ;
	    RECT 11.0000 84.8000 11.4000 85.2000 ;
	    RECT 11.0000 84.2000 11.3000 84.8000 ;
	    RECT 11.0000 83.8000 11.4000 84.2000 ;
	    RECT 18.2000 64.8000 18.6000 65.2000 ;
	    RECT 18.2000 56.2000 18.5000 64.8000 ;
	    RECT 18.2000 55.8000 18.6000 56.2000 ;
	    RECT 25.4000 56.1000 25.8000 56.2000 ;
	    RECT 26.2000 56.1000 26.6000 56.2000 ;
	    RECT 25.4000 55.8000 26.6000 56.1000 ;
	    RECT 11.0000 47.8000 11.4000 48.2000 ;
	    RECT 11.0000 47.2000 11.3000 47.8000 ;
	    RECT 11.0000 46.8000 11.4000 47.2000 ;
	    RECT 0.6000 45.8000 1.0000 46.2000 ;
	    RECT 0.6000 45.2000 0.9000 45.8000 ;
	    RECT 0.6000 44.8000 1.0000 45.2000 ;
         LAYER metal3 ;
	    RECT 2.2000 132.1000 2.6000 132.2000 ;
	    RECT 15.8000 132.1000 16.2000 132.2000 ;
	    RECT 21.4000 132.1000 21.8000 132.2000 ;
	    RECT 2.2000 131.8000 21.8000 132.1000 ;
	    RECT 2.2000 120.1000 2.6000 120.2000 ;
	    RECT 11.0000 120.1000 11.4000 120.2000 ;
	    RECT 2.2000 119.8000 11.4000 120.1000 ;
	    RECT 11.0000 84.8000 11.4000 85.2000 ;
	    RECT 11.0000 84.2000 11.3000 84.8000 ;
	    RECT 11.0000 83.8000 11.4000 84.2000 ;
	    RECT 11.0000 56.1000 11.4000 56.2000 ;
	    RECT 18.2000 56.1000 18.6000 56.2000 ;
	    RECT 25.4000 56.1000 25.8000 56.2000 ;
	    RECT 11.0000 55.8000 25.8000 56.1000 ;
	    RECT 11.0000 47.8000 11.4000 48.2000 ;
	    RECT 11.0000 47.2000 11.3000 47.8000 ;
	    RECT 11.0000 46.8000 11.4000 47.2000 ;
	    RECT 0.6000 45.8000 1.0000 46.2000 ;
	    RECT -2.6000 45.1000 -2.2000 45.2000 ;
	    RECT 0.6000 45.1000 0.9000 45.8000 ;
	    RECT 11.0000 45.1000 11.4000 45.2000 ;
	    RECT -2.6000 44.8000 11.4000 45.1000 ;
         LAYER metal4 ;
	    RECT 11.0000 119.8000 11.4000 120.2000 ;
	    RECT 11.0000 85.2000 11.3000 119.8000 ;
	    RECT 11.0000 84.8000 11.4000 85.2000 ;
	    RECT 11.0000 56.2000 11.3000 84.8000 ;
	    RECT 11.0000 55.8000 11.4000 56.2000 ;
	    RECT 11.0000 47.2000 11.3000 55.8000 ;
	    RECT 11.0000 46.8000 11.4000 47.2000 ;
	    RECT 11.0000 45.2000 11.3000 46.8000 ;
	    RECT 11.0000 44.8000 11.4000 45.2000 ;
      END
   END SEL_A[4]
   PIN SEL_A[3]
      PORT
         LAYER metal1 ;
	    RECT 5.4000 124.8000 5.8000 125.6000 ;
	    RECT 8.6000 124.8000 9.0000 125.6000 ;
	    RECT 11.8000 124.8000 12.2000 125.6000 ;
	    RECT 3.8000 66.8000 4.2000 67.6000 ;
	    RECT 11.8000 64.8000 12.2000 66.2000 ;
         LAYER metal2 ;
	    RECT 5.4000 124.8000 5.8000 125.2000 ;
	    RECT 8.6000 124.8000 9.0000 125.2000 ;
	    RECT 11.0000 125.1000 11.4000 125.2000 ;
	    RECT 11.8000 125.1000 12.2000 125.2000 ;
	    RECT 11.0000 124.8000 12.2000 125.1000 ;
	    RECT 5.4000 119.2000 5.7000 124.8000 ;
	    RECT 8.6000 124.2000 8.9000 124.8000 ;
	    RECT 8.6000 123.8000 9.0000 124.2000 ;
	    RECT 5.4000 118.8000 5.8000 119.2000 ;
	    RECT 3.8000 79.8000 4.2000 80.2000 ;
	    RECT 3.8000 67.2000 4.1000 79.8000 ;
	    RECT 3.8000 66.8000 4.2000 67.2000 ;
	    RECT 3.8000 66.2000 4.1000 66.8000 ;
	    RECT 3.8000 65.8000 4.2000 66.2000 ;
	    RECT 11.8000 66.1000 12.2000 66.2000 ;
	    RECT 12.6000 66.1000 13.0000 66.2000 ;
	    RECT 11.8000 65.8000 13.0000 66.1000 ;
         LAYER metal3 ;
	    RECT 5.4000 125.1000 5.8000 125.2000 ;
	    RECT 11.0000 125.1000 11.4000 125.2000 ;
	    RECT 5.4000 124.8000 11.4000 125.1000 ;
	    RECT 8.6000 124.2000 8.9000 124.8000 ;
	    RECT 8.6000 123.8000 9.0000 124.2000 ;
	    RECT 5.4000 118.8000 5.8000 119.2000 ;
	    RECT 5.4000 118.2000 5.7000 118.8000 ;
	    RECT 5.4000 117.8000 5.8000 118.2000 ;
	    RECT -2.6000 80.1000 -2.2000 80.2000 ;
	    RECT 3.8000 80.1000 4.2000 80.2000 ;
	    RECT 5.4000 80.1000 5.8000 80.2000 ;
	    RECT -2.6000 79.8000 5.8000 80.1000 ;
	    RECT 3.8000 66.1000 4.2000 66.2000 ;
	    RECT 12.6000 66.1000 13.0000 66.2000 ;
	    RECT 3.8000 65.8000 13.0000 66.1000 ;
         LAYER metal4 ;
	    RECT 5.4000 117.8000 5.8000 118.2000 ;
	    RECT 5.4000 80.2000 5.7000 117.8000 ;
	    RECT 5.4000 79.8000 5.8000 80.2000 ;
      END
   END SEL_A[3]
   PIN SEL_A[2]
      PORT
         LAYER metal1 ;
	    RECT 42.2000 154.4000 42.6000 155.2000 ;
	    RECT 54.2000 154.4000 54.6000 155.2000 ;
	    RECT 39.8000 114.4000 40.2000 115.2000 ;
	    RECT 60.6000 115.1000 61.0000 115.2000 ;
	    RECT 63.0000 115.1000 63.4000 115.2000 ;
	    RECT 60.6000 114.8000 63.4000 115.1000 ;
	    RECT 60.6000 114.4000 61.0000 114.8000 ;
	    RECT 63.0000 114.4000 63.4000 114.8000 ;
         LAYER metal2 ;
	    RECT 55.0000 164.1000 55.4000 164.2000 ;
	    RECT 54.2000 163.8000 55.4000 164.1000 ;
	    RECT 54.2000 156.2000 54.5000 163.8000 ;
	    RECT 42.2000 155.8000 42.6000 156.2000 ;
	    RECT 54.2000 155.8000 54.6000 156.2000 ;
	    RECT 42.2000 155.2000 42.5000 155.8000 ;
	    RECT 54.2000 155.2000 54.5000 155.8000 ;
	    RECT 42.2000 154.8000 42.6000 155.2000 ;
	    RECT 54.2000 154.8000 54.6000 155.2000 ;
	    RECT 54.2000 135.2000 54.5000 154.8000 ;
	    RECT 54.2000 134.8000 54.6000 135.2000 ;
	    RECT 39.8000 115.1000 40.2000 115.2000 ;
	    RECT 40.6000 115.1000 41.0000 115.2000 ;
	    RECT 39.8000 114.8000 41.0000 115.1000 ;
	    RECT 60.6000 115.1000 61.0000 115.2000 ;
	    RECT 61.4000 115.1000 61.8000 115.2000 ;
	    RECT 60.6000 114.8000 61.8000 115.1000 ;
         LAYER metal3 ;
	    RECT 42.2000 156.1000 42.6000 156.2000 ;
	    RECT 54.2000 156.1000 54.6000 156.2000 ;
	    RECT 42.2000 155.8000 54.6000 156.1000 ;
	    RECT 54.2000 135.1000 54.6000 135.2000 ;
	    RECT 55.0000 135.1000 55.4000 135.2000 ;
	    RECT 54.2000 134.8000 55.4000 135.1000 ;
	    RECT 40.6000 115.1000 41.0000 115.2000 ;
	    RECT 54.2000 115.1000 54.6000 115.2000 ;
	    RECT 61.4000 115.1000 61.8000 115.2000 ;
	    RECT 40.6000 114.8000 61.8000 115.1000 ;
         LAYER metal4 ;
	    RECT 55.0000 135.1000 55.4000 135.2000 ;
	    RECT 54.2000 134.8000 55.4000 135.1000 ;
	    RECT 54.2000 115.2000 54.5000 134.8000 ;
	    RECT 54.2000 114.8000 54.6000 115.2000 ;
      END
   END SEL_A[2]
   PIN SEL_A[1]
      PORT
         LAYER metal1 ;
	    RECT 51.0000 153.4000 51.4000 154.2000 ;
	    RECT 71.0000 153.4000 71.4000 154.2000 ;
	    RECT 80.6000 133.4000 81.0000 134.2000 ;
	    RECT 80.6000 126.8000 81.0000 127.6000 ;
	    RECT 55.8000 115.4000 56.2000 116.2000 ;
	    RECT 51.0000 104.8000 51.4000 105.6000 ;
	    RECT 87.0000 95.4000 87.4000 96.2000 ;
	    RECT 90.2000 95.4000 90.6000 96.2000 ;
	    RECT 70.2000 86.8000 70.6000 87.6000 ;
         LAYER metal2 ;
	    RECT 75.0000 163.8000 75.4000 164.2000 ;
	    RECT 75.0000 154.2000 75.3000 163.8000 ;
	    RECT 51.0000 153.8000 51.4000 154.2000 ;
	    RECT 70.2000 154.1000 70.6000 154.2000 ;
	    RECT 71.0000 154.1000 71.4000 154.2000 ;
	    RECT 70.2000 153.8000 71.4000 154.1000 ;
	    RECT 75.0000 153.8000 75.4000 154.2000 ;
	    RECT 80.6000 153.8000 81.0000 154.2000 ;
	    RECT 51.0000 153.2000 51.3000 153.8000 ;
	    RECT 51.0000 152.8000 51.4000 153.2000 ;
	    RECT 80.6000 134.2000 80.9000 153.8000 ;
	    RECT 80.6000 133.8000 81.0000 134.2000 ;
	    RECT 80.6000 127.2000 80.9000 133.8000 ;
	    RECT 80.6000 126.8000 81.0000 127.2000 ;
	    RECT 80.6000 119.2000 80.9000 126.8000 ;
	    RECT 55.8000 118.8000 56.2000 119.2000 ;
	    RECT 80.6000 118.8000 81.0000 119.2000 ;
	    RECT 55.8000 116.2000 56.1000 118.8000 ;
	    RECT 80.6000 117.2000 80.9000 118.8000 ;
	    RECT 80.6000 116.8000 81.0000 117.2000 ;
	    RECT 90.2000 116.8000 90.6000 117.2000 ;
	    RECT 55.8000 115.8000 56.2000 116.2000 ;
	    RECT 55.8000 109.2000 56.1000 115.8000 ;
	    RECT 51.0000 108.8000 51.4000 109.2000 ;
	    RECT 55.8000 108.8000 56.2000 109.2000 ;
	    RECT 51.0000 105.2000 51.3000 108.8000 ;
	    RECT 51.0000 104.8000 51.4000 105.2000 ;
	    RECT 90.2000 96.2000 90.5000 116.8000 ;
	    RECT 87.0000 96.1000 87.4000 96.2000 ;
	    RECT 87.8000 96.1000 88.2000 96.2000 ;
	    RECT 87.0000 95.8000 88.2000 96.1000 ;
	    RECT 90.2000 95.8000 90.6000 96.2000 ;
	    RECT 70.2000 92.8000 70.6000 93.2000 ;
	    RECT 70.2000 87.2000 70.5000 92.8000 ;
	    RECT 70.2000 86.8000 70.6000 87.2000 ;
         LAYER metal3 ;
	    RECT 70.2000 154.1000 70.6000 154.2000 ;
	    RECT 75.0000 154.1000 75.4000 154.2000 ;
	    RECT 80.6000 154.1000 81.0000 154.2000 ;
	    RECT 51.0000 153.8000 81.0000 154.1000 ;
	    RECT 51.0000 153.2000 51.3000 153.8000 ;
	    RECT 51.0000 152.8000 51.4000 153.2000 ;
	    RECT 55.8000 119.1000 56.2000 119.2000 ;
	    RECT 71.0000 119.1000 71.4000 119.2000 ;
	    RECT 80.6000 119.1000 81.0000 119.2000 ;
	    RECT 55.8000 118.8000 81.0000 119.1000 ;
	    RECT 80.6000 117.1000 81.0000 117.2000 ;
	    RECT 90.2000 117.1000 90.6000 117.2000 ;
	    RECT 80.6000 116.8000 90.6000 117.1000 ;
	    RECT 51.0000 109.1000 51.4000 109.2000 ;
	    RECT 55.8000 109.1000 56.2000 109.2000 ;
	    RECT 51.0000 108.8000 56.2000 109.1000 ;
	    RECT 87.8000 96.1000 88.2000 96.2000 ;
	    RECT 90.2000 96.1000 90.6000 96.2000 ;
	    RECT 87.8000 95.8000 90.6000 96.1000 ;
	    RECT 70.2000 93.1000 70.6000 93.2000 ;
	    RECT 71.0000 93.1000 71.4000 93.2000 ;
	    RECT 70.2000 92.8000 71.4000 93.1000 ;
         LAYER metal4 ;
	    RECT 71.0000 118.8000 71.4000 119.2000 ;
	    RECT 71.0000 93.2000 71.3000 118.8000 ;
	    RECT 71.0000 92.8000 71.4000 93.2000 ;
      END
   END SEL_A[1]
   PIN SEL_A[0]
      PORT
         LAYER metal1 ;
	    RECT 59.0000 144.8000 59.4000 145.6000 ;
	    RECT 67.8000 144.8000 68.2000 145.6000 ;
	    RECT 76.6000 125.1000 77.0000 125.2000 ;
	    RECT 77.4000 125.1000 77.8000 125.6000 ;
	    RECT 76.6000 124.8000 77.8000 125.1000 ;
	    RECT 76.6000 106.8000 77.0000 107.6000 ;
	    RECT 71.0000 104.8000 71.4000 105.6000 ;
         LAYER metal2 ;
	    RECT 71.0000 163.8000 71.4000 164.2000 ;
	    RECT 71.0000 159.2000 71.3000 163.8000 ;
	    RECT 67.8000 158.8000 68.2000 159.2000 ;
	    RECT 71.0000 158.8000 71.4000 159.2000 ;
	    RECT 67.8000 146.2000 68.1000 158.8000 ;
	    RECT 59.0000 145.8000 59.4000 146.2000 ;
	    RECT 67.8000 145.8000 68.2000 146.2000 ;
	    RECT 59.0000 145.2000 59.3000 145.8000 ;
	    RECT 67.8000 145.2000 68.1000 145.8000 ;
	    RECT 59.0000 144.8000 59.4000 145.2000 ;
	    RECT 67.8000 145.1000 68.2000 145.2000 ;
	    RECT 68.6000 145.1000 69.0000 145.2000 ;
	    RECT 67.8000 144.8000 69.0000 145.1000 ;
	    RECT 75.8000 144.8000 76.2000 145.2000 ;
	    RECT 75.8000 127.1000 76.1000 144.8000 ;
	    RECT 75.8000 126.8000 76.9000 127.1000 ;
	    RECT 76.6000 125.2000 76.9000 126.8000 ;
	    RECT 76.6000 124.8000 77.0000 125.2000 ;
	    RECT 76.6000 107.2000 76.9000 124.8000 ;
	    RECT 71.0000 106.8000 71.4000 107.2000 ;
	    RECT 76.6000 106.8000 77.0000 107.2000 ;
	    RECT 71.0000 105.2000 71.3000 106.8000 ;
	    RECT 71.0000 104.8000 71.4000 105.2000 ;
         LAYER metal3 ;
	    RECT 67.8000 159.1000 68.2000 159.2000 ;
	    RECT 71.0000 159.1000 71.4000 159.2000 ;
	    RECT 67.8000 158.8000 71.4000 159.1000 ;
	    RECT 59.0000 146.1000 59.4000 146.2000 ;
	    RECT 67.8000 146.1000 68.2000 146.2000 ;
	    RECT 59.0000 145.8000 68.2000 146.1000 ;
	    RECT 68.6000 145.1000 69.0000 145.2000 ;
	    RECT 75.8000 145.1000 76.2000 145.2000 ;
	    RECT 68.6000 144.8000 76.2000 145.1000 ;
	    RECT 71.0000 107.1000 71.4000 107.2000 ;
	    RECT 76.6000 107.1000 77.0000 107.2000 ;
	    RECT 71.0000 106.8000 77.0000 107.1000 ;
      END
   END SEL_A[0]
   PIN SEL_AB[3]
      PORT
         LAYER metal1 ;
	    RECT 40.6000 73.4000 41.0000 74.2000 ;
	    RECT 59.0000 55.4000 59.4000 56.2000 ;
	    RECT 73.4000 55.4000 73.8000 56.2000 ;
	    RECT 76.6000 56.1000 77.0000 56.2000 ;
	    RECT 77.4000 56.1000 77.8000 56.2000 ;
	    RECT 76.6000 55.8000 77.8000 56.1000 ;
	    RECT 76.6000 55.4000 77.0000 55.8000 ;
	    RECT 77.4000 55.4000 77.8000 55.8000 ;
         LAYER metal2 ;
	    RECT 40.6000 73.8000 41.0000 74.2000 ;
	    RECT 40.6000 64.2000 40.9000 73.8000 ;
	    RECT 40.6000 63.8000 41.0000 64.2000 ;
	    RECT 40.6000 60.2000 40.9000 63.8000 ;
	    RECT 59.0000 61.8000 59.4000 62.2000 ;
	    RECT 73.4000 61.8000 73.8000 62.2000 ;
	    RECT 59.0000 60.2000 59.3000 61.8000 ;
	    RECT 40.6000 59.8000 41.0000 60.2000 ;
	    RECT 59.0000 59.8000 59.4000 60.2000 ;
	    RECT 59.0000 56.2000 59.3000 59.8000 ;
	    RECT 73.4000 56.2000 73.7000 61.8000 ;
	    RECT 59.0000 55.8000 59.4000 56.2000 ;
	    RECT 73.4000 55.8000 73.8000 56.2000 ;
	    RECT 75.8000 56.1000 76.2000 56.2000 ;
	    RECT 76.6000 56.1000 77.0000 56.2000 ;
	    RECT 75.8000 55.8000 77.0000 56.1000 ;
         LAYER metal3 ;
	    RECT -2.6000 68.1000 -2.2000 68.2000 ;
	    RECT 0.6000 68.1000 1.0000 68.2000 ;
	    RECT -2.6000 67.8000 1.0000 68.1000 ;
	    RECT 0.6000 64.1000 1.0000 64.2000 ;
	    RECT 40.6000 64.1000 41.0000 64.2000 ;
	    RECT 0.6000 63.8000 41.0000 64.1000 ;
	    RECT 59.0000 62.1000 59.4000 62.2000 ;
	    RECT 73.4000 62.1000 73.8000 62.2000 ;
	    RECT 59.0000 61.8000 73.8000 62.1000 ;
	    RECT 40.6000 60.1000 41.0000 60.2000 ;
	    RECT 59.0000 60.1000 59.4000 60.2000 ;
	    RECT 40.6000 59.8000 59.4000 60.1000 ;
	    RECT 73.4000 56.1000 73.8000 56.2000 ;
	    RECT 75.8000 56.1000 76.2000 56.2000 ;
	    RECT 73.4000 55.8000 76.2000 56.1000 ;
         LAYER metal4 ;
	    RECT 0.6000 67.8000 1.0000 68.2000 ;
	    RECT 0.6000 64.2000 0.9000 67.8000 ;
	    RECT 0.6000 63.8000 1.0000 64.2000 ;
      END
   END SEL_AB[3]
   PIN SEL_AB[2]
      PORT
         LAYER metal1 ;
	    RECT 135.0000 55.4000 135.4000 56.2000 ;
	    RECT 134.2000 53.4000 134.6000 54.2000 ;
	    RECT 147.0000 44.8000 147.4000 45.6000 ;
	    RECT 151.0000 35.4000 151.4000 36.2000 ;
	    RECT 161.4000 35.4000 161.8000 36.2000 ;
         LAYER metal2 ;
	    RECT 135.0000 56.1000 135.4000 56.2000 ;
	    RECT 134.2000 55.8000 135.4000 56.1000 ;
	    RECT 134.2000 54.2000 134.5000 55.8000 ;
	    RECT 134.2000 53.8000 134.6000 54.2000 ;
	    RECT 134.2000 44.2000 134.5000 53.8000 ;
	    RECT 147.0000 44.8000 147.4000 45.2000 ;
	    RECT 147.0000 44.2000 147.3000 44.8000 ;
	    RECT 134.2000 43.8000 134.6000 44.2000 ;
	    RECT 147.0000 43.8000 147.4000 44.2000 ;
	    RECT 151.0000 43.8000 151.4000 44.2000 ;
	    RECT 151.0000 40.2000 151.3000 43.8000 ;
	    RECT 161.4000 41.8000 161.8000 42.2000 ;
	    RECT 161.4000 40.2000 161.7000 41.8000 ;
	    RECT 151.0000 39.8000 151.4000 40.2000 ;
	    RECT 161.4000 39.8000 161.8000 40.2000 ;
	    RECT 151.0000 36.2000 151.3000 39.8000 ;
	    RECT 161.4000 36.2000 161.7000 39.8000 ;
	    RECT 151.0000 35.8000 151.4000 36.2000 ;
	    RECT 161.4000 35.8000 161.8000 36.2000 ;
         LAYER metal3 ;
	    RECT 134.2000 44.1000 134.6000 44.2000 ;
	    RECT 147.0000 44.1000 147.4000 44.2000 ;
	    RECT 151.0000 44.1000 151.4000 44.2000 ;
	    RECT 134.2000 43.8000 151.4000 44.1000 ;
	    RECT 161.4000 42.1000 161.8000 42.2000 ;
	    RECT 172.6000 42.1000 173.0000 42.2000 ;
	    RECT 161.4000 41.8000 173.0000 42.1000 ;
	    RECT 151.0000 40.1000 151.4000 40.2000 ;
	    RECT 161.4000 40.1000 161.8000 40.2000 ;
	    RECT 151.0000 39.8000 161.8000 40.1000 ;
	    RECT 172.6000 36.1000 173.0000 36.2000 ;
	    RECT 175.8000 36.1000 176.2000 36.2000 ;
	    RECT 172.6000 35.8000 176.2000 36.1000 ;
         LAYER metal4 ;
	    RECT 172.6000 41.8000 173.0000 42.2000 ;
	    RECT 172.6000 36.2000 172.9000 41.8000 ;
	    RECT 172.6000 35.8000 173.0000 36.2000 ;
      END
   END SEL_AB[2]
   PIN SEL_AB[1]
      PORT
         LAYER metal1 ;
	    RECT 7.0000 53.4000 7.4000 54.2000 ;
	    RECT 23.8000 44.8000 24.2000 45.6000 ;
	    RECT 7.0000 35.4000 7.4000 36.2000 ;
	    RECT 12.6000 35.4000 13.0000 36.2000 ;
	    RECT 15.8000 35.4000 16.2000 36.2000 ;
         LAYER metal2 ;
	    RECT 7.0000 53.8000 7.4000 54.2000 ;
	    RECT 7.0000 50.2000 7.3000 53.8000 ;
	    RECT 7.0000 49.8000 7.4000 50.2000 ;
	    RECT 23.8000 44.8000 24.2000 45.2000 ;
	    RECT 23.8000 39.2000 24.1000 44.8000 ;
	    RECT 7.0000 38.8000 7.4000 39.2000 ;
	    RECT 12.6000 38.8000 13.0000 39.2000 ;
	    RECT 15.8000 38.8000 16.2000 39.2000 ;
	    RECT 23.8000 38.8000 24.2000 39.2000 ;
	    RECT 7.0000 36.2000 7.3000 38.8000 ;
	    RECT 12.6000 36.2000 12.9000 38.8000 ;
	    RECT 15.8000 36.2000 16.1000 38.8000 ;
	    RECT 7.0000 35.8000 7.4000 36.2000 ;
	    RECT 12.6000 35.8000 13.0000 36.2000 ;
	    RECT 15.8000 35.8000 16.2000 36.2000 ;
         LAYER metal3 ;
	    RECT 0.6000 50.1000 1.0000 50.2000 ;
	    RECT 7.0000 50.1000 7.4000 50.2000 ;
	    RECT 0.6000 49.8000 7.4000 50.1000 ;
	    RECT -2.6000 47.1000 -2.2000 47.2000 ;
	    RECT 0.6000 47.1000 1.0000 47.2000 ;
	    RECT -2.6000 46.8000 1.0000 47.1000 ;
	    RECT 0.6000 39.1000 1.0000 39.2000 ;
	    RECT 7.0000 39.1000 7.4000 39.2000 ;
	    RECT 12.6000 39.1000 13.0000 39.2000 ;
	    RECT 15.8000 39.1000 16.2000 39.2000 ;
	    RECT 23.8000 39.1000 24.2000 39.2000 ;
	    RECT 0.6000 38.8000 24.2000 39.1000 ;
         LAYER metal4 ;
	    RECT 0.6000 49.8000 1.0000 50.2000 ;
	    RECT 0.6000 47.2000 0.9000 49.8000 ;
	    RECT 0.6000 46.8000 1.0000 47.2000 ;
	    RECT 0.6000 39.2000 0.9000 46.8000 ;
	    RECT 0.6000 38.8000 1.0000 39.2000 ;
      END
   END SEL_AB[1]
   PIN SEL_AB[0]
      PORT
         LAYER metal1 ;
	    RECT 110.2000 56.1000 110.6000 56.2000 ;
	    RECT 111.0000 56.1000 111.4000 56.2000 ;
	    RECT 110.2000 55.8000 111.4000 56.1000 ;
	    RECT 111.0000 55.4000 111.4000 55.8000 ;
	    RECT 115.8000 55.4000 116.2000 56.2000 ;
	    RECT 100.6000 53.4000 101.0000 54.2000 ;
	    RECT 99.0000 44.8000 99.4000 45.6000 ;
	    RECT 107.8000 35.4000 108.2000 36.2000 ;
         LAYER metal2 ;
	    RECT 110.2000 55.8000 110.6000 56.2000 ;
	    RECT 115.0000 56.1000 115.4000 56.2000 ;
	    RECT 115.8000 56.1000 116.2000 56.2000 ;
	    RECT 115.0000 55.8000 116.2000 56.1000 ;
	    RECT 100.6000 53.8000 101.0000 54.2000 ;
	    RECT 100.6000 50.2000 100.9000 53.8000 ;
	    RECT 110.2000 50.2000 110.5000 55.8000 ;
	    RECT 99.0000 49.8000 99.4000 50.2000 ;
	    RECT 100.6000 49.8000 101.0000 50.2000 ;
	    RECT 107.8000 49.8000 108.2000 50.2000 ;
	    RECT 110.2000 49.8000 110.6000 50.2000 ;
	    RECT 99.0000 45.2000 99.3000 49.8000 ;
	    RECT 99.0000 44.8000 99.4000 45.2000 ;
	    RECT 107.8000 36.2000 108.1000 49.8000 ;
	    RECT 107.8000 36.1000 108.2000 36.2000 ;
	    RECT 108.6000 36.1000 109.0000 36.2000 ;
	    RECT 107.8000 35.8000 109.0000 36.1000 ;
	    RECT 116.6000 0.8000 117.0000 1.2000 ;
	    RECT 116.6000 -1.8000 116.9000 0.8000 ;
	    RECT 116.6000 -2.2000 117.0000 -1.8000 ;
         LAYER metal3 ;
	    RECT 110.2000 56.1000 110.6000 56.2000 ;
	    RECT 115.0000 56.1000 115.4000 56.2000 ;
	    RECT 110.2000 55.8000 115.4000 56.1000 ;
	    RECT 99.0000 50.1000 99.4000 50.2000 ;
	    RECT 100.6000 50.1000 101.0000 50.2000 ;
	    RECT 107.8000 50.1000 108.2000 50.2000 ;
	    RECT 110.2000 50.1000 110.6000 50.2000 ;
	    RECT 99.0000 49.8000 110.6000 50.1000 ;
	    RECT 107.8000 36.1000 108.2000 36.2000 ;
	    RECT 108.6000 36.1000 109.0000 36.2000 ;
	    RECT 107.8000 35.8000 109.0000 36.1000 ;
	    RECT 107.8000 1.1000 108.2000 1.2000 ;
	    RECT 116.6000 1.1000 117.0000 1.2000 ;
	    RECT 107.8000 0.8000 117.0000 1.1000 ;
         LAYER metal4 ;
	    RECT 107.8000 35.8000 108.2000 36.2000 ;
	    RECT 107.8000 1.2000 108.1000 35.8000 ;
	    RECT 107.8000 0.8000 108.2000 1.2000 ;
      END
   END SEL_AB[0]
   PIN SEL_B[11]
      PORT
         LAYER metal1 ;
	    RECT 60.6000 26.1000 61.0000 26.6000 ;
	    RECT 62.2000 26.1000 62.6000 26.2000 ;
	    RECT 60.6000 25.8000 62.6000 26.1000 ;
	    RECT 69.4000 25.8000 69.8000 26.6000 ;
	    RECT 80.6000 25.8000 81.0000 26.6000 ;
	    RECT 59.0000 5.8000 59.4000 6.6000 ;
	    RECT 79.0000 5.8000 79.4000 6.6000 ;
         LAYER metal2 ;
	    RECT 62.2000 26.1000 62.6000 26.2000 ;
	    RECT 63.0000 26.1000 63.4000 26.2000 ;
	    RECT 62.2000 25.8000 63.4000 26.1000 ;
	    RECT 68.6000 26.1000 69.0000 26.2000 ;
	    RECT 69.4000 26.1000 69.8000 26.2000 ;
	    RECT 68.6000 25.8000 69.8000 26.1000 ;
	    RECT 79.8000 26.1000 80.2000 26.2000 ;
	    RECT 80.6000 26.1000 81.0000 26.2000 ;
	    RECT 79.8000 25.8000 81.0000 26.1000 ;
	    RECT 62.2000 22.2000 62.5000 25.8000 ;
	    RECT 59.0000 21.8000 59.4000 22.2000 ;
	    RECT 62.2000 21.8000 62.6000 22.2000 ;
	    RECT 59.0000 6.2000 59.3000 21.8000 ;
	    RECT 59.0000 5.8000 59.4000 6.2000 ;
	    RECT 79.0000 6.1000 79.4000 6.2000 ;
	    RECT 79.8000 6.1000 80.1000 25.8000 ;
	    RECT 79.0000 5.8000 80.1000 6.1000 ;
	    RECT 79.8000 1.2000 80.1000 5.8000 ;
	    RECT 79.8000 0.8000 80.2000 1.2000 ;
	    RECT 81.4000 0.8000 81.8000 1.2000 ;
	    RECT 81.4000 -1.8000 81.7000 0.8000 ;
	    RECT 81.4000 -2.2000 81.8000 -1.8000 ;
         LAYER metal3 ;
	    RECT 63.0000 26.1000 63.4000 26.2000 ;
	    RECT 68.6000 26.1000 69.0000 26.2000 ;
	    RECT 79.8000 26.1000 80.2000 26.2000 ;
	    RECT 63.0000 25.8000 80.2000 26.1000 ;
	    RECT 59.0000 22.1000 59.4000 22.2000 ;
	    RECT 62.2000 22.1000 62.6000 22.2000 ;
	    RECT 59.0000 21.8000 62.6000 22.1000 ;
	    RECT 79.8000 1.1000 80.2000 1.2000 ;
	    RECT 81.4000 1.1000 81.8000 1.2000 ;
	    RECT 79.8000 0.8000 81.8000 1.1000 ;
      END
   END SEL_B[11]
   PIN SEL_B[10]
      PORT
         LAYER metal1 ;
	    RECT 71.0000 44.8000 71.4000 45.6000 ;
	    RECT 83.0000 45.1000 83.4000 45.2000 ;
	    RECT 83.8000 45.1000 84.2000 45.6000 ;
	    RECT 83.0000 44.8000 84.2000 45.1000 ;
	    RECT 59.0000 34.1000 59.4000 34.2000 ;
	    RECT 59.8000 34.1000 60.2000 34.2000 ;
	    RECT 59.0000 33.8000 60.2000 34.1000 ;
	    RECT 82.2000 34.1000 82.6000 34.2000 ;
	    RECT 83.0000 34.1000 83.4000 34.2000 ;
	    RECT 82.2000 33.8000 83.4000 34.1000 ;
	    RECT 59.0000 33.4000 59.4000 33.8000 ;
	    RECT 82.2000 33.4000 82.6000 33.8000 ;
	    RECT 64.6000 26.8000 65.0000 27.6000 ;
	    RECT 67.0000 26.8000 67.4000 27.6000 ;
	    RECT 78.2000 26.8000 78.6000 27.6000 ;
	    RECT 55.0000 24.8000 55.4000 25.6000 ;
	    RECT 84.6000 15.4000 85.0000 16.2000 ;
         LAYER metal2 ;
	    RECT 71.0000 45.1000 71.4000 45.2000 ;
	    RECT 71.8000 45.1000 72.2000 45.2000 ;
	    RECT 71.0000 44.8000 72.2000 45.1000 ;
	    RECT 83.0000 44.8000 83.4000 45.2000 ;
	    RECT 83.0000 34.2000 83.3000 44.8000 ;
	    RECT 59.8000 33.8000 60.2000 34.2000 ;
	    RECT 78.2000 33.8000 78.6000 34.2000 ;
	    RECT 83.0000 33.8000 83.4000 34.2000 ;
	    RECT 59.8000 27.2000 60.1000 33.8000 ;
	    RECT 78.2000 27.2000 78.5000 33.8000 ;
	    RECT 55.0000 26.8000 55.4000 27.2000 ;
	    RECT 59.8000 26.8000 60.2000 27.2000 ;
	    RECT 64.6000 27.1000 65.0000 27.2000 ;
	    RECT 65.4000 27.1000 65.8000 27.2000 ;
	    RECT 64.6000 26.8000 65.8000 27.1000 ;
	    RECT 67.0000 27.1000 67.4000 27.2000 ;
	    RECT 67.8000 27.1000 68.2000 27.2000 ;
	    RECT 67.0000 26.8000 68.2000 27.1000 ;
	    RECT 78.2000 26.8000 78.6000 27.2000 ;
	    RECT 84.6000 26.8000 85.0000 27.2000 ;
	    RECT 55.0000 25.2000 55.3000 26.8000 ;
	    RECT 55.0000 24.8000 55.4000 25.2000 ;
	    RECT 84.6000 16.2000 84.9000 26.8000 ;
	    RECT 84.6000 15.8000 85.0000 16.2000 ;
	    RECT 84.6000 12.1000 84.9000 15.8000 ;
	    RECT 85.4000 12.1000 85.8000 12.2000 ;
	    RECT 84.6000 11.8000 85.8000 12.1000 ;
	    RECT 83.8000 6.8000 84.2000 7.2000 ;
	    RECT 83.8000 -1.8000 84.1000 6.8000 ;
	    RECT 83.8000 -2.2000 84.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 71.8000 45.1000 72.2000 45.2000 ;
	    RECT 83.0000 45.1000 83.4000 45.2000 ;
	    RECT 71.8000 44.8000 83.4000 45.1000 ;
	    RECT 78.2000 34.1000 78.6000 34.2000 ;
	    RECT 83.0000 34.1000 83.4000 34.2000 ;
	    RECT 78.2000 33.8000 83.4000 34.1000 ;
	    RECT 55.0000 27.1000 55.4000 27.2000 ;
	    RECT 59.8000 27.1000 60.2000 27.2000 ;
	    RECT 65.4000 27.1000 65.8000 27.2000 ;
	    RECT 67.8000 27.1000 68.2000 27.2000 ;
	    RECT 78.2000 27.1000 78.6000 27.2000 ;
	    RECT 84.6000 27.1000 85.0000 27.2000 ;
	    RECT 55.0000 26.8000 85.0000 27.1000 ;
	    RECT 84.6000 12.1000 85.0000 12.2000 ;
	    RECT 85.4000 12.1000 85.8000 12.2000 ;
	    RECT 84.6000 11.8000 85.8000 12.1000 ;
	    RECT 83.8000 7.1000 84.2000 7.2000 ;
	    RECT 84.6000 7.1000 85.0000 7.2000 ;
	    RECT 83.8000 6.8000 85.0000 7.1000 ;
         LAYER metal4 ;
	    RECT 84.6000 11.8000 85.0000 12.2000 ;
	    RECT 84.6000 7.2000 84.9000 11.8000 ;
	    RECT 84.6000 6.8000 85.0000 7.2000 ;
      END
   END SEL_B[10]
   PIN SEL_B[9]
      PORT
         LAYER metal1 ;
	    RECT 69.4000 35.4000 69.8000 36.2000 ;
	    RECT 75.0000 35.4000 75.4000 36.2000 ;
	    RECT 61.4000 33.4000 61.8000 34.2000 ;
	    RECT 58.2000 24.8000 58.6000 25.6000 ;
	    RECT 81.4000 24.8000 81.8000 25.6000 ;
         LAYER metal2 ;
	    RECT 69.4000 35.8000 69.8000 36.2000 ;
	    RECT 75.0000 35.8000 75.4000 36.2000 ;
	    RECT 69.4000 35.2000 69.7000 35.8000 ;
	    RECT 75.0000 35.2000 75.3000 35.8000 ;
	    RECT 61.4000 34.8000 61.8000 35.2000 ;
	    RECT 69.4000 34.8000 69.8000 35.2000 ;
	    RECT 75.0000 34.8000 75.4000 35.2000 ;
	    RECT 61.4000 34.2000 61.7000 34.8000 ;
	    RECT 61.4000 33.8000 61.8000 34.2000 ;
	    RECT 61.4000 26.2000 61.7000 33.8000 ;
	    RECT 58.2000 25.8000 58.6000 26.2000 ;
	    RECT 61.4000 25.8000 61.8000 26.2000 ;
	    RECT 58.2000 25.2000 58.5000 25.8000 ;
	    RECT 58.2000 24.8000 58.6000 25.2000 ;
	    RECT 80.6000 25.1000 81.0000 25.2000 ;
	    RECT 81.4000 25.1000 81.8000 25.2000 ;
	    RECT 80.6000 24.8000 81.8000 25.1000 ;
	    RECT 79.0000 0.8000 79.4000 1.2000 ;
	    RECT 79.0000 -1.9000 79.3000 0.8000 ;
	    RECT 79.8000 -1.9000 80.2000 -1.8000 ;
	    RECT 79.0000 -2.2000 80.2000 -1.9000 ;
         LAYER metal3 ;
	    RECT 61.4000 35.1000 61.8000 35.2000 ;
	    RECT 69.4000 35.1000 69.8000 35.2000 ;
	    RECT 75.0000 35.1000 75.4000 35.2000 ;
	    RECT 61.4000 34.8000 75.4000 35.1000 ;
	    RECT 58.2000 26.1000 58.6000 26.2000 ;
	    RECT 61.4000 26.1000 61.8000 26.2000 ;
	    RECT 58.2000 25.8000 61.8000 26.1000 ;
	    RECT 75.0000 25.1000 75.4000 25.2000 ;
	    RECT 80.6000 25.1000 81.0000 25.2000 ;
	    RECT 75.0000 24.8000 81.0000 25.1000 ;
	    RECT 75.0000 1.1000 75.4000 1.2000 ;
	    RECT 79.0000 1.1000 79.4000 1.2000 ;
	    RECT 75.0000 0.8000 79.4000 1.1000 ;
         LAYER metal4 ;
	    RECT 75.0000 34.8000 75.4000 35.2000 ;
	    RECT 75.0000 25.2000 75.3000 34.8000 ;
	    RECT 75.0000 24.8000 75.4000 25.2000 ;
	    RECT 75.0000 1.2000 75.3000 24.8000 ;
	    RECT 75.0000 0.8000 75.4000 1.2000 ;
      END
   END SEL_B[9]
   PIN SEL_B[8]
      PORT
         LAYER metal1 ;
	    RECT 158.2000 34.4000 158.6000 35.2000 ;
	    RECT 160.6000 34.4000 161.0000 35.2000 ;
	    RECT 158.2000 25.8000 158.6000 26.6000 ;
	    RECT 171.0000 15.1000 171.4000 15.2000 ;
	    RECT 173.4000 15.1000 173.8000 15.2000 ;
	    RECT 171.0000 14.8000 173.8000 15.1000 ;
	    RECT 171.0000 14.4000 171.4000 14.8000 ;
	    RECT 168.6000 5.8000 169.0000 6.6000 ;
         LAYER metal2 ;
	    RECT 158.2000 35.1000 158.6000 35.2000 ;
	    RECT 159.0000 35.1000 159.4000 35.2000 ;
	    RECT 158.2000 34.8000 159.4000 35.1000 ;
	    RECT 160.6000 35.1000 161.0000 35.2000 ;
	    RECT 161.4000 35.1000 161.8000 35.2000 ;
	    RECT 160.6000 34.8000 161.8000 35.1000 ;
	    RECT 158.2000 26.2000 158.5000 34.8000 ;
	    RECT 158.2000 25.8000 158.6000 26.2000 ;
	    RECT 158.2000 19.2000 158.5000 25.8000 ;
	    RECT 158.2000 18.8000 158.6000 19.2000 ;
	    RECT 171.0000 18.8000 171.4000 19.2000 ;
	    RECT 171.0000 15.2000 171.3000 18.8000 ;
	    RECT 171.0000 14.8000 171.4000 15.2000 ;
	    RECT 173.4000 14.8000 173.8000 15.2000 ;
	    RECT 173.4000 6.2000 173.7000 14.8000 ;
	    RECT 168.6000 6.1000 169.0000 6.2000 ;
	    RECT 169.4000 6.1000 169.8000 6.2000 ;
	    RECT 168.6000 5.8000 169.8000 6.1000 ;
	    RECT 173.4000 5.8000 173.8000 6.2000 ;
         LAYER metal3 ;
	    RECT 159.0000 35.1000 159.4000 35.2000 ;
	    RECT 161.4000 35.1000 161.8000 35.2000 ;
	    RECT 159.0000 34.8000 161.8000 35.1000 ;
	    RECT 158.2000 19.1000 158.6000 19.2000 ;
	    RECT 171.0000 19.1000 171.4000 19.2000 ;
	    RECT 158.2000 18.8000 171.4000 19.1000 ;
	    RECT 169.4000 6.1000 169.8000 6.2000 ;
	    RECT 173.4000 6.1000 173.8000 6.2000 ;
	    RECT 175.8000 6.1000 176.2000 6.2000 ;
	    RECT 169.4000 5.8000 176.2000 6.1000 ;
      END
   END SEL_B[8]
   PIN SEL_B[7]
      PORT
         LAYER metal1 ;
	    RECT 144.6000 55.4000 145.0000 56.2000 ;
	    RECT 151.8000 53.4000 152.2000 54.2000 ;
	    RECT 167.8000 44.8000 168.2000 45.6000 ;
	    RECT 137.4000 26.8000 137.8000 27.6000 ;
	    RECT 147.8000 27.1000 148.2000 27.6000 ;
	    RECT 148.6000 27.1000 149.0000 27.6000 ;
	    RECT 147.8000 26.8000 149.0000 27.1000 ;
	    RECT 154.2000 26.8000 154.6000 27.6000 ;
	    RECT 148.6000 26.2000 148.9000 26.8000 ;
	    RECT 148.6000 25.8000 149.0000 26.2000 ;
	    RECT 124.6000 24.8000 125.0000 25.6000 ;
	    RECT 158.2000 15.4000 158.6000 16.2000 ;
         LAYER metal2 ;
	    RECT 144.6000 55.8000 145.0000 56.2000 ;
	    RECT 144.6000 54.2000 144.9000 55.8000 ;
	    RECT 144.6000 53.8000 145.0000 54.2000 ;
	    RECT 151.8000 53.8000 152.2000 54.2000 ;
	    RECT 151.8000 53.2000 152.1000 53.8000 ;
	    RECT 151.8000 52.8000 152.2000 53.2000 ;
	    RECT 167.8000 44.8000 168.2000 45.2000 ;
	    RECT 167.8000 44.2000 168.1000 44.8000 ;
	    RECT 167.8000 43.8000 168.2000 44.2000 ;
	    RECT 167.8000 38.2000 168.1000 43.8000 ;
	    RECT 167.8000 37.8000 168.2000 38.2000 ;
	    RECT 124.6000 28.8000 125.0000 29.2000 ;
	    RECT 124.6000 25.2000 124.9000 28.8000 ;
	    RECT 137.4000 27.8000 137.8000 28.2000 ;
	    RECT 137.4000 27.2000 137.7000 27.8000 ;
	    RECT 137.4000 26.8000 137.8000 27.2000 ;
	    RECT 148.6000 26.8000 149.0000 27.2000 ;
	    RECT 153.4000 27.1000 153.8000 27.2000 ;
	    RECT 154.2000 27.1000 154.6000 27.2000 ;
	    RECT 153.4000 26.8000 154.6000 27.1000 ;
	    RECT 148.6000 26.2000 148.9000 26.8000 ;
	    RECT 148.6000 25.8000 149.0000 26.2000 ;
	    RECT 124.6000 24.8000 125.0000 25.2000 ;
	    RECT 154.2000 16.2000 154.5000 26.8000 ;
	    RECT 154.2000 15.8000 154.6000 16.2000 ;
	    RECT 157.4000 16.1000 157.8000 16.2000 ;
	    RECT 158.2000 16.1000 158.6000 16.2000 ;
	    RECT 157.4000 15.8000 158.6000 16.1000 ;
         LAYER metal3 ;
	    RECT 144.6000 54.1000 145.0000 54.2000 ;
	    RECT 151.8000 54.1000 152.2000 54.2000 ;
	    RECT 144.6000 53.8000 152.2000 54.1000 ;
	    RECT 151.8000 53.2000 152.1000 53.8000 ;
	    RECT 151.8000 52.8000 152.2000 53.2000 ;
	    RECT 172.6000 47.1000 173.0000 47.2000 ;
	    RECT 175.8000 47.1000 176.2000 47.2000 ;
	    RECT 172.6000 46.8000 176.2000 47.1000 ;
	    RECT 167.8000 44.1000 168.2000 44.2000 ;
	    RECT 172.6000 44.1000 173.0000 44.2000 ;
	    RECT 167.8000 43.8000 173.0000 44.1000 ;
	    RECT 151.8000 38.1000 152.2000 38.2000 ;
	    RECT 167.8000 38.1000 168.2000 38.2000 ;
	    RECT 151.8000 37.8000 168.2000 38.1000 ;
	    RECT 124.6000 29.1000 125.0000 29.2000 ;
	    RECT 124.6000 28.8000 137.7000 29.1000 ;
	    RECT 137.4000 28.2000 137.7000 28.8000 ;
	    RECT 137.4000 28.1000 137.8000 28.2000 ;
	    RECT 137.4000 27.8000 148.9000 28.1000 ;
	    RECT 148.6000 27.2000 148.9000 27.8000 ;
	    RECT 148.6000 27.1000 149.0000 27.2000 ;
	    RECT 151.8000 27.1000 152.2000 27.2000 ;
	    RECT 153.4000 27.1000 153.8000 27.2000 ;
	    RECT 148.6000 26.8000 153.8000 27.1000 ;
	    RECT 154.2000 16.1000 154.6000 16.2000 ;
	    RECT 157.4000 16.1000 157.8000 16.2000 ;
	    RECT 154.2000 15.8000 157.8000 16.1000 ;
         LAYER metal4 ;
	    RECT 151.8000 53.8000 152.2000 54.2000 ;
	    RECT 151.8000 38.2000 152.1000 53.8000 ;
	    RECT 172.6000 46.8000 173.0000 47.2000 ;
	    RECT 172.6000 44.2000 172.9000 46.8000 ;
	    RECT 172.6000 43.8000 173.0000 44.2000 ;
	    RECT 151.8000 37.8000 152.2000 38.2000 ;
	    RECT 151.8000 27.2000 152.1000 37.8000 ;
	    RECT 151.8000 26.8000 152.2000 27.2000 ;
      END
   END SEL_B[7]
   PIN SEL_B[6]
      PORT
         LAYER metal1 ;
	    RECT 162.2000 44.8000 162.6000 45.6000 ;
	    RECT 136.6000 35.4000 137.0000 36.2000 ;
	    RECT 152.6000 33.4000 153.0000 34.2000 ;
	    RECT 134.2000 24.8000 134.6000 25.6000 ;
	    RECT 151.0000 24.8000 151.4000 25.6000 ;
         LAYER metal2 ;
	    RECT 162.2000 44.8000 162.6000 45.2000 ;
	    RECT 170.2000 44.8000 170.6000 45.2000 ;
	    RECT 162.2000 37.2000 162.5000 44.8000 ;
	    RECT 170.2000 37.2000 170.5000 44.8000 ;
	    RECT 162.2000 36.8000 162.6000 37.2000 ;
	    RECT 170.2000 36.8000 170.6000 37.2000 ;
	    RECT 162.2000 36.2000 162.5000 36.8000 ;
	    RECT 136.6000 36.1000 137.0000 36.2000 ;
	    RECT 137.4000 36.1000 137.8000 36.2000 ;
	    RECT 136.6000 35.8000 137.8000 36.1000 ;
	    RECT 152.6000 35.8000 153.0000 36.2000 ;
	    RECT 162.2000 35.8000 162.6000 36.2000 ;
	    RECT 136.6000 33.2000 136.9000 35.8000 ;
	    RECT 152.6000 34.2000 152.9000 35.8000 ;
	    RECT 152.6000 33.8000 153.0000 34.2000 ;
	    RECT 134.2000 32.8000 134.6000 33.2000 ;
	    RECT 136.6000 32.8000 137.0000 33.2000 ;
	    RECT 134.2000 25.2000 134.5000 32.8000 ;
	    RECT 152.6000 26.2000 152.9000 33.8000 ;
	    RECT 151.0000 25.8000 151.4000 26.2000 ;
	    RECT 152.6000 25.8000 153.0000 26.2000 ;
	    RECT 151.0000 25.2000 151.3000 25.8000 ;
	    RECT 134.2000 24.8000 134.6000 25.2000 ;
	    RECT 151.0000 24.8000 151.4000 25.2000 ;
         LAYER metal3 ;
	    RECT 170.2000 45.1000 170.6000 45.2000 ;
	    RECT 175.8000 45.1000 176.2000 45.2000 ;
	    RECT 170.2000 44.8000 176.2000 45.1000 ;
	    RECT 162.2000 37.1000 162.6000 37.2000 ;
	    RECT 170.2000 37.1000 170.6000 37.2000 ;
	    RECT 162.2000 36.8000 170.6000 37.1000 ;
	    RECT 137.4000 36.1000 137.8000 36.2000 ;
	    RECT 152.6000 36.1000 153.0000 36.2000 ;
	    RECT 162.2000 36.1000 162.6000 36.2000 ;
	    RECT 137.4000 35.8000 162.6000 36.1000 ;
	    RECT 134.2000 33.1000 134.6000 33.2000 ;
	    RECT 136.6000 33.1000 137.0000 33.2000 ;
	    RECT 134.2000 32.8000 137.0000 33.1000 ;
	    RECT 151.0000 26.1000 151.4000 26.2000 ;
	    RECT 152.6000 26.1000 153.0000 26.2000 ;
	    RECT 151.0000 25.8000 153.0000 26.1000 ;
      END
   END SEL_B[6]
   PIN SEL_B[5]
      PORT
         LAYER metal1 ;
	    RECT 12.6000 25.8000 13.0000 26.6000 ;
	    RECT 19.8000 25.8000 20.2000 26.6000 ;
	    RECT 28.6000 25.8000 29.0000 26.6000 ;
	    RECT 29.4000 14.4000 29.8000 15.2000 ;
	    RECT 19.8000 5.8000 20.2000 6.6000 ;
         LAYER metal2 ;
	    RECT 11.8000 26.1000 12.2000 26.2000 ;
	    RECT 12.6000 26.1000 13.0000 26.2000 ;
	    RECT 11.8000 25.8000 13.0000 26.1000 ;
	    RECT 19.0000 26.1000 19.4000 26.2000 ;
	    RECT 19.8000 26.1000 20.2000 26.2000 ;
	    RECT 19.0000 25.8000 20.2000 26.1000 ;
	    RECT 27.8000 26.1000 28.2000 26.2000 ;
	    RECT 28.6000 26.1000 29.0000 26.2000 ;
	    RECT 27.8000 25.8000 29.0000 26.1000 ;
	    RECT 29.4000 25.8000 29.8000 26.2000 ;
	    RECT 29.4000 15.2000 29.7000 25.8000 ;
	    RECT 29.4000 14.8000 29.8000 15.2000 ;
	    RECT 29.4000 6.2000 29.7000 14.8000 ;
	    RECT 19.8000 6.1000 20.2000 6.2000 ;
	    RECT 20.6000 6.1000 21.0000 6.2000 ;
	    RECT 19.8000 5.8000 21.0000 6.1000 ;
	    RECT 29.4000 5.8000 29.8000 6.2000 ;
	    RECT 29.4000 -1.8000 29.7000 5.8000 ;
	    RECT 29.4000 -2.2000 29.8000 -1.8000 ;
         LAYER metal3 ;
	    RECT 11.8000 26.1000 12.2000 26.2000 ;
	    RECT 19.0000 26.1000 19.4000 26.2000 ;
	    RECT 27.8000 26.1000 28.2000 26.2000 ;
	    RECT 29.4000 26.1000 29.8000 26.2000 ;
	    RECT 11.8000 25.8000 29.8000 26.1000 ;
	    RECT 20.6000 6.1000 21.0000 6.2000 ;
	    RECT 29.4000 6.1000 29.8000 6.2000 ;
	    RECT 20.6000 5.8000 29.8000 6.1000 ;
      END
   END SEL_B[5]
   PIN SEL_B[4]
      PORT
         LAYER metal1 ;
	    RECT 17.4000 44.8000 17.8000 45.6000 ;
	    RECT 32.6000 45.1000 33.0000 45.6000 ;
	    RECT 33.4000 45.1000 33.8000 45.2000 ;
	    RECT 32.6000 44.8000 33.8000 45.1000 ;
	    RECT 19.8000 33.4000 20.2000 34.2000 ;
	    RECT 14.2000 15.4000 14.6000 16.2000 ;
	    RECT 23.0000 15.4000 23.4000 16.2000 ;
	    RECT 2.2000 13.4000 2.6000 14.2000 ;
	    RECT 20.6000 13.4000 21.0000 14.2000 ;
	    RECT 4.6000 7.1000 5.0000 7.2000 ;
	    RECT 5.4000 7.1000 5.8000 7.6000 ;
	    RECT 4.6000 6.8000 5.8000 7.1000 ;
	    RECT 19.0000 6.8000 19.4000 7.6000 ;
         LAYER metal2 ;
	    RECT 17.4000 45.1000 17.8000 45.2000 ;
	    RECT 18.2000 45.1000 18.6000 45.2000 ;
	    RECT 17.4000 44.8000 18.6000 45.1000 ;
	    RECT 20.6000 44.8000 21.0000 45.2000 ;
	    RECT 32.6000 45.1000 33.0000 45.2000 ;
	    RECT 33.4000 45.1000 33.8000 45.2000 ;
	    RECT 32.6000 44.8000 33.8000 45.1000 ;
	    RECT 19.8000 34.1000 20.2000 34.2000 ;
	    RECT 20.6000 34.1000 20.9000 44.8000 ;
	    RECT 19.8000 33.8000 20.9000 34.1000 ;
	    RECT 20.6000 18.2000 20.9000 33.8000 ;
	    RECT 2.2000 17.8000 2.6000 18.2000 ;
	    RECT 14.2000 17.8000 14.6000 18.2000 ;
	    RECT 20.6000 17.8000 21.0000 18.2000 ;
	    RECT 2.2000 16.2000 2.5000 17.8000 ;
	    RECT 14.2000 16.2000 14.5000 17.8000 ;
	    RECT 20.6000 16.2000 20.9000 17.8000 ;
	    RECT 2.2000 15.8000 2.6000 16.2000 ;
	    RECT 14.2000 15.8000 14.6000 16.2000 ;
	    RECT 20.6000 15.8000 21.0000 16.2000 ;
	    RECT 23.0000 16.1000 23.4000 16.2000 ;
	    RECT 23.8000 16.1000 24.2000 16.2000 ;
	    RECT 23.0000 15.8000 24.2000 16.1000 ;
	    RECT 2.2000 14.2000 2.5000 15.8000 ;
	    RECT 20.6000 14.2000 20.9000 15.8000 ;
	    RECT 2.2000 13.8000 2.6000 14.2000 ;
	    RECT 20.6000 13.8000 21.0000 14.2000 ;
	    RECT 2.2000 8.2000 2.5000 13.8000 ;
	    RECT 2.2000 7.8000 2.6000 8.2000 ;
	    RECT 4.6000 7.8000 5.0000 8.2000 ;
	    RECT 4.6000 7.2000 4.9000 7.8000 ;
	    RECT 20.6000 7.2000 20.9000 13.8000 ;
	    RECT 4.6000 6.8000 5.0000 7.2000 ;
	    RECT 19.0000 7.1000 19.4000 7.2000 ;
	    RECT 19.8000 7.1000 20.2000 7.2000 ;
	    RECT 19.0000 6.8000 20.2000 7.1000 ;
	    RECT 20.6000 6.8000 21.0000 7.2000 ;
         LAYER metal3 ;
	    RECT 18.2000 45.1000 18.6000 45.2000 ;
	    RECT 20.6000 45.1000 21.0000 45.2000 ;
	    RECT 32.6000 45.1000 33.0000 45.2000 ;
	    RECT 18.2000 44.8000 33.0000 45.1000 ;
	    RECT 2.2000 18.1000 2.6000 18.2000 ;
	    RECT 14.2000 18.1000 14.6000 18.2000 ;
	    RECT 20.6000 18.1000 21.0000 18.2000 ;
	    RECT 2.2000 17.8000 21.0000 18.1000 ;
	    RECT -2.6000 16.1000 -2.2000 16.2000 ;
	    RECT 2.2000 16.1000 2.6000 16.2000 ;
	    RECT -2.6000 15.8000 2.6000 16.1000 ;
	    RECT 20.6000 16.1000 21.0000 16.2000 ;
	    RECT 23.8000 16.1000 24.2000 16.2000 ;
	    RECT 20.6000 15.8000 24.2000 16.1000 ;
	    RECT 2.2000 8.1000 2.6000 8.2000 ;
	    RECT 4.6000 8.1000 5.0000 8.2000 ;
	    RECT 2.2000 7.8000 5.0000 8.1000 ;
	    RECT 19.8000 7.1000 20.2000 7.2000 ;
	    RECT 20.6000 7.1000 21.0000 7.2000 ;
	    RECT 19.8000 6.8000 21.0000 7.1000 ;
      END
   END SEL_B[4]
   PIN SEL_B[3]
      PORT
         LAYER metal1 ;
	    RECT 29.4000 44.8000 29.8000 45.6000 ;
	    RECT 10.2000 24.8000 10.6000 25.6000 ;
	    RECT 13.4000 24.8000 13.8000 25.6000 ;
	    RECT 16.6000 24.8000 17.0000 25.6000 ;
	    RECT 13.4000 13.4000 13.8000 14.2000 ;
         LAYER metal2 ;
	    RECT 29.4000 44.8000 29.8000 45.2000 ;
	    RECT 29.4000 41.2000 29.7000 44.8000 ;
	    RECT 13.4000 40.8000 13.8000 41.2000 ;
	    RECT 29.4000 40.8000 29.8000 41.2000 ;
	    RECT 13.4000 25.2000 13.7000 40.8000 ;
	    RECT 10.2000 24.8000 10.6000 25.2000 ;
	    RECT 13.4000 24.8000 13.8000 25.2000 ;
	    RECT 15.8000 25.1000 16.2000 25.2000 ;
	    RECT 16.6000 25.1000 17.0000 25.2000 ;
	    RECT 15.8000 24.8000 17.0000 25.1000 ;
	    RECT 10.2000 24.2000 10.5000 24.8000 ;
	    RECT 13.4000 24.2000 13.7000 24.8000 ;
	    RECT 10.2000 23.8000 10.6000 24.2000 ;
	    RECT 13.4000 23.8000 13.8000 24.2000 ;
	    RECT 13.4000 14.2000 13.7000 23.8000 ;
	    RECT 13.4000 13.8000 13.8000 14.2000 ;
         LAYER metal3 ;
	    RECT 13.4000 41.1000 13.8000 41.2000 ;
	    RECT 29.4000 41.1000 29.8000 41.2000 ;
	    RECT 13.4000 40.8000 29.8000 41.1000 ;
	    RECT -2.6000 25.1000 -2.2000 25.2000 ;
	    RECT 10.2000 25.1000 10.6000 25.2000 ;
	    RECT -2.6000 24.8000 10.6000 25.1000 ;
	    RECT 13.4000 25.1000 13.8000 25.2000 ;
	    RECT 15.8000 25.1000 16.2000 25.2000 ;
	    RECT 13.4000 24.8000 16.2000 25.1000 ;
	    RECT 10.2000 24.1000 10.6000 24.2000 ;
	    RECT 13.4000 24.1000 13.8000 24.2000 ;
	    RECT 10.2000 23.8000 13.8000 24.1000 ;
      END
   END SEL_B[3]
   PIN SEL_B[2]
      PORT
         LAYER metal1 ;
	    RECT 115.0000 54.4000 115.4000 55.2000 ;
	    RECT 123.0000 54.4000 123.4000 55.2000 ;
	    RECT 111.8000 26.1000 112.2000 26.6000 ;
	    RECT 112.6000 26.1000 113.0000 26.2000 ;
	    RECT 111.8000 25.8000 113.0000 26.1000 ;
	    RECT 128.6000 14.4000 129.0000 15.2000 ;
	    RECT 121.4000 6.1000 121.8000 6.6000 ;
	    RECT 122.2000 6.1000 122.6000 6.2000 ;
	    RECT 121.4000 5.8000 122.6000 6.1000 ;
         LAYER metal2 ;
	    RECT 115.0000 55.1000 115.4000 55.2000 ;
	    RECT 115.8000 55.1000 116.2000 55.2000 ;
	    RECT 115.0000 54.8000 116.2000 55.1000 ;
	    RECT 122.2000 55.1000 122.6000 55.2000 ;
	    RECT 123.0000 55.1000 123.4000 55.2000 ;
	    RECT 122.2000 54.8000 123.4000 55.1000 ;
	    RECT 112.6000 26.8000 113.0000 27.2000 ;
	    RECT 112.6000 26.2000 112.9000 26.8000 ;
	    RECT 112.6000 25.8000 113.0000 26.2000 ;
	    RECT 127.8000 15.1000 128.2000 15.2000 ;
	    RECT 128.6000 15.1000 129.0000 15.2000 ;
	    RECT 127.8000 14.8000 129.0000 15.1000 ;
	    RECT 122.2000 5.8000 122.6000 6.2000 ;
	    RECT 122.2000 1.2000 122.5000 5.8000 ;
	    RECT 122.2000 0.8000 122.6000 1.2000 ;
	    RECT 123.8000 0.8000 124.2000 1.2000 ;
	    RECT 123.8000 -1.8000 124.1000 0.8000 ;
	    RECT 123.8000 -2.2000 124.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 115.8000 55.1000 116.2000 55.2000 ;
	    RECT 119.8000 55.1000 120.2000 55.2000 ;
	    RECT 122.2000 55.1000 122.6000 55.2000 ;
	    RECT 115.8000 54.8000 122.6000 55.1000 ;
	    RECT 112.6000 26.8000 113.0000 27.2000 ;
	    RECT 112.6000 26.1000 112.9000 26.8000 ;
	    RECT 119.8000 26.1000 120.2000 26.2000 ;
	    RECT 112.6000 25.8000 120.2000 26.1000 ;
	    RECT 119.8000 15.1000 120.2000 15.2000 ;
	    RECT 127.8000 15.1000 128.2000 15.2000 ;
	    RECT 128.6000 15.1000 129.0000 15.2000 ;
	    RECT 119.8000 14.8000 129.0000 15.1000 ;
	    RECT 122.2000 1.1000 122.6000 1.2000 ;
	    RECT 123.8000 1.1000 124.2000 1.2000 ;
	    RECT 128.6000 1.1000 129.0000 1.2000 ;
	    RECT 122.2000 0.8000 129.0000 1.1000 ;
         LAYER metal4 ;
	    RECT 119.8000 54.8000 120.2000 55.2000 ;
	    RECT 119.8000 26.2000 120.1000 54.8000 ;
	    RECT 119.8000 25.8000 120.2000 26.2000 ;
	    RECT 119.8000 15.2000 120.1000 25.8000 ;
	    RECT 119.8000 14.8000 120.2000 15.2000 ;
	    RECT 128.6000 14.8000 129.0000 15.2000 ;
	    RECT 128.6000 1.2000 128.9000 14.8000 ;
	    RECT 128.6000 0.8000 129.0000 1.2000 ;
      END
   END SEL_B[2]
   PIN SEL_B[1]
      PORT
         LAYER metal1 ;
	    RECT 103.8000 46.8000 104.2000 47.6000 ;
	    RECT 113.4000 46.8000 113.8000 47.6000 ;
	    RECT 115.8000 44.8000 116.2000 45.6000 ;
	    RECT 125.4000 44.8000 125.8000 45.6000 ;
	    RECT 118.2000 26.8000 118.6000 27.6000 ;
	    RECT 125.4000 26.8000 125.8000 27.6000 ;
	    RECT 103.8000 15.4000 104.2000 16.2000 ;
	    RECT 115.0000 15.4000 115.4000 16.2000 ;
	    RECT 102.2000 6.8000 102.6000 7.6000 ;
         LAYER metal2 ;
	    RECT 103.0000 47.1000 103.4000 47.2000 ;
	    RECT 103.8000 47.1000 104.2000 47.2000 ;
	    RECT 103.0000 46.8000 104.2000 47.1000 ;
	    RECT 113.4000 46.8000 113.8000 47.2000 ;
	    RECT 113.4000 45.2000 113.7000 46.8000 ;
	    RECT 113.4000 44.8000 113.8000 45.2000 ;
	    RECT 115.0000 45.1000 115.4000 45.2000 ;
	    RECT 115.8000 45.1000 116.2000 45.2000 ;
	    RECT 115.0000 44.8000 116.2000 45.1000 ;
	    RECT 124.6000 45.1000 125.0000 45.2000 ;
	    RECT 125.4000 45.1000 125.8000 45.2000 ;
	    RECT 124.6000 44.8000 125.8000 45.1000 ;
	    RECT 115.0000 27.2000 115.3000 44.8000 ;
	    RECT 115.0000 26.8000 115.4000 27.2000 ;
	    RECT 117.4000 27.1000 117.8000 27.2000 ;
	    RECT 118.2000 27.1000 118.6000 27.2000 ;
	    RECT 117.4000 26.8000 118.6000 27.1000 ;
	    RECT 125.4000 27.1000 125.8000 27.2000 ;
	    RECT 126.2000 27.1000 126.6000 27.2000 ;
	    RECT 125.4000 26.8000 126.6000 27.1000 ;
	    RECT 117.4000 18.2000 117.7000 26.8000 ;
	    RECT 115.0000 17.8000 115.4000 18.2000 ;
	    RECT 117.4000 17.8000 117.8000 18.2000 ;
	    RECT 115.0000 16.2000 115.3000 17.8000 ;
	    RECT 102.2000 15.8000 102.6000 16.2000 ;
	    RECT 103.8000 16.1000 104.2000 16.2000 ;
	    RECT 104.6000 16.1000 105.0000 16.2000 ;
	    RECT 103.8000 15.8000 105.0000 16.1000 ;
	    RECT 115.0000 15.8000 115.4000 16.2000 ;
	    RECT 102.2000 7.2000 102.5000 15.8000 ;
	    RECT 102.2000 6.8000 102.6000 7.2000 ;
	    RECT 102.2000 2.2000 102.5000 6.8000 ;
	    RECT 102.2000 1.8000 102.6000 2.2000 ;
	    RECT 103.8000 1.8000 104.2000 2.2000 ;
	    RECT 103.8000 -1.8000 104.1000 1.8000 ;
	    RECT 103.8000 -2.2000 104.2000 -1.8000 ;
         LAYER metal3 ;
	    RECT 103.0000 47.1000 103.4000 47.2000 ;
	    RECT 113.4000 47.1000 113.8000 47.2000 ;
	    RECT 103.0000 46.8000 113.8000 47.1000 ;
	    RECT 113.4000 45.1000 113.8000 45.2000 ;
	    RECT 115.0000 45.1000 115.4000 45.2000 ;
	    RECT 124.6000 45.1000 125.0000 45.2000 ;
	    RECT 113.4000 44.8000 125.0000 45.1000 ;
	    RECT 115.0000 27.1000 115.4000 27.2000 ;
	    RECT 117.4000 27.1000 117.8000 27.2000 ;
	    RECT 126.2000 27.1000 126.6000 27.2000 ;
	    RECT 115.0000 26.8000 126.6000 27.1000 ;
	    RECT 115.0000 18.1000 115.4000 18.2000 ;
	    RECT 117.4000 18.1000 117.8000 18.2000 ;
	    RECT 115.0000 17.8000 117.8000 18.1000 ;
	    RECT 102.2000 16.1000 102.6000 16.2000 ;
	    RECT 104.6000 16.1000 105.0000 16.2000 ;
	    RECT 115.0000 16.1000 115.4000 16.2000 ;
	    RECT 102.2000 15.8000 115.4000 16.1000 ;
	    RECT 102.2000 2.1000 102.6000 2.2000 ;
	    RECT 103.8000 2.1000 104.2000 2.2000 ;
	    RECT 102.2000 1.8000 104.2000 2.1000 ;
      END
   END SEL_B[1]
   PIN SEL_B[0]
      PORT
         LAYER metal1 ;
	    RECT 122.2000 45.1000 122.6000 45.6000 ;
	    RECT 123.0000 45.1000 123.4000 45.2000 ;
	    RECT 122.2000 44.8000 123.4000 45.1000 ;
	    RECT 123.0000 33.4000 123.4000 34.2000 ;
	    RECT 99.0000 25.1000 99.4000 25.6000 ;
	    RECT 99.8000 25.1000 100.2000 25.6000 ;
	    RECT 99.0000 24.8000 100.2000 25.1000 ;
	    RECT 107.0000 25.1000 107.4000 25.6000 ;
	    RECT 107.8000 25.1000 108.2000 25.2000 ;
	    RECT 107.0000 24.8000 108.2000 25.1000 ;
         LAYER metal2 ;
	    RECT 123.0000 44.8000 123.4000 45.2000 ;
	    RECT 123.0000 34.2000 123.3000 44.8000 ;
	    RECT 123.0000 33.8000 123.4000 34.2000 ;
	    RECT 123.0000 33.2000 123.3000 33.8000 ;
	    RECT 108.6000 32.8000 109.0000 33.2000 ;
	    RECT 123.0000 32.8000 123.4000 33.2000 ;
	    RECT 108.6000 27.1000 108.9000 32.8000 ;
	    RECT 107.8000 26.8000 108.9000 27.1000 ;
	    RECT 107.8000 25.2000 108.1000 26.8000 ;
	    RECT 99.8000 25.1000 100.2000 25.2000 ;
	    RECT 100.6000 25.1000 101.0000 25.2000 ;
	    RECT 99.8000 24.8000 101.0000 25.1000 ;
	    RECT 107.8000 24.8000 108.2000 25.2000 ;
	    RECT 110.2000 1.8000 110.6000 2.2000 ;
	    RECT 110.2000 -1.8000 110.5000 1.8000 ;
	    RECT 110.2000 -2.2000 110.6000 -1.8000 ;
         LAYER metal3 ;
	    RECT 108.6000 33.1000 109.0000 33.2000 ;
	    RECT 123.0000 33.1000 123.4000 33.2000 ;
	    RECT 108.6000 32.8000 123.4000 33.1000 ;
	    RECT 100.6000 25.1000 101.0000 25.2000 ;
	    RECT 107.8000 25.1000 108.2000 25.2000 ;
	    RECT 109.4000 25.1000 109.8000 25.2000 ;
	    RECT 100.6000 24.8000 109.8000 25.1000 ;
	    RECT 109.4000 2.1000 109.8000 2.2000 ;
	    RECT 110.2000 2.1000 110.6000 2.2000 ;
	    RECT 109.4000 1.8000 110.6000 2.1000 ;
         LAYER metal4 ;
	    RECT 109.4000 24.8000 109.8000 25.2000 ;
	    RECT 109.4000 2.2000 109.7000 24.8000 ;
	    RECT 109.4000 1.8000 109.8000 2.2000 ;
      END
   END SEL_B[0]
   OBS
         LAYER metal1 ;
	    RECT 1.4000 156.1000 1.8000 159.9000 ;
	    RECT 2.2000 156.1000 2.6000 156.6000 ;
	    RECT 1.4000 155.8000 2.6000 156.1000 ;
	    RECT 1.4000 151.1000 1.8000 155.8000 ;
	    RECT 3.0000 153.1000 3.4000 159.9000 ;
	    RECT 3.8000 154.1000 4.2000 154.2000 ;
	    RECT 4.6000 154.1000 5.0000 154.2000 ;
	    RECT 3.8000 153.8000 5.0000 154.1000 ;
	    RECT 3.8000 153.4000 4.2000 153.8000 ;
	    RECT 4.6000 153.4000 5.0000 153.8000 ;
	    RECT 2.5000 152.8000 3.4000 153.1000 ;
	    RECT 5.4000 153.1000 5.8000 159.9000 ;
	    RECT 7.0000 154.1000 7.4000 159.9000 ;
	    RECT 9.9000 156.2000 10.3000 159.9000 ;
	    RECT 10.6000 156.8000 11.0000 157.2000 ;
	    RECT 10.7000 156.2000 11.0000 156.8000 ;
	    RECT 9.9000 155.9000 10.4000 156.2000 ;
	    RECT 10.7000 155.9000 11.4000 156.2000 ;
	    RECT 9.4000 154.4000 9.8000 155.2000 ;
	    RECT 10.1000 154.2000 10.4000 155.9000 ;
	    RECT 11.0000 155.8000 11.4000 155.9000 ;
	    RECT 11.0000 155.1000 11.3000 155.8000 ;
	    RECT 12.6000 155.1000 13.0000 159.9000 ;
	    RECT 11.0000 154.8000 13.0000 155.1000 ;
	    RECT 8.6000 154.1000 9.0000 154.2000 ;
	    RECT 10.1000 154.1000 11.4000 154.2000 ;
	    RECT 11.8000 154.1000 12.2000 154.2000 ;
	    RECT 7.0000 153.8000 9.4000 154.1000 ;
	    RECT 10.1000 153.8000 12.2000 154.1000 ;
	    RECT 5.4000 152.8000 6.3000 153.1000 ;
	    RECT 2.5000 152.2000 2.9000 152.8000 ;
	    RECT 2.2000 151.8000 2.9000 152.2000 ;
	    RECT 2.5000 151.1000 2.9000 151.8000 ;
	    RECT 5.9000 152.2000 6.3000 152.8000 ;
	    RECT 5.9000 151.8000 6.6000 152.2000 ;
	    RECT 5.9000 151.1000 6.3000 151.8000 ;
	    RECT 7.0000 151.1000 7.4000 153.8000 ;
	    RECT 9.0000 153.6000 9.4000 153.8000 ;
	    RECT 8.7000 153.1000 10.5000 153.3000 ;
	    RECT 11.0000 153.1000 11.3000 153.8000 ;
	    RECT 12.6000 153.1000 13.0000 154.8000 ;
	    RECT 13.4000 153.4000 13.8000 154.2000 ;
	    RECT 14.2000 153.4000 14.6000 154.2000 ;
	    RECT 8.6000 153.0000 10.6000 153.1000 ;
	    RECT 8.6000 151.1000 9.0000 153.0000 ;
	    RECT 10.2000 151.1000 10.6000 153.0000 ;
	    RECT 11.0000 151.1000 11.4000 153.1000 ;
	    RECT 12.1000 152.8000 13.0000 153.1000 ;
	    RECT 15.0000 153.1000 15.4000 159.9000 ;
	    RECT 16.6000 155.9000 17.0000 159.9000 ;
	    RECT 18.2000 156.2000 18.6000 159.9000 ;
	    RECT 17.5000 155.9000 18.6000 156.2000 ;
	    RECT 16.6000 154.8000 16.9000 155.9000 ;
	    RECT 17.5000 155.6000 17.8000 155.9000 ;
	    RECT 17.2000 155.2000 17.8000 155.6000 ;
	    RECT 15.8000 154.1000 16.2000 154.2000 ;
	    RECT 16.6000 154.1000 17.0000 154.8000 ;
	    RECT 15.8000 153.8000 17.0000 154.1000 ;
	    RECT 15.0000 152.8000 15.9000 153.1000 ;
	    RECT 12.1000 151.1000 12.5000 152.8000 ;
	    RECT 15.5000 152.2000 15.9000 152.8000 ;
	    RECT 15.0000 151.8000 15.9000 152.2000 ;
	    RECT 15.5000 151.1000 15.9000 151.8000 ;
	    RECT 16.6000 151.1000 17.0000 153.8000 ;
	    RECT 17.5000 153.7000 17.8000 155.2000 ;
	    RECT 17.5000 153.4000 18.6000 153.7000 ;
	    RECT 19.0000 153.4000 19.4000 154.2000 ;
	    RECT 18.2000 151.1000 18.6000 153.4000 ;
	    RECT 19.8000 153.1000 20.2000 159.9000 ;
	    RECT 21.4000 153.4000 21.8000 154.2000 ;
	    RECT 22.2000 153.1000 22.6000 159.9000 ;
	    RECT 23.0000 156.1000 23.4000 156.6000 ;
	    RECT 23.8000 156.1000 24.2000 159.9000 ;
	    RECT 23.0000 155.8000 24.2000 156.1000 ;
	    RECT 19.8000 152.8000 20.7000 153.1000 ;
	    RECT 22.2000 152.8000 23.1000 153.1000 ;
	    RECT 20.3000 152.2000 20.7000 152.8000 ;
	    RECT 22.7000 152.2000 23.1000 152.8000 ;
	    RECT 20.3000 151.8000 21.0000 152.2000 ;
	    RECT 22.2000 151.8000 23.1000 152.2000 ;
	    RECT 20.3000 151.1000 20.7000 151.8000 ;
	    RECT 22.7000 151.1000 23.1000 151.8000 ;
	    RECT 23.8000 151.1000 24.2000 155.8000 ;
	    RECT 25.4000 153.4000 25.8000 154.2000 ;
	    RECT 26.2000 153.1000 26.6000 159.9000 ;
	    RECT 27.8000 154.1000 28.2000 154.2000 ;
	    RECT 28.6000 154.1000 29.0000 159.9000 ;
	    RECT 27.8000 153.8000 29.0000 154.1000 ;
	    RECT 26.2000 152.8000 27.1000 153.1000 ;
	    RECT 26.7000 152.2000 27.1000 152.8000 ;
	    RECT 26.7000 151.8000 27.4000 152.2000 ;
	    RECT 26.7000 151.1000 27.1000 151.8000 ;
	    RECT 28.6000 151.1000 29.0000 153.8000 ;
	    RECT 29.4000 151.1000 29.8000 159.9000 ;
	    RECT 31.8000 151.1000 32.2000 159.9000 ;
	    RECT 33.9000 156.2000 34.3000 159.9000 ;
	    RECT 34.6000 156.8000 35.0000 157.2000 ;
	    RECT 34.7000 156.2000 35.0000 156.8000 ;
	    RECT 33.9000 155.9000 34.4000 156.2000 ;
	    RECT 34.7000 155.9000 35.4000 156.2000 ;
	    RECT 33.4000 154.4000 33.8000 155.2000 ;
	    RECT 34.1000 154.2000 34.4000 155.9000 ;
	    RECT 35.0000 155.8000 35.4000 155.9000 ;
	    RECT 35.0000 155.1000 35.3000 155.8000 ;
	    RECT 36.6000 155.1000 37.0000 159.9000 ;
	    RECT 35.0000 154.8000 37.0000 155.1000 ;
	    RECT 32.6000 154.1000 33.0000 154.2000 ;
	    RECT 34.1000 154.1000 35.4000 154.2000 ;
	    RECT 35.8000 154.1000 36.2000 154.2000 ;
	    RECT 32.6000 153.8000 33.4000 154.1000 ;
	    RECT 34.1000 153.8000 36.2000 154.1000 ;
	    RECT 33.0000 153.6000 33.4000 153.8000 ;
	    RECT 32.7000 153.1000 34.5000 153.3000 ;
	    RECT 35.0000 153.1000 35.3000 153.8000 ;
	    RECT 36.6000 153.1000 37.0000 154.8000 ;
	    RECT 37.4000 153.4000 37.8000 154.2000 ;
	    RECT 39.0000 153.1000 39.4000 159.9000 ;
	    RECT 40.6000 155.9000 41.0000 159.9000 ;
	    RECT 42.2000 156.2000 42.6000 159.9000 ;
	    RECT 41.5000 155.9000 42.6000 156.2000 ;
	    RECT 40.6000 154.8000 40.9000 155.9000 ;
	    RECT 41.5000 155.6000 41.8000 155.9000 ;
	    RECT 41.2000 155.2000 41.8000 155.6000 ;
	    RECT 39.8000 153.4000 40.2000 154.2000 ;
	    RECT 32.6000 153.0000 34.6000 153.1000 ;
	    RECT 32.6000 151.1000 33.0000 153.0000 ;
	    RECT 34.2000 151.1000 34.6000 153.0000 ;
	    RECT 35.0000 151.1000 35.4000 153.1000 ;
	    RECT 36.1000 152.8000 37.0000 153.1000 ;
	    RECT 38.5000 152.8000 39.4000 153.1000 ;
	    RECT 36.1000 151.1000 36.5000 152.8000 ;
	    RECT 38.5000 152.2000 38.9000 152.8000 ;
	    RECT 38.5000 151.8000 39.4000 152.2000 ;
	    RECT 38.5000 151.1000 38.9000 151.8000 ;
	    RECT 40.6000 151.1000 41.0000 154.8000 ;
	    RECT 41.5000 153.7000 41.8000 155.2000 ;
	    RECT 41.5000 153.4000 42.6000 153.7000 ;
	    RECT 43.0000 153.4000 43.4000 154.2000 ;
	    RECT 42.2000 151.1000 42.6000 153.4000 ;
	    RECT 43.8000 153.1000 44.2000 159.9000 ;
	    RECT 45.4000 153.4000 45.8000 154.2000 ;
	    RECT 46.2000 153.1000 46.6000 159.9000 ;
	    RECT 47.0000 156.1000 47.4000 156.6000 ;
	    RECT 47.8000 156.1000 48.2000 159.9000 ;
	    RECT 47.0000 155.8000 48.2000 156.1000 ;
	    RECT 49.4000 155.8000 49.8000 156.6000 ;
	    RECT 43.8000 152.8000 44.7000 153.1000 ;
	    RECT 46.2000 152.8000 47.1000 153.1000 ;
	    RECT 44.3000 152.2000 44.7000 152.8000 ;
	    RECT 43.8000 151.8000 44.7000 152.2000 ;
	    RECT 44.3000 151.1000 44.7000 151.8000 ;
	    RECT 46.7000 152.2000 47.1000 152.8000 ;
	    RECT 46.7000 151.8000 47.4000 152.2000 ;
	    RECT 46.7000 151.1000 47.1000 151.8000 ;
	    RECT 47.8000 151.1000 48.2000 155.8000 ;
	    RECT 50.2000 153.1000 50.6000 159.9000 ;
	    RECT 51.8000 153.4000 52.2000 154.2000 ;
	    RECT 49.7000 152.8000 50.6000 153.1000 ;
	    RECT 52.6000 153.1000 53.0000 159.9000 ;
	    RECT 54.2000 156.2000 54.6000 159.9000 ;
	    RECT 54.2000 155.9000 55.3000 156.2000 ;
	    RECT 55.8000 155.9000 56.2000 159.9000 ;
	    RECT 55.0000 155.6000 55.3000 155.9000 ;
	    RECT 55.0000 155.2000 55.6000 155.6000 ;
	    RECT 55.0000 153.7000 55.3000 155.2000 ;
	    RECT 55.9000 154.8000 56.2000 155.9000 ;
	    RECT 54.2000 153.4000 55.3000 153.7000 ;
	    RECT 52.6000 152.8000 53.5000 153.1000 ;
	    RECT 49.7000 152.2000 50.1000 152.8000 ;
	    RECT 53.1000 152.2000 53.5000 152.8000 ;
	    RECT 49.7000 151.8000 50.6000 152.2000 ;
	    RECT 53.1000 151.8000 53.8000 152.2000 ;
	    RECT 49.7000 151.1000 50.1000 151.8000 ;
	    RECT 53.1000 151.1000 53.5000 151.8000 ;
	    RECT 54.2000 151.1000 54.6000 153.4000 ;
	    RECT 55.8000 151.1000 56.2000 154.8000 ;
	    RECT 57.4000 154.1000 57.8000 159.9000 ;
	    RECT 59.5000 156.2000 59.9000 159.9000 ;
	    RECT 60.2000 156.8000 60.6000 157.2000 ;
	    RECT 60.3000 156.2000 60.6000 156.8000 ;
	    RECT 59.5000 155.9000 60.0000 156.2000 ;
	    RECT 60.3000 156.1000 61.0000 156.2000 ;
	    RECT 61.4000 156.1000 61.8000 156.2000 ;
	    RECT 60.3000 155.9000 61.8000 156.1000 ;
	    RECT 59.0000 154.4000 59.4000 155.2000 ;
	    RECT 59.7000 155.1000 60.0000 155.9000 ;
	    RECT 60.6000 155.8000 61.8000 155.9000 ;
	    RECT 62.2000 155.1000 62.6000 155.2000 ;
	    RECT 59.7000 154.8000 62.6000 155.1000 ;
	    RECT 59.7000 154.2000 60.0000 154.8000 ;
	    RECT 58.2000 154.1000 58.6000 154.2000 ;
	    RECT 57.4000 153.8000 59.0000 154.1000 ;
	    RECT 59.7000 153.8000 61.0000 154.2000 ;
	    RECT 61.4000 154.1000 61.8000 154.2000 ;
	    RECT 63.8000 154.1000 64.2000 159.9000 ;
	    RECT 61.4000 153.8000 64.2000 154.1000 ;
	    RECT 57.4000 151.1000 57.8000 153.8000 ;
	    RECT 58.6000 153.6000 59.0000 153.8000 ;
	    RECT 58.3000 153.1000 60.1000 153.3000 ;
	    RECT 60.6000 153.1000 60.9000 153.8000 ;
	    RECT 63.8000 153.1000 64.2000 153.8000 ;
	    RECT 64.6000 154.1000 65.0000 154.2000 ;
	    RECT 65.4000 154.1000 65.8000 154.2000 ;
	    RECT 64.6000 153.8000 65.8000 154.1000 ;
	    RECT 64.6000 153.4000 65.0000 153.8000 ;
	    RECT 65.4000 153.4000 65.8000 153.8000 ;
	    RECT 58.2000 153.0000 60.2000 153.1000 ;
	    RECT 58.2000 151.1000 58.6000 153.0000 ;
	    RECT 59.8000 151.1000 60.2000 153.0000 ;
	    RECT 60.6000 151.1000 61.0000 153.1000 ;
	    RECT 63.3000 152.8000 64.2000 153.1000 ;
	    RECT 66.2000 153.1000 66.6000 159.9000 ;
	    RECT 67.0000 156.1000 67.4000 156.6000 ;
	    RECT 67.8000 156.1000 68.2000 159.9000 ;
	    RECT 67.0000 155.8000 68.2000 156.1000 ;
	    RECT 69.4000 155.8000 69.8000 156.6000 ;
	    RECT 66.2000 152.8000 67.1000 153.1000 ;
	    RECT 63.3000 151.1000 63.7000 152.8000 ;
	    RECT 66.7000 152.2000 67.1000 152.8000 ;
	    RECT 66.2000 151.8000 67.1000 152.2000 ;
	    RECT 66.7000 151.1000 67.1000 151.8000 ;
	    RECT 67.8000 151.1000 68.2000 155.8000 ;
	    RECT 70.2000 153.1000 70.6000 159.9000 ;
	    RECT 71.8000 153.4000 72.2000 154.2000 ;
	    RECT 69.7000 152.8000 70.6000 153.1000 ;
	    RECT 72.6000 153.1000 73.0000 159.9000 ;
	    RECT 73.4000 156.1000 73.8000 156.6000 ;
	    RECT 74.2000 156.1000 74.6000 159.9000 ;
	    RECT 73.4000 155.8000 74.6000 156.1000 ;
	    RECT 76.1000 156.3000 76.5000 159.9000 ;
	    RECT 76.1000 155.9000 77.0000 156.3000 ;
	    RECT 72.6000 152.8000 73.5000 153.1000 ;
	    RECT 69.7000 152.2000 70.1000 152.8000 ;
	    RECT 69.4000 151.8000 70.1000 152.2000 ;
	    RECT 69.7000 151.1000 70.1000 151.8000 ;
	    RECT 73.1000 152.2000 73.5000 152.8000 ;
	    RECT 73.1000 151.8000 73.8000 152.2000 ;
	    RECT 73.1000 151.1000 73.5000 151.8000 ;
	    RECT 74.2000 151.1000 74.6000 155.8000 ;
	    RECT 75.8000 154.8000 76.2000 155.6000 ;
	    RECT 76.6000 154.2000 76.9000 155.9000 ;
	    RECT 78.2000 155.8000 78.6000 156.6000 ;
	    RECT 76.6000 153.8000 77.0000 154.2000 ;
	    RECT 75.8000 153.1000 76.2000 153.2000 ;
	    RECT 76.6000 153.1000 76.9000 153.8000 ;
	    RECT 75.8000 152.8000 76.9000 153.1000 ;
	    RECT 76.6000 152.1000 76.9000 152.8000 ;
	    RECT 77.4000 152.4000 77.8000 153.2000 ;
	    RECT 79.0000 153.1000 79.4000 159.9000 ;
	    RECT 80.6000 155.6000 81.0000 159.9000 ;
	    RECT 82.7000 157.9000 83.3000 159.9000 ;
	    RECT 85.0000 157.9000 85.4000 159.9000 ;
	    RECT 87.2000 158.2000 87.6000 159.9000 ;
	    RECT 87.2000 157.9000 88.2000 158.2000 ;
	    RECT 83.0000 157.5000 83.4000 157.9000 ;
	    RECT 85.1000 157.6000 85.4000 157.9000 ;
	    RECT 84.7000 157.3000 86.5000 157.6000 ;
	    RECT 87.8000 157.5000 88.2000 157.9000 ;
	    RECT 84.7000 157.2000 85.1000 157.3000 ;
	    RECT 86.1000 157.2000 86.5000 157.3000 ;
	    RECT 82.6000 156.6000 83.3000 157.0000 ;
	    RECT 83.0000 156.1000 83.3000 156.6000 ;
	    RECT 84.1000 156.5000 85.2000 156.8000 ;
	    RECT 84.1000 156.4000 84.5000 156.5000 ;
	    RECT 83.0000 155.8000 84.2000 156.1000 ;
	    RECT 80.6000 155.3000 82.7000 155.6000 ;
	    RECT 79.8000 154.1000 80.2000 154.2000 ;
	    RECT 80.6000 154.1000 81.0000 155.3000 ;
	    RECT 82.3000 155.2000 82.7000 155.3000 ;
	    RECT 81.5000 154.9000 81.9000 155.0000 ;
	    RECT 81.5000 154.6000 83.4000 154.9000 ;
	    RECT 83.0000 154.5000 83.4000 154.6000 ;
	    RECT 79.8000 153.8000 81.0000 154.1000 ;
	    RECT 83.9000 154.2000 84.2000 155.8000 ;
	    RECT 84.9000 155.9000 85.2000 156.5000 ;
	    RECT 85.5000 156.5000 85.9000 156.6000 ;
	    RECT 87.8000 156.5000 88.2000 156.6000 ;
	    RECT 85.5000 156.2000 88.2000 156.5000 ;
	    RECT 84.9000 155.7000 87.3000 155.9000 ;
	    RECT 89.4000 155.7000 89.8000 159.9000 ;
	    RECT 84.9000 155.6000 89.8000 155.7000 ;
	    RECT 86.9000 155.5000 89.8000 155.6000 ;
	    RECT 87.0000 155.4000 89.8000 155.5000 ;
	    RECT 86.2000 155.1000 86.6000 155.2000 ;
	    RECT 90.2000 155.1000 90.6000 159.9000 ;
	    RECT 93.1000 155.9000 94.1000 159.9000 ;
	    RECT 97.1000 156.2000 98.1000 159.9000 ;
	    RECT 100.1000 156.3000 100.5000 159.9000 ;
	    RECT 97.1000 155.9000 98.6000 156.2000 ;
	    RECT 100.1000 155.9000 101.0000 156.3000 ;
	    RECT 86.2000 154.8000 88.7000 155.1000 ;
	    RECT 87.0000 154.7000 87.4000 154.8000 ;
	    RECT 88.3000 154.7000 88.7000 154.8000 ;
	    RECT 90.2000 154.8000 92.1000 155.1000 ;
	    RECT 87.5000 154.2000 87.9000 154.3000 ;
	    RECT 83.9000 153.9000 89.4000 154.2000 ;
	    RECT 84.1000 153.8000 84.5000 153.9000 ;
	    RECT 79.8000 153.4000 80.2000 153.8000 ;
	    RECT 80.6000 153.6000 81.0000 153.8000 ;
	    RECT 78.5000 152.8000 79.4000 153.1000 ;
	    RECT 80.6000 153.3000 82.6000 153.6000 ;
	    RECT 78.5000 152.2000 78.9000 152.8000 ;
	    RECT 76.6000 151.1000 77.0000 152.1000 ;
	    RECT 78.5000 151.8000 79.4000 152.2000 ;
	    RECT 78.5000 151.1000 78.9000 151.8000 ;
	    RECT 80.6000 151.1000 81.0000 153.3000 ;
	    RECT 82.1000 153.2000 82.6000 153.3000 ;
	    RECT 82.2000 153.1000 82.6000 153.2000 ;
	    RECT 83.8000 153.1000 84.2000 153.2000 ;
	    RECT 82.2000 152.8000 84.2000 153.1000 ;
	    RECT 87.0000 152.8000 87.3000 153.9000 ;
	    RECT 88.6000 153.8000 89.4000 153.9000 ;
	    RECT 86.1000 152.7000 86.5000 152.8000 ;
	    RECT 83.0000 152.1000 83.4000 152.5000 ;
	    RECT 85.1000 152.4000 86.5000 152.7000 ;
	    RECT 87.0000 152.4000 87.4000 152.8000 ;
	    RECT 85.1000 152.1000 85.4000 152.4000 ;
	    RECT 87.8000 152.1000 88.2000 152.5000 ;
	    RECT 82.7000 151.8000 83.4000 152.1000 ;
	    RECT 82.7000 151.1000 83.3000 151.8000 ;
	    RECT 85.0000 151.1000 85.4000 152.1000 ;
	    RECT 87.2000 151.8000 88.2000 152.1000 ;
	    RECT 87.2000 151.1000 87.6000 151.8000 ;
	    RECT 89.4000 151.1000 89.8000 153.5000 ;
	    RECT 90.2000 151.1000 90.6000 154.8000 ;
	    RECT 91.8000 154.2000 92.1000 154.8000 ;
	    RECT 92.6000 154.4000 93.0000 155.2000 ;
	    RECT 93.4000 154.2000 93.7000 155.9000 ;
	    RECT 97.4000 155.8000 98.6000 155.9000 ;
	    RECT 94.2000 154.4000 94.6000 155.2000 ;
	    RECT 91.0000 153.4000 91.4000 154.2000 ;
	    RECT 91.8000 154.1000 92.2000 154.2000 ;
	    RECT 93.4000 154.1000 93.8000 154.2000 ;
	    RECT 91.8000 153.8000 92.6000 154.1000 ;
	    RECT 93.4000 153.8000 94.6000 154.1000 ;
	    RECT 95.0000 153.8000 95.4000 154.6000 ;
	    RECT 96.6000 154.4000 97.0000 155.2000 ;
	    RECT 97.4000 154.2000 97.7000 155.8000 ;
	    RECT 98.2000 154.4000 98.6000 155.2000 ;
	    RECT 99.8000 154.8000 100.2000 155.6000 ;
	    RECT 95.8000 154.1000 96.2000 154.2000 ;
	    RECT 97.4000 154.1000 97.8000 154.2000 ;
	    RECT 99.0000 154.1000 99.4000 154.6000 ;
	    RECT 100.6000 154.2000 100.9000 155.9000 ;
	    RECT 99.8000 154.1000 100.2000 154.2000 ;
	    RECT 95.8000 153.8000 96.6000 154.1000 ;
	    RECT 97.4000 153.8000 98.6000 154.1000 ;
	    RECT 99.0000 153.8000 100.2000 154.1000 ;
	    RECT 100.6000 154.1000 101.0000 154.2000 ;
	    RECT 102.2000 154.1000 102.6000 154.2000 ;
	    RECT 100.6000 153.8000 102.6000 154.1000 ;
	    RECT 92.2000 153.6000 92.6000 153.8000 ;
	    RECT 91.9000 153.1000 93.7000 153.3000 ;
	    RECT 94.3000 153.1000 94.6000 153.8000 ;
	    RECT 96.2000 153.6000 96.6000 153.8000 ;
	    RECT 95.9000 153.1000 97.7000 153.3000 ;
	    RECT 98.3000 153.1000 98.6000 153.8000 ;
	    RECT 91.8000 153.0000 93.8000 153.1000 ;
	    RECT 91.8000 151.1000 92.2000 153.0000 ;
	    RECT 93.4000 151.4000 93.8000 153.0000 ;
	    RECT 94.2000 151.7000 94.6000 153.1000 ;
	    RECT 95.0000 151.4000 95.4000 153.1000 ;
	    RECT 93.4000 151.1000 95.4000 151.4000 ;
	    RECT 95.8000 153.0000 97.8000 153.1000 ;
	    RECT 95.8000 151.1000 96.2000 153.0000 ;
	    RECT 97.4000 151.4000 97.8000 153.0000 ;
	    RECT 98.2000 151.7000 98.6000 153.1000 ;
	    RECT 99.0000 151.4000 99.4000 153.1000 ;
	    RECT 97.4000 151.1000 99.4000 151.4000 ;
	    RECT 100.6000 152.1000 100.9000 153.8000 ;
	    RECT 102.2000 153.4000 102.6000 153.8000 ;
	    RECT 101.4000 152.4000 101.8000 153.2000 ;
	    RECT 103.0000 153.1000 103.4000 159.9000 ;
	    RECT 103.8000 156.1000 104.2000 156.6000 ;
	    RECT 104.6000 156.1000 105.0000 159.9000 ;
	    RECT 103.8000 155.8000 105.0000 156.1000 ;
	    RECT 105.4000 156.2000 105.8000 159.9000 ;
	    RECT 107.0000 156.2000 107.4000 159.9000 ;
	    RECT 105.4000 155.9000 107.4000 156.2000 ;
	    RECT 107.8000 155.8000 108.2000 156.6000 ;
	    RECT 104.7000 155.2000 105.0000 155.8000 ;
	    RECT 106.6000 155.2000 107.0000 155.4000 ;
	    RECT 104.6000 154.9000 105.8000 155.2000 ;
	    RECT 106.6000 155.1000 107.4000 155.2000 ;
	    RECT 108.6000 155.1000 109.0000 159.9000 ;
	    RECT 110.5000 156.3000 110.9000 159.9000 ;
	    RECT 106.6000 154.9000 109.0000 155.1000 ;
	    RECT 104.6000 154.8000 105.0000 154.9000 ;
	    RECT 103.0000 152.8000 103.9000 153.1000 ;
	    RECT 104.6000 152.8000 105.0000 153.2000 ;
	    RECT 105.5000 153.1000 105.8000 154.9000 ;
	    RECT 107.0000 154.8000 109.0000 154.9000 ;
	    RECT 109.4000 155.8000 109.8000 156.2000 ;
	    RECT 110.5000 155.9000 111.4000 156.3000 ;
	    RECT 115.0000 156.1000 115.4000 159.9000 ;
	    RECT 115.8000 156.8000 116.2000 157.2000 ;
	    RECT 115.8000 156.1000 116.1000 156.8000 ;
	    RECT 109.4000 155.1000 109.7000 155.8000 ;
	    RECT 110.2000 155.1000 110.6000 155.6000 ;
	    RECT 109.4000 154.8000 110.6000 155.1000 ;
	    RECT 106.2000 153.8000 106.6000 154.6000 ;
	    RECT 108.6000 153.1000 109.0000 154.8000 ;
	    RECT 111.0000 154.2000 111.3000 155.9000 ;
	    RECT 115.0000 155.8000 116.1000 156.1000 ;
	    RECT 109.4000 153.4000 109.8000 154.2000 ;
	    RECT 111.0000 154.1000 111.4000 154.2000 ;
	    RECT 113.4000 154.1000 113.8000 154.2000 ;
	    RECT 111.0000 153.8000 113.8000 154.1000 ;
	    RECT 103.5000 152.2000 103.9000 152.8000 ;
	    RECT 104.7000 152.4000 105.1000 152.8000 ;
	    RECT 100.6000 151.1000 101.0000 152.1000 ;
	    RECT 103.0000 151.8000 103.9000 152.2000 ;
	    RECT 103.5000 151.1000 103.9000 151.8000 ;
	    RECT 105.4000 151.1000 105.8000 153.1000 ;
	    RECT 108.1000 152.8000 109.0000 153.1000 ;
	    RECT 108.1000 151.1000 108.5000 152.8000 ;
	    RECT 111.0000 152.1000 111.3000 153.8000 ;
	    RECT 111.8000 152.4000 112.2000 153.2000 ;
	    RECT 113.4000 153.1000 113.8000 153.2000 ;
	    RECT 114.2000 153.1000 114.6000 153.2000 ;
	    RECT 113.4000 152.8000 114.6000 153.1000 ;
	    RECT 114.2000 152.4000 114.6000 152.8000 ;
	    RECT 111.0000 151.1000 111.4000 152.1000 ;
	    RECT 115.0000 151.1000 115.4000 155.8000 ;
	    RECT 115.8000 155.1000 116.2000 155.2000 ;
	    RECT 116.6000 155.1000 117.0000 159.9000 ;
	    RECT 117.4000 155.8000 117.8000 156.6000 ;
	    RECT 118.2000 156.2000 118.6000 159.9000 ;
	    RECT 119.8000 159.6000 121.8000 159.9000 ;
	    RECT 119.8000 156.2000 120.2000 159.6000 ;
	    RECT 118.2000 155.9000 120.2000 156.2000 ;
	    RECT 120.6000 155.9000 121.0000 159.3000 ;
	    RECT 121.4000 155.9000 121.8000 159.6000 ;
	    RECT 122.2000 156.9000 122.6000 159.9000 ;
	    RECT 122.3000 156.6000 122.6000 156.9000 ;
	    RECT 123.8000 159.6000 125.8000 159.9000 ;
	    RECT 123.8000 156.9000 124.2000 159.6000 ;
	    RECT 124.6000 156.9000 125.0000 159.3000 ;
	    RECT 125.4000 157.0000 125.8000 159.6000 ;
	    RECT 126.3000 159.6000 128.1000 159.9000 ;
	    RECT 126.3000 159.5000 126.6000 159.6000 ;
	    RECT 123.8000 156.6000 124.1000 156.9000 ;
	    RECT 122.3000 156.3000 124.1000 156.6000 ;
	    RECT 124.7000 156.7000 125.0000 156.9000 ;
	    RECT 126.2000 156.7000 126.6000 159.5000 ;
	    RECT 127.8000 159.5000 128.1000 159.6000 ;
	    RECT 124.7000 156.5000 126.6000 156.7000 ;
	    RECT 127.0000 156.5000 127.4000 159.3000 ;
	    RECT 127.8000 156.5000 128.2000 159.5000 ;
	    RECT 124.7000 156.4000 126.5000 156.5000 ;
	    RECT 127.0000 156.2000 127.3000 156.5000 ;
	    RECT 127.0000 156.1000 127.4000 156.2000 ;
	    RECT 120.6000 155.6000 120.9000 155.9000 ;
	    RECT 125.7000 155.8000 127.4000 156.1000 ;
	    RECT 118.6000 155.2000 119.0000 155.4000 ;
	    RECT 119.9000 155.3000 120.9000 155.6000 ;
	    RECT 119.9000 155.2000 120.2000 155.3000 ;
	    RECT 115.8000 154.8000 117.0000 155.1000 ;
	    RECT 118.2000 154.9000 119.0000 155.2000 ;
	    RECT 118.2000 154.8000 118.6000 154.9000 ;
	    RECT 119.8000 154.8000 120.2000 155.2000 ;
	    RECT 121.4000 155.1000 121.8000 155.6000 ;
	    RECT 122.2000 155.1000 122.6000 155.2000 ;
	    RECT 121.4000 154.8000 122.6000 155.1000 ;
	    RECT 124.6000 154.8000 125.4000 155.2000 ;
	    RECT 115.8000 153.4000 116.2000 154.2000 ;
	    RECT 116.6000 153.1000 117.0000 154.8000 ;
	    RECT 117.4000 154.1000 117.8000 154.2000 ;
	    RECT 119.0000 154.1000 119.4000 154.6000 ;
	    RECT 117.4000 153.8000 119.4000 154.1000 ;
	    RECT 119.9000 153.1000 120.2000 154.8000 ;
	    RECT 120.5000 154.4000 120.9000 154.8000 ;
	    RECT 120.6000 154.2000 120.9000 154.4000 ;
	    RECT 120.6000 154.1000 121.0000 154.2000 ;
	    RECT 121.4000 154.1000 121.8000 154.2000 ;
	    RECT 120.6000 153.8000 121.8000 154.1000 ;
	    RECT 123.8000 153.8000 124.6000 154.2000 ;
	    RECT 116.6000 152.8000 117.5000 153.1000 ;
	    RECT 117.1000 151.1000 117.5000 152.8000 ;
	    RECT 119.7000 152.2000 120.5000 153.1000 ;
	    RECT 123.0000 152.8000 123.9000 153.2000 ;
	    RECT 124.6000 153.1000 125.0000 153.2000 ;
	    RECT 125.7000 153.1000 126.0000 155.8000 ;
	    RECT 129.4000 155.1000 129.8000 159.9000 ;
	    RECT 130.6000 156.8000 131.0000 157.2000 ;
	    RECT 130.6000 156.2000 130.9000 156.8000 ;
	    RECT 131.3000 156.2000 131.7000 159.9000 ;
	    RECT 130.2000 155.9000 130.9000 156.2000 ;
	    RECT 131.2000 155.9000 131.7000 156.2000 ;
	    RECT 133.4000 155.9000 133.8000 159.9000 ;
	    RECT 134.2000 156.2000 134.6000 159.9000 ;
	    RECT 135.8000 156.2000 136.2000 159.9000 ;
	    RECT 137.0000 156.8000 137.4000 157.2000 ;
	    RECT 137.0000 156.2000 137.3000 156.8000 ;
	    RECT 137.7000 156.2000 138.1000 159.9000 ;
	    RECT 134.2000 155.9000 136.2000 156.2000 ;
	    RECT 136.6000 155.9000 137.3000 156.2000 ;
	    RECT 137.6000 155.9000 138.1000 156.2000 ;
	    RECT 140.1000 157.2000 140.5000 159.9000 ;
	    RECT 140.1000 156.8000 141.0000 157.2000 ;
	    RECT 140.1000 156.3000 140.5000 156.8000 ;
	    RECT 140.1000 155.9000 141.0000 156.3000 ;
	    RECT 142.2000 155.9000 142.6000 159.9000 ;
	    RECT 143.0000 156.2000 143.4000 159.9000 ;
	    RECT 144.6000 156.2000 145.0000 159.9000 ;
	    RECT 143.0000 155.9000 145.0000 156.2000 ;
	    RECT 130.2000 155.8000 130.6000 155.9000 ;
	    RECT 130.2000 155.1000 130.6000 155.2000 ;
	    RECT 129.4000 154.8000 130.6000 155.1000 ;
	    RECT 124.6000 152.8000 126.0000 153.1000 ;
	    RECT 125.7000 152.5000 126.0000 152.8000 ;
	    RECT 124.0000 152.2000 126.0000 152.5000 ;
	    RECT 128.6000 152.4000 129.0000 153.2000 ;
	    RECT 119.7000 151.8000 121.0000 152.2000 ;
	    RECT 124.0000 152.1000 124.3000 152.2000 ;
	    RECT 123.8000 151.8000 124.3000 152.1000 ;
	    RECT 125.4000 152.1000 126.0000 152.2000 ;
	    RECT 119.7000 151.1000 120.5000 151.8000 ;
	    RECT 123.8000 151.1000 124.2000 151.8000 ;
	    RECT 125.4000 151.1000 125.8000 152.1000 ;
	    RECT 129.4000 151.1000 129.8000 154.8000 ;
	    RECT 131.2000 154.2000 131.5000 155.9000 ;
	    RECT 133.5000 155.2000 133.8000 155.9000 ;
	    RECT 136.6000 155.8000 137.0000 155.9000 ;
	    RECT 135.4000 155.2000 135.8000 155.4000 ;
	    RECT 131.8000 154.4000 132.2000 155.2000 ;
	    RECT 133.4000 154.9000 134.6000 155.2000 ;
	    RECT 135.4000 155.1000 136.2000 155.2000 ;
	    RECT 137.6000 155.1000 137.9000 155.9000 ;
	    RECT 135.4000 154.9000 137.9000 155.1000 ;
	    RECT 133.4000 154.8000 133.8000 154.9000 ;
	    RECT 130.2000 153.8000 131.5000 154.2000 ;
	    RECT 132.6000 154.1000 133.0000 154.2000 ;
	    RECT 132.2000 153.8000 133.0000 154.1000 ;
	    RECT 130.3000 153.1000 130.6000 153.8000 ;
	    RECT 132.2000 153.6000 132.6000 153.8000 ;
	    RECT 131.1000 153.1000 132.9000 153.3000 ;
	    RECT 134.3000 153.2000 134.6000 154.9000 ;
	    RECT 135.8000 154.8000 137.9000 154.9000 ;
	    RECT 135.0000 153.8000 135.4000 154.6000 ;
	    RECT 137.6000 154.2000 137.9000 154.8000 ;
	    RECT 138.2000 154.4000 138.6000 155.2000 ;
	    RECT 139.8000 155.1000 140.2000 155.6000 ;
	    RECT 139.0000 154.8000 140.2000 155.1000 ;
	    RECT 136.6000 153.8000 137.9000 154.2000 ;
	    RECT 139.0000 154.2000 139.3000 154.8000 ;
	    RECT 140.6000 154.2000 140.9000 155.9000 ;
	    RECT 142.3000 155.2000 142.6000 155.9000 ;
	    RECT 145.4000 155.8000 145.8000 156.6000 ;
	    RECT 144.2000 155.2000 144.6000 155.4000 ;
	    RECT 142.2000 154.9000 143.4000 155.2000 ;
	    RECT 144.2000 154.9000 145.0000 155.2000 ;
	    RECT 142.2000 154.8000 142.6000 154.9000 ;
	    RECT 143.0000 154.8000 143.4000 154.9000 ;
	    RECT 144.6000 154.8000 145.0000 154.9000 ;
	    RECT 146.2000 155.1000 146.6000 159.9000 ;
	    RECT 148.6000 157.9000 149.0000 159.9000 ;
	    RECT 148.7000 157.8000 149.0000 157.9000 ;
	    RECT 150.2000 157.9000 150.6000 159.9000 ;
	    RECT 151.0000 157.9000 151.4000 159.9000 ;
	    RECT 150.2000 157.8000 150.5000 157.9000 ;
	    RECT 148.7000 157.5000 150.5000 157.8000 ;
	    RECT 150.2000 157.2000 150.5000 157.5000 ;
	    RECT 151.1000 157.8000 151.4000 157.9000 ;
	    RECT 152.6000 157.9000 153.0000 159.9000 ;
	    RECT 152.6000 157.8000 152.9000 157.9000 ;
	    RECT 151.1000 157.5000 152.9000 157.8000 ;
	    RECT 147.0000 157.1000 147.4000 157.2000 ;
	    RECT 149.4000 157.1000 149.8000 157.2000 ;
	    RECT 147.0000 156.8000 149.8000 157.1000 ;
	    RECT 149.4000 156.4000 149.8000 156.8000 ;
	    RECT 150.2000 156.8000 150.6000 157.2000 ;
	    RECT 150.2000 156.2000 150.5000 156.8000 ;
	    RECT 151.1000 156.2000 151.4000 157.5000 ;
	    RECT 151.8000 156.4000 152.2000 157.2000 ;
	    RECT 147.0000 155.8000 147.4000 156.2000 ;
	    RECT 147.0000 155.1000 147.3000 155.8000 ;
	    RECT 147.8000 155.4000 148.2000 156.2000 ;
	    RECT 150.2000 155.8000 150.6000 156.2000 ;
	    RECT 151.0000 155.8000 151.4000 156.2000 ;
	    RECT 146.2000 154.8000 147.3000 155.1000 ;
	    RECT 148.6000 154.8000 149.4000 155.2000 ;
	    RECT 139.0000 154.1000 139.4000 154.2000 ;
	    RECT 138.6000 153.8000 139.4000 154.1000 ;
	    RECT 140.6000 153.8000 141.0000 154.2000 ;
	    RECT 130.2000 151.1000 130.6000 153.1000 ;
	    RECT 131.0000 153.0000 133.0000 153.1000 ;
	    RECT 131.0000 151.1000 131.4000 153.0000 ;
	    RECT 132.6000 151.1000 133.0000 153.0000 ;
	    RECT 133.4000 152.8000 133.8000 153.2000 ;
	    RECT 133.5000 152.4000 133.9000 152.8000 ;
	    RECT 134.2000 151.1000 134.6000 153.2000 ;
	    RECT 136.7000 153.1000 137.0000 153.8000 ;
	    RECT 138.6000 153.6000 139.0000 153.8000 ;
	    RECT 137.5000 153.1000 139.3000 153.3000 ;
	    RECT 136.6000 151.1000 137.0000 153.1000 ;
	    RECT 137.4000 153.0000 139.4000 153.1000 ;
	    RECT 137.4000 151.1000 137.8000 153.0000 ;
	    RECT 139.0000 151.1000 139.4000 153.0000 ;
	    RECT 140.6000 152.1000 140.9000 153.8000 ;
	    RECT 141.4000 152.4000 141.8000 153.2000 ;
	    RECT 142.2000 152.8000 142.6000 153.2000 ;
	    RECT 143.1000 153.1000 143.4000 154.8000 ;
	    RECT 143.8000 153.8000 144.2000 154.6000 ;
	    RECT 146.2000 153.1000 146.6000 154.8000 ;
	    RECT 150.2000 154.2000 150.5000 155.8000 ;
	    RECT 147.0000 153.4000 147.4000 154.2000 ;
	    RECT 149.7000 154.1000 150.5000 154.2000 ;
	    RECT 149.6000 153.9000 150.5000 154.1000 ;
	    RECT 151.1000 154.2000 151.4000 155.8000 ;
	    RECT 153.4000 155.4000 153.8000 156.2000 ;
	    RECT 152.2000 154.8000 153.0000 155.2000 ;
	    RECT 151.1000 153.9000 152.2000 154.2000 ;
	    RECT 142.3000 152.4000 142.7000 152.8000 ;
	    RECT 140.6000 151.1000 141.0000 152.1000 ;
	    RECT 143.0000 151.1000 143.4000 153.1000 ;
	    RECT 145.7000 152.8000 146.6000 153.1000 ;
	    RECT 145.7000 151.1000 146.1000 152.8000 ;
	    RECT 149.6000 151.1000 150.0000 153.9000 ;
	    RECT 151.6000 153.8000 152.2000 153.9000 ;
	    RECT 151.6000 151.1000 152.0000 153.8000 ;
	    RECT 154.2000 153.4000 154.6000 154.2000 ;
	    RECT 155.0000 154.1000 155.4000 159.9000 ;
	    RECT 155.8000 155.8000 156.2000 156.6000 ;
	    RECT 157.9000 156.2000 158.3000 159.9000 ;
	    RECT 158.6000 156.8000 159.0000 157.2000 ;
	    RECT 158.7000 156.2000 159.0000 156.8000 ;
	    RECT 157.9000 155.9000 158.4000 156.2000 ;
	    RECT 158.7000 155.9000 159.4000 156.2000 ;
	    RECT 157.4000 154.4000 157.8000 155.2000 ;
	    RECT 158.1000 155.1000 158.4000 155.9000 ;
	    RECT 159.0000 155.8000 159.4000 155.9000 ;
	    RECT 159.0000 155.1000 159.4000 155.2000 ;
	    RECT 158.1000 154.8000 159.4000 155.1000 ;
	    RECT 158.1000 154.2000 158.4000 154.8000 ;
	    RECT 156.6000 154.1000 157.0000 154.2000 ;
	    RECT 155.0000 153.8000 157.4000 154.1000 ;
	    RECT 158.1000 153.8000 159.4000 154.2000 ;
	    RECT 155.0000 153.1000 155.4000 153.8000 ;
	    RECT 157.0000 153.6000 157.4000 153.8000 ;
	    RECT 156.7000 153.1000 158.5000 153.3000 ;
	    RECT 159.0000 153.1000 159.3000 153.8000 ;
	    RECT 159.8000 153.4000 160.2000 154.2000 ;
	    RECT 160.6000 153.1000 161.0000 159.9000 ;
	    RECT 161.4000 155.8000 161.8000 156.6000 ;
	    RECT 162.2000 155.7000 162.6000 159.9000 ;
	    RECT 164.4000 158.2000 164.8000 159.9000 ;
	    RECT 163.8000 157.9000 164.8000 158.2000 ;
	    RECT 166.6000 157.9000 167.0000 159.9000 ;
	    RECT 168.7000 157.9000 169.3000 159.9000 ;
	    RECT 163.8000 157.5000 164.2000 157.9000 ;
	    RECT 166.6000 157.6000 166.9000 157.9000 ;
	    RECT 165.5000 157.3000 167.3000 157.6000 ;
	    RECT 168.6000 157.5000 169.0000 157.9000 ;
	    RECT 165.5000 157.2000 165.9000 157.3000 ;
	    RECT 166.9000 157.2000 167.3000 157.3000 ;
	    RECT 163.8000 156.5000 164.2000 156.6000 ;
	    RECT 166.1000 156.5000 166.5000 156.6000 ;
	    RECT 163.8000 156.2000 166.5000 156.5000 ;
	    RECT 166.8000 156.5000 167.9000 156.8000 ;
	    RECT 166.8000 155.9000 167.1000 156.5000 ;
	    RECT 167.5000 156.4000 167.9000 156.5000 ;
	    RECT 168.7000 156.6000 169.4000 157.0000 ;
	    RECT 168.7000 156.1000 169.0000 156.6000 ;
	    RECT 164.7000 155.7000 167.1000 155.9000 ;
	    RECT 162.2000 155.6000 167.1000 155.7000 ;
	    RECT 167.8000 155.8000 169.0000 156.1000 ;
	    RECT 162.2000 155.5000 165.1000 155.6000 ;
	    RECT 162.2000 155.4000 165.0000 155.5000 ;
	    RECT 165.4000 155.1000 165.8000 155.2000 ;
	    RECT 163.3000 154.8000 165.8000 155.1000 ;
	    RECT 163.3000 154.7000 163.7000 154.8000 ;
	    RECT 164.6000 154.7000 165.0000 154.8000 ;
	    RECT 164.1000 154.2000 164.5000 154.3000 ;
	    RECT 167.8000 154.2000 168.1000 155.8000 ;
	    RECT 171.0000 155.6000 171.4000 159.9000 ;
	    RECT 169.3000 155.3000 171.4000 155.6000 ;
	    RECT 169.3000 155.2000 169.7000 155.3000 ;
	    RECT 170.1000 154.9000 170.5000 155.0000 ;
	    RECT 168.6000 154.6000 170.5000 154.9000 ;
	    RECT 168.6000 154.5000 169.0000 154.6000 ;
	    RECT 162.6000 153.9000 168.1000 154.2000 ;
	    RECT 162.6000 153.8000 163.4000 153.9000 ;
	    RECT 155.0000 152.8000 155.9000 153.1000 ;
	    RECT 155.5000 151.1000 155.9000 152.8000 ;
	    RECT 156.6000 153.0000 158.6000 153.1000 ;
	    RECT 156.6000 151.1000 157.0000 153.0000 ;
	    RECT 158.2000 151.1000 158.6000 153.0000 ;
	    RECT 159.0000 151.1000 159.4000 153.1000 ;
	    RECT 160.6000 152.8000 161.5000 153.1000 ;
	    RECT 161.1000 152.2000 161.5000 152.8000 ;
	    RECT 161.1000 151.8000 161.8000 152.2000 ;
	    RECT 161.1000 151.1000 161.5000 151.8000 ;
	    RECT 162.2000 151.1000 162.6000 153.5000 ;
	    RECT 164.7000 152.8000 165.0000 153.9000 ;
	    RECT 165.4000 153.8000 165.8000 153.9000 ;
	    RECT 167.5000 153.8000 167.9000 153.9000 ;
	    RECT 171.0000 153.6000 171.4000 155.3000 ;
	    RECT 169.4000 153.3000 171.4000 153.6000 ;
	    RECT 169.4000 153.2000 169.9000 153.3000 ;
	    RECT 167.8000 153.1000 168.2000 153.2000 ;
	    RECT 169.4000 153.1000 169.8000 153.2000 ;
	    RECT 167.8000 152.8000 169.8000 153.1000 ;
	    RECT 163.8000 152.1000 164.2000 152.5000 ;
	    RECT 164.6000 152.4000 165.0000 152.8000 ;
	    RECT 165.5000 152.7000 165.9000 152.8000 ;
	    RECT 165.5000 152.4000 166.9000 152.7000 ;
	    RECT 166.6000 152.1000 166.9000 152.4000 ;
	    RECT 168.6000 152.1000 169.0000 152.5000 ;
	    RECT 163.8000 151.8000 164.8000 152.1000 ;
	    RECT 164.4000 151.1000 164.8000 151.8000 ;
	    RECT 166.6000 151.1000 167.0000 152.1000 ;
	    RECT 168.6000 151.8000 169.3000 152.1000 ;
	    RECT 168.7000 151.1000 169.3000 151.8000 ;
	    RECT 171.0000 151.1000 171.4000 153.3000 ;
	    RECT 1.2000 147.1000 1.6000 149.9000 ;
	    RECT 0.7000 146.9000 1.6000 147.1000 ;
	    RECT 3.8000 147.9000 4.2000 149.9000 ;
	    RECT 5.4000 148.9000 5.8000 149.9000 ;
	    RECT 0.7000 146.8000 1.5000 146.9000 ;
	    RECT 0.7000 145.2000 1.0000 146.8000 ;
	    RECT 3.8000 146.2000 4.1000 147.9000 ;
	    RECT 5.4000 147.8000 5.7000 148.9000 ;
	    RECT 6.2000 147.8000 6.6000 148.6000 ;
	    RECT 7.0000 147.9000 7.4000 149.9000 ;
	    RECT 7.8000 148.0000 8.2000 149.9000 ;
	    RECT 9.4000 148.0000 9.8000 149.9000 ;
	    RECT 7.8000 147.9000 9.8000 148.0000 ;
	    RECT 4.5000 147.5000 5.7000 147.8000 ;
	    RECT 1.8000 145.8000 2.6000 146.2000 ;
	    RECT 3.8000 145.8000 4.2000 146.2000 ;
	    RECT 4.5000 146.0000 4.8000 147.5000 ;
	    RECT 7.1000 147.2000 7.4000 147.9000 ;
	    RECT 7.9000 147.7000 9.7000 147.9000 ;
	    RECT 9.0000 147.2000 9.4000 147.4000 ;
	    RECT 7.0000 146.8000 8.3000 147.2000 ;
	    RECT 9.0000 147.1000 9.8000 147.2000 ;
	    RECT 10.2000 147.1000 10.6000 149.9000 ;
	    RECT 11.8000 147.6000 12.2000 149.9000 ;
	    RECT 11.8000 147.3000 12.9000 147.6000 ;
	    RECT 9.0000 146.9000 10.6000 147.1000 ;
	    RECT 9.4000 146.8000 10.6000 146.9000 ;
	    RECT 7.0000 146.2000 7.3000 146.8000 ;
	    RECT 0.6000 144.8000 1.0000 145.2000 ;
	    RECT 3.0000 144.8000 3.4000 145.6000 ;
	    RECT 3.8000 145.1000 4.1000 145.8000 ;
	    RECT 4.5000 145.7000 4.9000 146.0000 ;
	    RECT 7.0000 145.8000 7.4000 146.2000 ;
	    RECT 4.5000 145.6000 6.6000 145.7000 ;
	    RECT 4.6000 145.4000 6.6000 145.6000 ;
	    RECT 3.8000 144.8000 4.5000 145.1000 ;
	    RECT 0.7000 143.5000 1.0000 144.8000 ;
	    RECT 1.4000 143.8000 1.8000 144.6000 ;
	    RECT 0.7000 143.2000 2.5000 143.5000 ;
	    RECT 0.7000 143.1000 1.0000 143.2000 ;
	    RECT 0.6000 141.1000 1.0000 143.1000 ;
	    RECT 2.2000 143.1000 2.5000 143.2000 ;
	    RECT 2.2000 141.1000 2.6000 143.1000 ;
	    RECT 4.1000 141.1000 4.5000 144.8000 ;
	    RECT 6.2000 141.1000 6.6000 145.4000 ;
	    RECT 7.0000 145.1000 7.4000 145.2000 ;
	    RECT 8.0000 145.1000 8.3000 146.8000 ;
	    RECT 8.6000 145.8000 9.0000 146.6000 ;
	    RECT 7.0000 144.8000 7.7000 145.1000 ;
	    RECT 8.0000 144.8000 8.5000 145.1000 ;
	    RECT 7.4000 144.2000 7.7000 144.8000 ;
	    RECT 7.4000 143.8000 7.8000 144.2000 ;
	    RECT 8.1000 141.1000 8.5000 144.8000 ;
	    RECT 10.2000 141.1000 10.6000 146.8000 ;
	    RECT 12.6000 145.8000 12.9000 147.3000 ;
	    RECT 13.4000 146.2000 13.8000 149.9000 ;
	    RECT 14.2000 147.9000 14.6000 149.9000 ;
	    RECT 15.0000 148.0000 15.4000 149.9000 ;
	    RECT 16.6000 148.0000 17.0000 149.9000 ;
	    RECT 15.0000 147.9000 17.0000 148.0000 ;
	    RECT 14.3000 147.2000 14.6000 147.9000 ;
	    RECT 15.1000 147.7000 16.9000 147.9000 ;
	    RECT 16.2000 147.2000 16.6000 147.4000 ;
	    RECT 14.2000 146.8000 15.5000 147.2000 ;
	    RECT 16.2000 146.9000 17.0000 147.2000 ;
	    RECT 16.6000 146.8000 17.0000 146.9000 ;
	    RECT 12.6000 145.4000 13.2000 145.8000 ;
	    RECT 12.6000 145.1000 12.9000 145.4000 ;
	    RECT 13.5000 145.1000 13.8000 146.2000 ;
	    RECT 11.8000 144.8000 12.9000 145.1000 ;
	    RECT 11.8000 141.1000 12.2000 144.8000 ;
	    RECT 13.4000 141.1000 13.8000 145.1000 ;
	    RECT 14.2000 145.1000 14.6000 145.2000 ;
	    RECT 15.2000 145.1000 15.5000 146.8000 ;
	    RECT 15.8000 145.8000 16.2000 146.6000 ;
	    RECT 14.2000 144.8000 14.9000 145.1000 ;
	    RECT 15.2000 144.8000 15.7000 145.1000 ;
	    RECT 14.6000 144.2000 14.9000 144.8000 ;
	    RECT 14.6000 143.8000 15.0000 144.2000 ;
	    RECT 15.3000 142.2000 15.7000 144.8000 ;
	    RECT 15.3000 141.8000 16.2000 142.2000 ;
	    RECT 15.3000 141.1000 15.7000 141.8000 ;
	    RECT 17.4000 141.1000 17.8000 149.9000 ;
	    RECT 19.0000 147.1000 19.4000 149.9000 ;
	    RECT 18.2000 146.8000 19.4000 147.1000 ;
	    RECT 22.4000 147.1000 22.8000 149.9000 ;
	    RECT 23.8000 147.9000 24.2000 149.9000 ;
	    RECT 25.4000 148.9000 25.8000 149.9000 ;
	    RECT 23.8000 147.2000 24.1000 147.9000 ;
	    RECT 25.4000 147.8000 25.7000 148.9000 ;
	    RECT 26.2000 147.8000 26.6000 148.6000 ;
	    RECT 27.0000 147.9000 27.4000 149.9000 ;
	    RECT 27.8000 148.0000 28.2000 149.9000 ;
	    RECT 29.4000 148.0000 29.8000 149.9000 ;
	    RECT 27.8000 147.9000 29.8000 148.0000 ;
	    RECT 24.5000 147.5000 25.7000 147.8000 ;
	    RECT 22.4000 146.9000 23.3000 147.1000 ;
	    RECT 22.5000 146.8000 23.3000 146.9000 ;
	    RECT 18.2000 146.2000 18.5000 146.8000 ;
	    RECT 18.2000 145.8000 18.6000 146.2000 ;
	    RECT 19.0000 141.1000 19.4000 146.8000 ;
	    RECT 21.4000 145.8000 22.2000 146.2000 ;
	    RECT 19.8000 145.1000 20.2000 145.2000 ;
	    RECT 20.6000 145.1000 21.0000 145.6000 ;
	    RECT 19.8000 144.8000 21.0000 145.1000 ;
	    RECT 23.0000 145.2000 23.3000 146.8000 ;
	    RECT 23.8000 146.8000 24.2000 147.2000 ;
	    RECT 23.8000 146.2000 24.1000 146.8000 ;
	    RECT 23.8000 145.8000 24.2000 146.2000 ;
	    RECT 24.5000 146.0000 24.8000 147.5000 ;
	    RECT 27.1000 147.2000 27.4000 147.9000 ;
	    RECT 27.9000 147.7000 29.7000 147.9000 ;
	    RECT 29.0000 147.2000 29.4000 147.4000 ;
	    RECT 27.0000 146.8000 28.3000 147.2000 ;
	    RECT 29.0000 146.9000 29.8000 147.2000 ;
	    RECT 29.4000 146.8000 29.8000 146.9000 ;
	    RECT 23.0000 144.8000 23.4000 145.2000 ;
	    RECT 23.8000 145.1000 24.1000 145.8000 ;
	    RECT 24.5000 145.7000 24.9000 146.0000 ;
	    RECT 24.5000 145.6000 26.6000 145.7000 ;
	    RECT 24.6000 145.4000 26.6000 145.6000 ;
	    RECT 23.8000 144.8000 24.5000 145.1000 ;
	    RECT 22.2000 143.8000 22.6000 144.6000 ;
	    RECT 23.0000 143.5000 23.3000 144.8000 ;
	    RECT 21.5000 143.2000 23.3000 143.5000 ;
	    RECT 21.5000 143.1000 21.8000 143.2000 ;
	    RECT 21.4000 141.1000 21.8000 143.1000 ;
	    RECT 23.0000 143.1000 23.3000 143.2000 ;
	    RECT 23.0000 141.1000 23.4000 143.1000 ;
	    RECT 24.1000 141.1000 24.5000 144.8000 ;
	    RECT 26.2000 141.1000 26.6000 145.4000 ;
	    RECT 27.0000 145.1000 27.4000 145.2000 ;
	    RECT 28.0000 145.1000 28.3000 146.8000 ;
	    RECT 28.6000 145.8000 29.0000 146.6000 ;
	    RECT 27.0000 144.8000 27.7000 145.1000 ;
	    RECT 28.0000 144.8000 28.5000 145.1000 ;
	    RECT 27.4000 144.2000 27.7000 144.8000 ;
	    RECT 27.4000 143.8000 27.8000 144.2000 ;
	    RECT 28.1000 142.2000 28.5000 144.8000 ;
	    RECT 28.1000 141.8000 29.0000 142.2000 ;
	    RECT 28.1000 141.1000 28.5000 141.8000 ;
	    RECT 30.2000 141.1000 30.6000 149.9000 ;
	    RECT 31.8000 147.9000 32.2000 149.9000 ;
	    RECT 32.6000 148.0000 33.0000 149.9000 ;
	    RECT 34.2000 148.0000 34.6000 149.9000 ;
	    RECT 32.6000 147.9000 34.6000 148.0000 ;
	    RECT 31.9000 147.2000 32.2000 147.9000 ;
	    RECT 32.7000 147.7000 34.5000 147.9000 ;
	    RECT 33.8000 147.2000 34.2000 147.4000 ;
	    RECT 31.8000 146.8000 33.1000 147.2000 ;
	    RECT 33.8000 147.1000 34.6000 147.2000 ;
	    RECT 35.0000 147.1000 35.4000 149.9000 ;
	    RECT 36.6000 148.0000 37.0000 149.9000 ;
	    RECT 38.2000 148.0000 38.6000 149.9000 ;
	    RECT 36.6000 147.9000 38.6000 148.0000 ;
	    RECT 39.0000 147.9000 39.4000 149.9000 ;
	    RECT 36.7000 147.7000 38.5000 147.9000 ;
	    RECT 37.0000 147.2000 37.4000 147.4000 ;
	    RECT 39.0000 147.2000 39.3000 147.9000 ;
	    RECT 33.8000 146.9000 35.4000 147.1000 ;
	    RECT 34.2000 146.8000 35.4000 146.9000 ;
	    RECT 35.8000 147.1000 36.2000 147.2000 ;
	    RECT 36.6000 147.1000 37.4000 147.2000 ;
	    RECT 35.8000 146.9000 37.4000 147.1000 ;
	    RECT 35.8000 146.8000 37.0000 146.9000 ;
	    RECT 38.1000 146.8000 39.4000 147.2000 ;
	    RECT 31.8000 145.1000 32.2000 145.2000 ;
	    RECT 32.8000 145.1000 33.1000 146.8000 ;
	    RECT 33.4000 145.8000 33.8000 146.6000 ;
	    RECT 31.8000 144.8000 32.5000 145.1000 ;
	    RECT 32.8000 144.8000 33.3000 145.1000 ;
	    RECT 32.2000 144.2000 32.5000 144.8000 ;
	    RECT 32.2000 143.8000 32.6000 144.2000 ;
	    RECT 32.9000 142.2000 33.3000 144.8000 ;
	    RECT 32.9000 141.8000 33.8000 142.2000 ;
	    RECT 32.9000 141.1000 33.3000 141.8000 ;
	    RECT 35.0000 141.1000 35.4000 146.8000 ;
	    RECT 37.4000 145.8000 37.8000 146.6000 ;
	    RECT 38.1000 145.1000 38.4000 146.8000 ;
	    RECT 39.8000 146.2000 40.2000 149.9000 ;
	    RECT 41.4000 147.6000 41.8000 149.9000 ;
	    RECT 40.7000 147.3000 41.8000 147.6000 ;
	    RECT 39.0000 145.1000 39.4000 145.2000 ;
	    RECT 37.9000 144.8000 38.4000 145.1000 ;
	    RECT 38.7000 144.8000 39.4000 145.1000 ;
	    RECT 39.8000 145.1000 40.1000 146.2000 ;
	    RECT 40.7000 145.8000 41.0000 147.3000 ;
	    RECT 40.4000 145.4000 41.0000 145.8000 ;
	    RECT 40.7000 145.1000 41.0000 145.4000 ;
	    RECT 43.0000 147.1000 43.4000 149.9000 ;
	    RECT 43.8000 148.0000 44.2000 149.9000 ;
	    RECT 45.4000 148.0000 45.8000 149.9000 ;
	    RECT 43.8000 147.9000 45.8000 148.0000 ;
	    RECT 46.2000 147.9000 46.6000 149.9000 ;
	    RECT 47.8000 148.9000 48.2000 149.9000 ;
	    RECT 43.9000 147.7000 45.7000 147.9000 ;
	    RECT 44.2000 147.2000 44.6000 147.4000 ;
	    RECT 46.2000 147.2000 46.5000 147.9000 ;
	    RECT 47.0000 147.8000 47.4000 148.6000 ;
	    RECT 47.9000 147.8000 48.2000 148.9000 ;
	    RECT 49.4000 147.9000 49.8000 149.9000 ;
	    RECT 47.9000 147.5000 49.1000 147.8000 ;
	    RECT 43.8000 147.1000 44.6000 147.2000 ;
	    RECT 43.0000 146.9000 44.6000 147.1000 ;
	    RECT 43.0000 146.8000 44.2000 146.9000 ;
	    RECT 45.3000 146.8000 46.6000 147.2000 ;
	    RECT 37.9000 142.2000 38.3000 144.8000 ;
	    RECT 38.7000 144.2000 39.0000 144.8000 ;
	    RECT 38.6000 143.8000 39.0000 144.2000 ;
	    RECT 37.4000 141.8000 38.3000 142.2000 ;
	    RECT 37.9000 141.1000 38.3000 141.8000 ;
	    RECT 39.8000 141.1000 40.2000 145.1000 ;
	    RECT 40.7000 144.8000 41.8000 145.1000 ;
	    RECT 41.4000 141.1000 41.8000 144.8000 ;
	    RECT 43.0000 141.1000 43.4000 146.8000 ;
	    RECT 44.6000 145.8000 45.0000 146.6000 ;
	    RECT 45.3000 145.1000 45.6000 146.8000 ;
	    RECT 48.8000 146.0000 49.1000 147.5000 ;
	    RECT 49.5000 146.2000 49.8000 147.9000 ;
	    RECT 48.7000 145.7000 49.1000 146.0000 ;
	    RECT 49.4000 146.1000 49.8000 146.2000 ;
	    RECT 50.2000 146.8000 50.6000 147.2000 ;
	    RECT 50.2000 146.1000 50.5000 146.8000 ;
	    RECT 49.4000 145.8000 50.5000 146.1000 ;
	    RECT 47.0000 145.6000 49.1000 145.7000 ;
	    RECT 47.0000 145.4000 49.0000 145.6000 ;
	    RECT 46.2000 145.1000 46.6000 145.2000 ;
	    RECT 45.1000 144.8000 45.6000 145.1000 ;
	    RECT 45.9000 144.8000 46.6000 145.1000 ;
	    RECT 45.1000 142.2000 45.5000 144.8000 ;
	    RECT 45.9000 144.2000 46.2000 144.8000 ;
	    RECT 45.8000 143.8000 46.2000 144.2000 ;
	    RECT 44.6000 141.8000 45.5000 142.2000 ;
	    RECT 45.1000 141.1000 45.5000 141.8000 ;
	    RECT 47.0000 141.1000 47.4000 145.4000 ;
	    RECT 49.5000 145.1000 49.8000 145.8000 ;
	    RECT 49.1000 144.8000 49.8000 145.1000 ;
	    RECT 49.1000 141.1000 49.5000 144.8000 ;
	    RECT 51.0000 141.1000 51.4000 149.9000 ;
	    RECT 52.4000 147.1000 52.8000 149.9000 ;
	    RECT 53.4000 147.8000 53.8000 148.2000 ;
	    RECT 53.4000 147.1000 53.7000 147.8000 ;
	    RECT 51.9000 146.8000 53.7000 147.1000 ;
	    RECT 51.9000 145.2000 52.2000 146.8000 ;
	    RECT 53.0000 145.8000 53.8000 146.2000 ;
	    RECT 51.8000 144.8000 52.2000 145.2000 ;
	    RECT 54.2000 145.1000 54.6000 145.6000 ;
	    RECT 55.0000 145.1000 55.4000 145.2000 ;
	    RECT 54.2000 144.8000 55.4000 145.1000 ;
	    RECT 51.9000 143.5000 52.2000 144.8000 ;
	    RECT 52.6000 143.8000 53.0000 144.6000 ;
	    RECT 51.9000 143.2000 53.7000 143.5000 ;
	    RECT 51.9000 143.1000 52.2000 143.2000 ;
	    RECT 51.8000 141.1000 52.2000 143.1000 ;
	    RECT 53.4000 143.1000 53.7000 143.2000 ;
	    RECT 53.4000 141.1000 53.8000 143.1000 ;
	    RECT 55.8000 141.1000 56.2000 149.9000 ;
	    RECT 57.2000 147.1000 57.6000 149.9000 ;
	    RECT 62.2000 148.9000 62.6000 149.9000 ;
	    RECT 60.6000 148.1000 61.0000 148.2000 ;
	    RECT 61.4000 148.1000 61.8000 148.6000 ;
	    RECT 60.6000 147.8000 61.8000 148.1000 ;
	    RECT 62.3000 147.8000 62.6000 148.9000 ;
	    RECT 63.8000 147.9000 64.2000 149.9000 ;
	    RECT 62.3000 147.5000 63.5000 147.8000 ;
	    RECT 56.7000 146.9000 57.6000 147.1000 ;
	    RECT 56.7000 146.8000 57.5000 146.9000 ;
	    RECT 56.7000 145.2000 57.0000 146.8000 ;
	    RECT 57.8000 145.8000 58.6000 146.2000 ;
	    RECT 63.2000 146.0000 63.5000 147.5000 ;
	    RECT 63.9000 147.2000 64.2000 147.9000 ;
	    RECT 63.8000 146.8000 64.2000 147.2000 ;
	    RECT 66.4000 147.2000 66.8000 149.9000 ;
	    RECT 66.4000 146.9000 67.4000 147.2000 ;
	    RECT 69.6000 147.1000 70.0000 149.9000 ;
	    RECT 69.6000 146.9000 70.5000 147.1000 ;
	    RECT 66.5000 146.8000 67.4000 146.9000 ;
	    RECT 69.7000 146.8000 70.5000 146.9000 ;
	    RECT 63.9000 146.2000 64.2000 146.8000 ;
	    RECT 63.1000 145.7000 63.5000 146.0000 ;
	    RECT 63.8000 145.8000 64.2000 146.2000 ;
	    RECT 65.4000 145.8000 66.2000 146.2000 ;
	    RECT 56.6000 144.8000 57.0000 145.2000 ;
	    RECT 56.7000 143.5000 57.0000 144.8000 ;
	    RECT 61.4000 145.6000 63.5000 145.7000 ;
	    RECT 61.4000 145.4000 63.4000 145.6000 ;
	    RECT 57.4000 143.8000 57.8000 144.6000 ;
	    RECT 56.7000 143.2000 58.5000 143.5000 ;
	    RECT 56.7000 143.1000 57.0000 143.2000 ;
	    RECT 56.6000 141.1000 57.0000 143.1000 ;
	    RECT 58.2000 143.1000 58.5000 143.2000 ;
	    RECT 58.2000 141.1000 58.6000 143.1000 ;
	    RECT 61.4000 141.1000 61.8000 145.4000 ;
	    RECT 63.9000 145.1000 64.2000 145.8000 ;
	    RECT 63.5000 144.8000 64.2000 145.1000 ;
	    RECT 64.6000 144.8000 65.0000 145.6000 ;
	    RECT 67.0000 145.2000 67.3000 146.8000 ;
	    RECT 68.6000 145.8000 69.4000 146.2000 ;
	    RECT 70.2000 145.2000 70.5000 146.8000 ;
	    RECT 67.0000 144.8000 67.4000 145.2000 ;
	    RECT 70.2000 144.8000 70.6000 145.2000 ;
	    RECT 63.5000 141.1000 63.9000 144.8000 ;
	    RECT 66.2000 143.8000 66.6000 144.6000 ;
	    RECT 67.0000 143.5000 67.3000 144.8000 ;
	    RECT 69.4000 143.8000 69.8000 144.6000 ;
	    RECT 70.2000 143.5000 70.5000 144.8000 ;
	    RECT 65.5000 143.2000 67.3000 143.5000 ;
	    RECT 65.5000 143.1000 65.8000 143.2000 ;
	    RECT 65.4000 141.1000 65.8000 143.1000 ;
	    RECT 67.0000 143.1000 67.3000 143.2000 ;
	    RECT 68.7000 143.2000 70.5000 143.5000 ;
	    RECT 68.7000 143.1000 69.0000 143.2000 ;
	    RECT 67.0000 141.1000 67.4000 143.1000 ;
	    RECT 68.6000 141.1000 69.0000 143.1000 ;
	    RECT 70.2000 143.1000 70.5000 143.2000 ;
	    RECT 70.2000 141.1000 70.6000 143.1000 ;
	    RECT 71.8000 141.1000 72.2000 149.9000 ;
	    RECT 74.2000 147.9000 74.6000 149.9000 ;
	    RECT 76.6000 148.9000 77.0000 149.9000 ;
	    RECT 74.9000 148.2000 75.3000 148.6000 ;
	    RECT 73.4000 146.4000 73.8000 147.2000 ;
	    RECT 72.6000 146.1000 73.0000 146.2000 ;
	    RECT 74.2000 146.1000 74.5000 147.9000 ;
	    RECT 75.0000 147.8000 75.4000 148.2000 ;
	    RECT 75.8000 147.8000 76.2000 148.6000 ;
	    RECT 76.7000 147.2000 77.0000 148.9000 ;
	    RECT 79.5000 148.2000 79.9000 149.9000 ;
	    RECT 79.0000 147.9000 79.9000 148.2000 ;
	    RECT 75.0000 147.1000 75.4000 147.2000 ;
	    RECT 76.6000 147.1000 77.0000 147.2000 ;
	    RECT 75.0000 146.8000 77.0000 147.1000 ;
	    RECT 78.2000 146.8000 78.6000 147.6000 ;
	    RECT 75.0000 146.1000 75.4000 146.2000 ;
	    RECT 72.6000 145.8000 73.4000 146.1000 ;
	    RECT 74.2000 145.8000 75.4000 146.1000 ;
	    RECT 73.0000 145.6000 73.4000 145.8000 ;
	    RECT 75.0000 145.1000 75.3000 145.8000 ;
	    RECT 76.7000 145.1000 77.0000 146.8000 ;
	    RECT 77.4000 145.4000 77.8000 146.2000 ;
	    RECT 79.0000 146.1000 79.4000 147.9000 ;
	    RECT 82.4000 147.1000 82.8000 149.9000 ;
	    RECT 83.8000 147.8000 84.2000 148.6000 ;
	    RECT 82.4000 146.9000 83.3000 147.1000 ;
	    RECT 82.5000 146.8000 83.3000 146.9000 ;
	    RECT 79.0000 145.8000 81.0000 146.1000 ;
	    RECT 81.4000 145.8000 82.2000 146.2000 ;
	    RECT 72.6000 144.8000 74.6000 145.1000 ;
	    RECT 72.6000 141.1000 73.0000 144.8000 ;
	    RECT 74.2000 141.1000 74.6000 144.8000 ;
	    RECT 75.0000 141.1000 75.4000 145.1000 ;
	    RECT 76.6000 144.7000 77.5000 145.1000 ;
	    RECT 77.1000 141.1000 77.5000 144.7000 ;
	    RECT 79.0000 141.1000 79.4000 145.8000 ;
	    RECT 79.8000 144.4000 80.2000 145.2000 ;
	    RECT 80.6000 144.8000 81.0000 145.8000 ;
	    RECT 83.0000 145.2000 83.3000 146.8000 ;
	    RECT 83.8000 146.1000 84.2000 146.2000 ;
	    RECT 84.6000 146.1000 85.0000 149.9000 ;
	    RECT 85.4000 146.8000 85.8000 147.6000 ;
	    RECT 83.8000 145.8000 85.0000 146.1000 ;
	    RECT 83.0000 144.8000 83.4000 145.2000 ;
	    RECT 82.2000 143.8000 82.6000 144.6000 ;
	    RECT 83.0000 143.5000 83.3000 144.8000 ;
	    RECT 81.5000 143.2000 83.3000 143.5000 ;
	    RECT 81.5000 143.1000 81.8000 143.2000 ;
	    RECT 81.4000 141.1000 81.8000 143.1000 ;
	    RECT 83.0000 143.1000 83.3000 143.2000 ;
	    RECT 83.0000 141.1000 83.4000 143.1000 ;
	    RECT 84.6000 141.1000 85.0000 145.8000 ;
	    RECT 86.2000 141.1000 86.6000 149.9000 ;
	    RECT 88.5000 147.9000 89.3000 149.9000 ;
	    RECT 87.8000 146.4000 88.2000 147.2000 ;
	    RECT 88.7000 146.2000 89.0000 147.9000 ;
	    RECT 89.4000 146.8000 89.8000 147.2000 ;
	    RECT 89.4000 146.6000 89.7000 146.8000 ;
	    RECT 89.3000 146.2000 89.7000 146.6000 ;
	    RECT 87.0000 146.1000 87.4000 146.2000 ;
	    RECT 87.0000 145.8000 87.8000 146.1000 ;
	    RECT 88.6000 145.8000 89.0000 146.2000 ;
	    RECT 87.4000 145.6000 87.8000 145.8000 ;
	    RECT 88.7000 145.7000 89.0000 145.8000 ;
	    RECT 88.7000 145.4000 89.7000 145.7000 ;
	    RECT 90.2000 145.4000 90.6000 146.2000 ;
	    RECT 89.4000 145.1000 89.7000 145.4000 ;
	    RECT 87.0000 144.8000 89.0000 145.1000 ;
	    RECT 87.0000 141.1000 87.4000 144.8000 ;
	    RECT 88.6000 141.4000 89.0000 144.8000 ;
	    RECT 89.4000 141.7000 89.8000 145.1000 ;
	    RECT 90.2000 141.4000 90.6000 145.1000 ;
	    RECT 88.6000 141.1000 90.6000 141.4000 ;
	    RECT 91.0000 141.1000 91.4000 149.9000 ;
	    RECT 91.8000 146.8000 92.2000 147.6000 ;
	    RECT 93.2000 147.1000 93.6000 149.9000 ;
	    RECT 97.1000 148.2000 97.5000 149.9000 ;
	    RECT 96.6000 147.9000 97.5000 148.2000 ;
	    RECT 99.0000 148.8000 99.4000 149.9000 ;
	    RECT 101.2000 149.1000 101.6000 149.9000 ;
	    RECT 101.2000 148.8000 102.5000 149.1000 ;
	    RECT 92.7000 146.9000 93.6000 147.1000 ;
	    RECT 92.7000 146.8000 93.5000 146.9000 ;
	    RECT 95.8000 146.8000 96.2000 147.6000 ;
	    RECT 96.6000 147.1000 97.0000 147.9000 ;
	    RECT 99.0000 147.2000 99.3000 148.8000 ;
	    RECT 99.8000 147.8000 100.2000 148.6000 ;
	    RECT 98.2000 147.1000 98.6000 147.2000 ;
	    RECT 96.6000 146.8000 98.6000 147.1000 ;
	    RECT 99.0000 146.8000 99.4000 147.2000 ;
	    RECT 101.2000 147.1000 101.6000 148.8000 ;
	    RECT 102.2000 148.2000 102.5000 148.8000 ;
	    RECT 102.2000 147.8000 102.6000 148.2000 ;
	    RECT 100.7000 146.9000 101.6000 147.1000 ;
	    RECT 100.7000 146.8000 101.5000 146.9000 ;
	    RECT 103.8000 146.8000 104.2000 147.6000 ;
	    RECT 92.7000 145.2000 93.0000 146.8000 ;
	    RECT 93.8000 145.8000 94.6000 146.2000 ;
	    RECT 92.6000 144.8000 93.0000 145.2000 ;
	    RECT 95.0000 144.8000 95.4000 145.6000 ;
	    RECT 92.7000 143.5000 93.0000 144.8000 ;
	    RECT 93.4000 143.8000 93.8000 144.6000 ;
	    RECT 92.7000 143.2000 94.5000 143.5000 ;
	    RECT 92.7000 143.1000 93.0000 143.2000 ;
	    RECT 92.6000 141.1000 93.0000 143.1000 ;
	    RECT 94.2000 141.1000 94.6000 143.2000 ;
	    RECT 96.6000 141.1000 97.0000 146.8000 ;
	    RECT 98.2000 145.4000 98.6000 146.2000 ;
	    RECT 97.4000 144.4000 97.8000 145.2000 ;
	    RECT 99.0000 145.1000 99.3000 146.8000 ;
	    RECT 100.7000 145.2000 101.0000 146.8000 ;
	    RECT 101.8000 145.8000 102.6000 146.2000 ;
	    RECT 104.6000 146.1000 105.0000 149.9000 ;
	    RECT 106.2000 147.9000 106.6000 149.9000 ;
	    RECT 107.0000 148.0000 107.4000 149.9000 ;
	    RECT 108.6000 148.0000 109.0000 149.9000 ;
	    RECT 107.0000 147.9000 109.0000 148.0000 ;
	    RECT 109.4000 147.9000 109.8000 149.9000 ;
	    RECT 110.2000 148.0000 110.6000 149.9000 ;
	    RECT 111.8000 148.0000 112.2000 149.9000 ;
	    RECT 110.2000 147.9000 112.2000 148.0000 ;
	    RECT 106.3000 147.2000 106.6000 147.9000 ;
	    RECT 107.1000 147.7000 108.9000 147.9000 ;
	    RECT 108.2000 147.2000 108.6000 147.4000 ;
	    RECT 109.5000 147.2000 109.8000 147.9000 ;
	    RECT 110.3000 147.7000 112.1000 147.9000 ;
	    RECT 111.4000 147.2000 111.8000 147.4000 ;
	    RECT 106.2000 146.8000 107.5000 147.2000 ;
	    RECT 108.2000 146.9000 109.0000 147.2000 ;
	    RECT 108.6000 146.8000 109.0000 146.9000 ;
	    RECT 109.4000 146.8000 110.7000 147.2000 ;
	    RECT 111.4000 146.9000 112.2000 147.2000 ;
	    RECT 114.8000 147.1000 115.2000 149.9000 ;
	    RECT 117.4000 148.0000 117.8000 149.9000 ;
	    RECT 119.0000 148.0000 119.4000 149.9000 ;
	    RECT 117.4000 147.9000 119.4000 148.0000 ;
	    RECT 119.8000 147.9000 120.2000 149.9000 ;
	    RECT 120.6000 147.9000 121.0000 149.9000 ;
	    RECT 121.4000 148.0000 121.8000 149.9000 ;
	    RECT 123.0000 148.0000 123.4000 149.9000 ;
	    RECT 121.4000 147.9000 123.4000 148.0000 ;
	    RECT 117.5000 147.7000 119.3000 147.9000 ;
	    RECT 117.8000 147.2000 118.2000 147.4000 ;
	    RECT 119.8000 147.2000 120.1000 147.9000 ;
	    RECT 120.7000 147.2000 121.0000 147.9000 ;
	    RECT 121.5000 147.7000 123.3000 147.9000 ;
	    RECT 122.6000 147.2000 123.0000 147.4000 ;
	    RECT 125.6000 147.2000 126.0000 149.9000 ;
	    RECT 127.1000 148.2000 127.5000 148.6000 ;
	    RECT 127.0000 147.8000 127.4000 148.2000 ;
	    RECT 127.8000 147.9000 128.2000 149.9000 ;
	    RECT 130.2000 147.9000 130.6000 149.9000 ;
	    RECT 131.0000 148.0000 131.4000 149.9000 ;
	    RECT 132.6000 148.0000 133.0000 149.9000 ;
	    RECT 135.8000 148.9000 136.2000 149.9000 ;
	    RECT 137.4000 149.2000 137.8000 149.9000 ;
	    RECT 131.0000 147.9000 133.0000 148.0000 ;
	    RECT 135.6000 148.8000 136.2000 148.9000 ;
	    RECT 137.3000 148.8000 137.8000 149.2000 ;
	    RECT 135.6000 148.5000 137.6000 148.8000 ;
	    RECT 111.8000 146.8000 112.2000 146.9000 ;
	    RECT 114.3000 146.9000 115.2000 147.1000 ;
	    RECT 117.4000 146.9000 118.2000 147.2000 ;
	    RECT 114.3000 146.8000 115.1000 146.9000 ;
	    RECT 117.4000 146.8000 117.8000 146.9000 ;
	    RECT 118.9000 146.8000 120.2000 147.2000 ;
	    RECT 120.6000 146.8000 121.9000 147.2000 ;
	    RECT 122.6000 146.9000 123.4000 147.2000 ;
	    RECT 123.0000 146.8000 123.4000 146.9000 ;
	    RECT 125.4000 147.1000 126.0000 147.2000 ;
	    RECT 125.4000 146.8000 126.5000 147.1000 ;
	    RECT 105.4000 146.1000 105.8000 146.2000 ;
	    RECT 104.6000 145.8000 105.8000 146.1000 ;
	    RECT 98.5000 144.7000 99.4000 145.1000 ;
	    RECT 100.6000 144.8000 101.0000 145.2000 ;
	    RECT 103.0000 144.8000 103.4000 145.6000 ;
	    RECT 98.5000 141.1000 98.9000 144.7000 ;
	    RECT 100.7000 143.5000 101.0000 144.8000 ;
	    RECT 101.4000 143.8000 101.8000 144.6000 ;
	    RECT 100.7000 143.2000 102.5000 143.5000 ;
	    RECT 100.7000 143.1000 101.0000 143.2000 ;
	    RECT 100.6000 141.1000 101.0000 143.1000 ;
	    RECT 102.2000 143.1000 102.5000 143.2000 ;
	    RECT 102.2000 141.1000 102.6000 143.1000 ;
	    RECT 104.6000 141.1000 105.0000 145.8000 ;
	    RECT 106.2000 145.1000 106.6000 145.2000 ;
	    RECT 107.2000 145.1000 107.5000 146.8000 ;
	    RECT 107.8000 145.8000 108.2000 146.6000 ;
	    RECT 109.4000 145.1000 109.8000 145.2000 ;
	    RECT 110.4000 145.1000 110.7000 146.8000 ;
	    RECT 111.0000 146.1000 111.4000 146.6000 ;
	    RECT 113.4000 146.1000 113.8000 146.2000 ;
	    RECT 111.0000 145.8000 113.8000 146.1000 ;
	    RECT 114.3000 145.2000 114.6000 146.8000 ;
	    RECT 115.4000 145.8000 116.2000 146.2000 ;
	    RECT 118.2000 145.8000 118.6000 146.6000 ;
	    RECT 106.2000 144.8000 106.9000 145.1000 ;
	    RECT 107.2000 144.8000 107.7000 145.1000 ;
	    RECT 109.4000 144.8000 110.1000 145.1000 ;
	    RECT 110.4000 144.8000 110.9000 145.1000 ;
	    RECT 114.2000 144.8000 114.6000 145.2000 ;
	    RECT 116.6000 144.8000 117.0000 145.6000 ;
	    RECT 118.9000 145.1000 119.2000 146.8000 ;
	    RECT 120.6000 146.2000 120.9000 146.8000 ;
	    RECT 120.6000 145.8000 121.0000 146.2000 ;
	    RECT 119.8000 145.1000 120.2000 145.2000 ;
	    RECT 118.7000 144.8000 119.2000 145.1000 ;
	    RECT 119.5000 144.8000 120.2000 145.1000 ;
	    RECT 120.6000 145.1000 121.0000 145.2000 ;
	    RECT 121.6000 145.1000 121.9000 146.8000 ;
	    RECT 122.2000 145.8000 122.6000 146.6000 ;
	    RECT 124.6000 145.8000 125.4000 146.2000 ;
	    RECT 120.6000 144.8000 121.3000 145.1000 ;
	    RECT 121.6000 144.8000 122.1000 145.1000 ;
	    RECT 123.8000 144.8000 124.2000 145.6000 ;
	    RECT 126.2000 145.2000 126.5000 146.8000 ;
	    RECT 127.0000 146.1000 127.4000 146.2000 ;
	    RECT 127.9000 146.1000 128.2000 147.9000 ;
	    RECT 130.3000 147.2000 130.6000 147.9000 ;
	    RECT 131.1000 147.7000 132.9000 147.9000 ;
	    RECT 132.2000 147.2000 132.6000 147.4000 ;
	    RECT 128.6000 147.1000 129.0000 147.2000 ;
	    RECT 129.4000 147.1000 129.8000 147.2000 ;
	    RECT 128.6000 146.8000 129.8000 147.1000 ;
	    RECT 130.2000 146.8000 131.5000 147.2000 ;
	    RECT 132.2000 146.9000 133.0000 147.2000 ;
	    RECT 132.6000 146.8000 133.0000 146.9000 ;
	    RECT 128.6000 146.4000 129.0000 146.8000 ;
	    RECT 129.4000 146.1000 129.8000 146.2000 ;
	    RECT 131.2000 146.1000 131.5000 146.8000 ;
	    RECT 127.0000 145.8000 128.2000 146.1000 ;
	    RECT 129.0000 145.8000 131.5000 146.1000 ;
	    RECT 131.8000 145.8000 132.2000 146.6000 ;
	    RECT 127.1000 145.2000 127.4000 145.8000 ;
	    RECT 129.0000 145.6000 129.4000 145.8000 ;
	    RECT 126.2000 144.8000 126.6000 145.2000 ;
	    RECT 106.6000 144.2000 106.9000 144.8000 ;
	    RECT 107.3000 144.2000 107.7000 144.8000 ;
	    RECT 109.8000 144.2000 110.1000 144.8000 ;
	    RECT 106.6000 143.8000 107.0000 144.2000 ;
	    RECT 107.3000 143.8000 108.2000 144.2000 ;
	    RECT 109.8000 143.8000 110.2000 144.2000 ;
	    RECT 107.3000 141.1000 107.7000 143.8000 ;
	    RECT 110.5000 141.1000 110.9000 144.8000 ;
	    RECT 114.3000 143.5000 114.6000 144.8000 ;
	    RECT 115.0000 143.8000 115.4000 144.6000 ;
	    RECT 114.3000 143.2000 116.1000 143.5000 ;
	    RECT 114.3000 143.1000 114.6000 143.2000 ;
	    RECT 114.2000 141.1000 114.6000 143.1000 ;
	    RECT 115.8000 141.1000 116.2000 143.2000 ;
	    RECT 118.7000 141.1000 119.1000 144.8000 ;
	    RECT 119.5000 144.2000 119.8000 144.8000 ;
	    RECT 119.4000 143.8000 119.8000 144.2000 ;
	    RECT 121.0000 144.2000 121.3000 144.8000 ;
	    RECT 121.0000 143.8000 121.4000 144.2000 ;
	    RECT 121.7000 141.1000 122.1000 144.8000 ;
	    RECT 125.4000 143.8000 125.8000 144.6000 ;
	    RECT 126.2000 143.5000 126.5000 144.8000 ;
	    RECT 124.7000 143.2000 126.5000 143.5000 ;
	    RECT 124.7000 143.1000 125.0000 143.2000 ;
	    RECT 124.6000 141.1000 125.0000 143.1000 ;
	    RECT 126.2000 143.1000 126.5000 143.2000 ;
	    RECT 126.2000 141.1000 126.6000 143.1000 ;
	    RECT 127.0000 141.1000 127.4000 145.2000 ;
	    RECT 130.2000 145.1000 130.6000 145.2000 ;
	    RECT 131.2000 145.1000 131.5000 145.8000 ;
	    RECT 135.6000 145.2000 135.9000 148.5000 ;
	    RECT 137.7000 147.8000 138.6000 148.2000 ;
	    RECT 139.8000 148.0000 140.2000 149.9000 ;
	    RECT 141.4000 148.0000 141.8000 149.9000 ;
	    RECT 139.8000 147.9000 141.8000 148.0000 ;
	    RECT 142.2000 147.9000 142.6000 149.9000 ;
	    RECT 144.3000 147.9000 145.1000 149.9000 ;
	    RECT 148.3000 147.9000 149.1000 149.9000 ;
	    RECT 151.8000 148.9000 152.2000 149.9000 ;
	    RECT 137.0000 146.8000 137.8000 147.2000 ;
	    RECT 138.2000 147.1000 138.5000 147.8000 ;
	    RECT 139.9000 147.7000 141.7000 147.9000 ;
	    RECT 140.2000 147.2000 140.6000 147.4000 ;
	    RECT 142.2000 147.2000 142.5000 147.9000 ;
	    RECT 139.8000 147.1000 140.6000 147.2000 ;
	    RECT 138.2000 146.9000 140.6000 147.1000 ;
	    RECT 141.3000 147.1000 142.6000 147.2000 ;
	    RECT 143.0000 147.1000 143.4000 147.2000 ;
	    RECT 138.2000 146.8000 140.2000 146.9000 ;
	    RECT 141.3000 146.8000 143.4000 147.1000 ;
	    RECT 143.8000 146.8000 144.2000 147.2000 ;
	    RECT 136.2000 145.8000 137.0000 146.2000 ;
	    RECT 137.4000 146.1000 137.7000 146.8000 ;
	    RECT 140.6000 146.1000 141.0000 146.6000 ;
	    RECT 137.4000 145.8000 141.0000 146.1000 ;
	    RECT 127.8000 144.8000 129.8000 145.1000 ;
	    RECT 130.2000 144.8000 130.9000 145.1000 ;
	    RECT 131.2000 144.8000 131.7000 145.1000 ;
	    RECT 134.2000 144.9000 135.9000 145.2000 ;
	    RECT 141.3000 145.1000 141.6000 146.8000 ;
	    RECT 143.9000 146.6000 144.2000 146.8000 ;
	    RECT 143.9000 146.2000 144.3000 146.6000 ;
	    RECT 144.6000 146.2000 144.9000 147.9000 ;
	    RECT 145.4000 147.1000 145.8000 147.2000 ;
	    RECT 147.8000 147.1000 148.2000 147.2000 ;
	    RECT 145.4000 146.8000 148.2000 147.1000 ;
	    RECT 145.4000 146.4000 145.8000 146.8000 ;
	    RECT 147.9000 146.6000 148.2000 146.8000 ;
	    RECT 147.9000 146.2000 148.3000 146.6000 ;
	    RECT 148.6000 146.2000 148.9000 147.9000 ;
	    RECT 151.0000 147.8000 151.4000 148.6000 ;
	    RECT 151.9000 147.2000 152.2000 148.9000 ;
	    RECT 149.4000 146.4000 149.8000 147.2000 ;
	    RECT 151.8000 146.8000 152.2000 147.2000 ;
	    RECT 155.2000 147.1000 155.6000 149.9000 ;
	    RECT 156.6000 148.0000 157.0000 149.9000 ;
	    RECT 158.2000 148.0000 158.6000 149.9000 ;
	    RECT 156.6000 147.9000 158.6000 148.0000 ;
	    RECT 159.0000 147.9000 159.4000 149.9000 ;
	    RECT 160.6000 148.8000 161.0000 149.9000 ;
	    RECT 156.7000 147.7000 158.5000 147.9000 ;
	    RECT 157.0000 147.2000 157.4000 147.4000 ;
	    RECT 159.0000 147.2000 159.3000 147.9000 ;
	    RECT 159.8000 147.8000 160.2000 148.6000 ;
	    RECT 160.7000 147.2000 161.0000 148.8000 ;
	    RECT 162.2000 147.5000 162.6000 149.9000 ;
	    RECT 164.4000 149.2000 164.8000 149.9000 ;
	    RECT 163.8000 148.9000 164.8000 149.2000 ;
	    RECT 166.6000 148.9000 167.0000 149.9000 ;
	    RECT 168.7000 149.2000 169.3000 149.9000 ;
	    RECT 168.6000 148.9000 169.3000 149.2000 ;
	    RECT 163.8000 148.5000 164.2000 148.9000 ;
	    RECT 166.6000 148.6000 166.9000 148.9000 ;
	    RECT 164.6000 148.2000 165.0000 148.6000 ;
	    RECT 165.5000 148.3000 166.9000 148.6000 ;
	    RECT 168.6000 148.5000 169.0000 148.9000 ;
	    RECT 165.5000 148.2000 165.9000 148.3000 ;
	    RECT 155.2000 146.9000 156.1000 147.1000 ;
	    RECT 155.3000 146.8000 156.1000 146.9000 ;
	    RECT 156.6000 146.9000 157.4000 147.2000 ;
	    RECT 156.6000 146.8000 157.0000 146.9000 ;
	    RECT 158.1000 146.8000 159.4000 147.2000 ;
	    RECT 160.6000 146.8000 161.0000 147.2000 ;
	    RECT 162.6000 147.1000 163.4000 147.2000 ;
	    RECT 164.7000 147.1000 165.0000 148.2000 ;
	    RECT 169.5000 147.7000 169.9000 147.8000 ;
	    RECT 171.0000 147.7000 171.4000 149.9000 ;
	    RECT 169.5000 147.4000 171.4000 147.7000 ;
	    RECT 165.4000 147.1000 165.8000 147.2000 ;
	    RECT 167.5000 147.1000 167.9000 147.2000 ;
	    RECT 162.6000 146.8000 168.1000 147.1000 ;
	    RECT 143.0000 145.4000 143.4000 146.2000 ;
	    RECT 144.6000 145.8000 145.0000 146.2000 ;
	    RECT 146.2000 146.1000 146.6000 146.2000 ;
	    RECT 147.0000 146.1000 147.4000 146.2000 ;
	    RECT 145.8000 145.8000 147.4000 146.1000 ;
	    RECT 144.6000 145.7000 144.9000 145.8000 ;
	    RECT 143.9000 145.4000 144.9000 145.7000 ;
	    RECT 145.8000 145.6000 146.2000 145.8000 ;
	    RECT 147.0000 145.4000 147.4000 145.8000 ;
	    RECT 148.6000 145.8000 149.0000 146.2000 ;
	    RECT 150.2000 146.1000 150.6000 146.2000 ;
	    RECT 149.8000 145.8000 150.6000 146.1000 ;
	    RECT 148.6000 145.7000 148.9000 145.8000 ;
	    RECT 147.9000 145.4000 148.9000 145.7000 ;
	    RECT 149.8000 145.6000 150.2000 145.8000 ;
	    RECT 142.2000 145.1000 142.6000 145.2000 ;
	    RECT 143.9000 145.1000 144.2000 145.4000 ;
	    RECT 147.9000 145.1000 148.2000 145.4000 ;
	    RECT 151.9000 145.1000 152.2000 146.8000 ;
	    RECT 152.6000 145.4000 153.0000 146.2000 ;
	    RECT 154.2000 145.8000 155.0000 146.2000 ;
	    RECT 134.2000 144.8000 134.6000 144.9000 ;
	    RECT 127.8000 141.1000 128.2000 144.8000 ;
	    RECT 129.4000 141.1000 129.8000 144.8000 ;
	    RECT 130.6000 144.2000 130.9000 144.8000 ;
	    RECT 130.6000 143.8000 131.0000 144.2000 ;
	    RECT 131.3000 141.1000 131.7000 144.8000 ;
	    RECT 134.3000 144.5000 134.6000 144.8000 ;
	    RECT 141.1000 144.8000 141.6000 145.1000 ;
	    RECT 141.9000 144.8000 142.6000 145.1000 ;
	    RECT 135.1000 144.5000 136.9000 144.6000 ;
	    RECT 133.4000 141.5000 133.8000 144.5000 ;
	    RECT 134.2000 141.7000 134.6000 144.5000 ;
	    RECT 135.0000 144.3000 136.9000 144.5000 ;
	    RECT 133.5000 141.4000 133.8000 141.5000 ;
	    RECT 135.0000 141.5000 135.4000 144.3000 ;
	    RECT 136.6000 144.1000 136.9000 144.3000 ;
	    RECT 137.5000 144.4000 139.3000 144.7000 ;
	    RECT 137.5000 144.1000 137.8000 144.4000 ;
	    RECT 135.0000 141.4000 135.3000 141.5000 ;
	    RECT 133.5000 141.1000 135.3000 141.4000 ;
	    RECT 135.8000 141.4000 136.2000 144.0000 ;
	    RECT 136.6000 141.7000 137.0000 144.1000 ;
	    RECT 137.4000 141.4000 137.8000 144.1000 ;
	    RECT 135.8000 141.1000 137.8000 141.4000 ;
	    RECT 139.0000 144.1000 139.3000 144.4000 ;
	    RECT 139.0000 141.1000 139.4000 144.1000 ;
	    RECT 141.1000 141.1000 141.5000 144.8000 ;
	    RECT 141.9000 144.2000 142.2000 144.8000 ;
	    RECT 141.8000 143.8000 142.2000 144.2000 ;
	    RECT 143.0000 141.4000 143.4000 145.1000 ;
	    RECT 143.8000 141.7000 144.2000 145.1000 ;
	    RECT 144.6000 144.8000 146.6000 145.1000 ;
	    RECT 144.6000 141.4000 145.0000 144.8000 ;
	    RECT 143.0000 141.1000 145.0000 141.4000 ;
	    RECT 146.2000 141.1000 146.6000 144.8000 ;
	    RECT 147.0000 141.4000 147.4000 145.1000 ;
	    RECT 147.8000 141.7000 148.2000 145.1000 ;
	    RECT 148.6000 144.8000 150.6000 145.1000 ;
	    RECT 148.6000 141.4000 149.0000 144.8000 ;
	    RECT 147.0000 141.1000 149.0000 141.4000 ;
	    RECT 150.2000 141.1000 150.6000 144.8000 ;
	    RECT 151.8000 144.7000 152.7000 145.1000 ;
	    RECT 152.3000 144.1000 152.7000 144.7000 ;
	    RECT 153.4000 144.8000 153.8000 145.6000 ;
	    RECT 155.8000 145.2000 156.1000 146.8000 ;
	    RECT 157.4000 145.8000 157.8000 146.6000 ;
	    RECT 155.8000 144.8000 156.2000 145.2000 ;
	    RECT 158.1000 145.1000 158.4000 146.8000 ;
	    RECT 159.0000 145.1000 159.4000 145.2000 ;
	    RECT 160.7000 145.1000 161.0000 146.8000 ;
	    RECT 164.1000 146.7000 164.5000 146.8000 ;
	    RECT 163.3000 146.2000 163.7000 146.3000 ;
	    RECT 161.4000 145.4000 161.8000 146.2000 ;
	    RECT 163.3000 145.9000 165.8000 146.2000 ;
	    RECT 165.4000 145.8000 165.8000 145.9000 ;
	    RECT 162.2000 145.5000 165.0000 145.6000 ;
	    RECT 162.2000 145.4000 165.1000 145.5000 ;
	    RECT 162.2000 145.3000 167.1000 145.4000 ;
	    RECT 157.9000 144.8000 158.4000 145.1000 ;
	    RECT 158.7000 144.8000 159.4000 145.1000 ;
	    RECT 153.4000 144.1000 153.7000 144.8000 ;
	    RECT 152.3000 143.8000 153.7000 144.1000 ;
	    RECT 155.0000 143.8000 155.4000 144.6000 ;
	    RECT 152.3000 141.1000 152.7000 143.8000 ;
	    RECT 155.8000 143.5000 156.1000 144.8000 ;
	    RECT 154.3000 143.2000 156.1000 143.5000 ;
	    RECT 154.3000 143.1000 154.6000 143.2000 ;
	    RECT 154.2000 141.1000 154.6000 143.1000 ;
	    RECT 155.8000 143.1000 156.1000 143.2000 ;
	    RECT 155.8000 141.1000 156.2000 143.1000 ;
	    RECT 157.9000 142.2000 158.3000 144.8000 ;
	    RECT 158.7000 144.2000 159.0000 144.8000 ;
	    RECT 160.6000 144.7000 161.5000 145.1000 ;
	    RECT 158.6000 143.8000 159.0000 144.2000 ;
	    RECT 157.4000 141.8000 158.3000 142.2000 ;
	    RECT 157.9000 141.1000 158.3000 141.8000 ;
	    RECT 161.1000 141.1000 161.5000 144.7000 ;
	    RECT 162.2000 141.1000 162.6000 145.3000 ;
	    RECT 164.7000 145.1000 167.1000 145.3000 ;
	    RECT 163.8000 144.5000 166.5000 144.8000 ;
	    RECT 163.8000 144.4000 164.2000 144.5000 ;
	    RECT 166.1000 144.4000 166.5000 144.5000 ;
	    RECT 166.8000 144.5000 167.1000 145.1000 ;
	    RECT 167.8000 145.2000 168.1000 146.8000 ;
	    RECT 168.6000 146.4000 169.0000 146.5000 ;
	    RECT 168.6000 146.1000 170.5000 146.4000 ;
	    RECT 170.1000 146.0000 170.5000 146.1000 ;
	    RECT 169.3000 145.7000 169.7000 145.8000 ;
	    RECT 171.0000 145.7000 171.4000 147.4000 ;
	    RECT 169.3000 145.4000 171.4000 145.7000 ;
	    RECT 167.8000 144.9000 169.0000 145.2000 ;
	    RECT 167.5000 144.5000 167.9000 144.6000 ;
	    RECT 166.8000 144.2000 167.9000 144.5000 ;
	    RECT 168.7000 144.4000 169.0000 144.9000 ;
	    RECT 168.7000 144.0000 169.4000 144.4000 ;
	    RECT 165.5000 143.7000 165.9000 143.8000 ;
	    RECT 166.9000 143.7000 167.3000 143.8000 ;
	    RECT 163.8000 143.1000 164.2000 143.5000 ;
	    RECT 165.5000 143.4000 167.3000 143.7000 ;
	    RECT 166.6000 143.1000 166.9000 143.4000 ;
	    RECT 168.6000 143.1000 169.0000 143.5000 ;
	    RECT 163.8000 142.8000 164.8000 143.1000 ;
	    RECT 164.4000 141.1000 164.8000 142.8000 ;
	    RECT 166.6000 141.1000 167.0000 143.1000 ;
	    RECT 168.7000 141.1000 169.3000 143.1000 ;
	    RECT 171.0000 141.1000 171.4000 145.4000 ;
	    RECT 0.6000 136.2000 1.0000 139.9000 ;
	    RECT 0.6000 135.9000 1.7000 136.2000 ;
	    RECT 2.2000 135.9000 2.6000 139.9000 ;
	    RECT 1.4000 135.6000 1.7000 135.9000 ;
	    RECT 1.4000 135.2000 2.0000 135.6000 ;
	    RECT 1.4000 133.7000 1.7000 135.2000 ;
	    RECT 2.3000 134.8000 2.6000 135.9000 ;
	    RECT 0.6000 133.4000 1.7000 133.7000 ;
	    RECT 0.6000 131.1000 1.0000 133.4000 ;
	    RECT 2.2000 131.1000 2.6000 134.8000 ;
	    RECT 3.8000 133.1000 4.2000 139.9000 ;
	    RECT 4.6000 135.8000 5.0000 136.6000 ;
	    RECT 5.4000 135.6000 5.8000 139.9000 ;
	    RECT 7.5000 136.2000 7.9000 139.9000 ;
	    RECT 9.4000 137.9000 9.8000 139.9000 ;
	    RECT 9.5000 137.8000 9.8000 137.9000 ;
	    RECT 11.0000 137.9000 11.4000 139.9000 ;
	    RECT 11.0000 137.8000 11.3000 137.9000 ;
	    RECT 9.5000 137.5000 11.3000 137.8000 ;
	    RECT 10.2000 136.4000 10.6000 137.2000 ;
	    RECT 11.0000 136.2000 11.3000 137.5000 ;
	    RECT 12.6000 137.1000 13.0000 139.9000 ;
	    RECT 11.8000 136.8000 13.0000 137.1000 ;
	    RECT 11.8000 136.2000 12.1000 136.8000 ;
	    RECT 7.5000 135.9000 8.2000 136.2000 ;
	    RECT 5.4000 135.4000 7.4000 135.6000 ;
	    RECT 5.4000 135.3000 7.5000 135.4000 ;
	    RECT 7.1000 135.0000 7.5000 135.3000 ;
	    RECT 7.9000 135.2000 8.2000 135.9000 ;
	    RECT 8.6000 135.4000 9.0000 136.2000 ;
	    RECT 11.0000 135.8000 11.4000 136.2000 ;
	    RECT 11.8000 135.8000 12.2000 136.2000 ;
	    RECT 7.2000 133.5000 7.5000 135.0000 ;
	    RECT 7.8000 134.8000 8.2000 135.2000 ;
	    RECT 9.4000 134.8000 10.2000 135.2000 ;
	    RECT 7.9000 134.2000 8.2000 134.8000 ;
	    RECT 11.0000 134.2000 11.3000 135.8000 ;
	    RECT 7.8000 133.8000 8.2000 134.2000 ;
	    RECT 10.5000 134.1000 11.3000 134.2000 ;
	    RECT 6.3000 133.2000 7.5000 133.5000 ;
	    RECT 3.8000 132.8000 4.7000 133.1000 ;
	    RECT 4.3000 132.2000 4.7000 132.8000 ;
	    RECT 5.4000 132.4000 5.8000 133.2000 ;
	    RECT 3.8000 131.8000 4.7000 132.2000 ;
	    RECT 6.3000 132.1000 6.6000 133.2000 ;
	    RECT 7.9000 133.1000 8.2000 133.8000 ;
	    RECT 4.3000 131.1000 4.7000 131.8000 ;
	    RECT 6.2000 131.1000 6.6000 132.1000 ;
	    RECT 7.8000 131.1000 8.2000 133.1000 ;
	    RECT 10.4000 133.9000 11.3000 134.1000 ;
	    RECT 9.4000 132.1000 9.8000 132.2000 ;
	    RECT 10.4000 132.1000 10.8000 133.9000 ;
	    RECT 11.8000 133.4000 12.2000 134.2000 ;
	    RECT 12.6000 133.1000 13.0000 136.8000 ;
	    RECT 13.4000 135.8000 13.8000 136.6000 ;
	    RECT 14.2000 135.8000 14.6000 136.6000 ;
	    RECT 15.0000 133.1000 15.4000 139.9000 ;
	    RECT 16.6000 135.8000 17.0000 136.6000 ;
	    RECT 17.4000 133.1000 17.8000 139.9000 ;
	    RECT 19.0000 135.8000 19.4000 136.6000 ;
	    RECT 18.2000 133.4000 18.6000 134.2000 ;
	    RECT 19.8000 133.1000 20.2000 139.9000 ;
	    RECT 12.6000 132.8000 13.5000 133.1000 ;
	    RECT 9.4000 131.8000 10.8000 132.1000 ;
	    RECT 10.4000 131.1000 10.8000 131.8000 ;
	    RECT 13.1000 131.1000 13.5000 132.8000 ;
	    RECT 14.5000 132.8000 15.4000 133.1000 ;
	    RECT 16.9000 132.8000 17.8000 133.1000 ;
	    RECT 19.3000 132.8000 20.2000 133.1000 ;
	    RECT 22.2000 133.1000 22.6000 139.9000 ;
	    RECT 23.0000 135.8000 23.4000 136.6000 ;
	    RECT 23.8000 136.2000 24.2000 139.9000 ;
	    RECT 23.8000 135.9000 24.9000 136.2000 ;
	    RECT 25.4000 135.9000 25.8000 139.9000 ;
	    RECT 24.6000 135.6000 24.9000 135.9000 ;
	    RECT 24.6000 135.2000 25.2000 135.6000 ;
	    RECT 24.6000 133.7000 24.9000 135.2000 ;
	    RECT 25.5000 134.8000 25.8000 135.9000 ;
	    RECT 23.8000 133.4000 24.9000 133.7000 ;
	    RECT 22.2000 132.8000 23.1000 133.1000 ;
	    RECT 14.5000 132.2000 14.9000 132.8000 ;
	    RECT 16.9000 132.2000 17.3000 132.8000 ;
	    RECT 19.3000 132.2000 19.7000 132.8000 ;
	    RECT 22.7000 132.2000 23.1000 132.8000 ;
	    RECT 14.2000 131.8000 14.9000 132.2000 ;
	    RECT 16.6000 131.8000 17.3000 132.2000 ;
	    RECT 19.0000 131.8000 19.7000 132.2000 ;
	    RECT 22.2000 131.8000 23.1000 132.2000 ;
	    RECT 14.5000 131.1000 14.9000 131.8000 ;
	    RECT 16.9000 131.1000 17.3000 131.8000 ;
	    RECT 19.3000 131.1000 19.7000 131.8000 ;
	    RECT 22.7000 131.1000 23.1000 131.8000 ;
	    RECT 23.8000 131.1000 24.2000 133.4000 ;
	    RECT 25.4000 131.1000 25.8000 134.8000 ;
	    RECT 26.2000 131.1000 26.6000 139.9000 ;
	    RECT 27.8000 135.8000 28.2000 136.6000 ;
	    RECT 28.6000 133.1000 29.0000 139.9000 ;
	    RECT 29.4000 133.4000 29.8000 134.2000 ;
	    RECT 28.1000 132.8000 29.0000 133.1000 ;
	    RECT 31.0000 133.1000 31.4000 139.9000 ;
	    RECT 31.8000 135.8000 32.2000 136.6000 ;
	    RECT 32.6000 135.6000 33.0000 139.9000 ;
	    RECT 34.7000 136.2000 35.1000 139.9000 ;
	    RECT 34.7000 135.9000 35.4000 136.2000 ;
	    RECT 32.6000 135.4000 34.6000 135.6000 ;
	    RECT 32.6000 135.3000 34.7000 135.4000 ;
	    RECT 34.3000 135.0000 34.7000 135.3000 ;
	    RECT 35.1000 135.2000 35.4000 135.9000 ;
	    RECT 34.4000 133.5000 34.7000 135.0000 ;
	    RECT 35.0000 134.8000 35.4000 135.2000 ;
	    RECT 33.5000 133.2000 34.7000 133.5000 ;
	    RECT 31.0000 132.8000 31.9000 133.1000 ;
	    RECT 28.1000 132.2000 28.5000 132.8000 ;
	    RECT 31.5000 132.2000 31.9000 132.8000 ;
	    RECT 32.6000 132.4000 33.0000 133.2000 ;
	    RECT 28.1000 131.8000 29.0000 132.2000 ;
	    RECT 31.5000 131.8000 32.2000 132.2000 ;
	    RECT 33.5000 132.1000 33.8000 133.2000 ;
	    RECT 35.1000 133.1000 35.4000 134.8000 ;
	    RECT 28.1000 131.1000 28.5000 131.8000 ;
	    RECT 31.5000 131.1000 31.9000 131.8000 ;
	    RECT 33.4000 131.1000 33.8000 132.1000 ;
	    RECT 35.0000 131.1000 35.4000 133.1000 ;
	    RECT 36.6000 133.1000 37.0000 139.9000 ;
	    RECT 37.4000 135.8000 37.8000 136.6000 ;
	    RECT 39.0000 134.1000 39.4000 139.9000 ;
	    RECT 41.1000 136.2000 41.5000 139.9000 ;
	    RECT 41.8000 136.8000 42.2000 137.2000 ;
	    RECT 41.9000 136.2000 42.2000 136.8000 ;
	    RECT 40.6000 135.8000 41.6000 136.2000 ;
	    RECT 41.9000 136.1000 42.6000 136.2000 ;
	    RECT 43.8000 136.1000 44.2000 139.9000 ;
	    RECT 41.9000 135.9000 44.2000 136.1000 ;
	    RECT 42.2000 135.8000 44.2000 135.9000 ;
	    RECT 40.6000 134.4000 41.0000 135.2000 ;
	    RECT 41.3000 134.2000 41.6000 135.8000 ;
	    RECT 39.8000 134.1000 40.2000 134.2000 ;
	    RECT 39.0000 133.8000 40.6000 134.1000 ;
	    RECT 41.3000 133.8000 42.6000 134.2000 ;
	    RECT 36.6000 132.8000 37.5000 133.1000 ;
	    RECT 37.1000 132.2000 37.5000 132.8000 ;
	    RECT 36.6000 131.8000 37.5000 132.2000 ;
	    RECT 37.1000 131.1000 37.5000 131.8000 ;
	    RECT 39.0000 131.1000 39.4000 133.8000 ;
	    RECT 40.2000 133.6000 40.6000 133.8000 ;
	    RECT 39.9000 133.1000 41.7000 133.3000 ;
	    RECT 42.2000 133.1000 42.5000 133.8000 ;
	    RECT 43.0000 133.4000 43.4000 134.2000 ;
	    RECT 43.8000 133.1000 44.2000 135.8000 ;
	    RECT 46.2000 134.1000 46.6000 139.9000 ;
	    RECT 48.3000 136.2000 48.7000 139.9000 ;
	    RECT 49.0000 136.8000 49.4000 137.2000 ;
	    RECT 49.1000 136.2000 49.4000 136.8000 ;
	    RECT 48.3000 135.9000 48.8000 136.2000 ;
	    RECT 49.1000 135.9000 49.8000 136.2000 ;
	    RECT 47.8000 134.4000 48.2000 135.2000 ;
	    RECT 48.5000 134.2000 48.8000 135.9000 ;
	    RECT 49.4000 135.8000 49.8000 135.9000 ;
	    RECT 49.4000 135.1000 49.7000 135.8000 ;
	    RECT 51.0000 135.1000 51.4000 139.9000 ;
	    RECT 51.8000 136.1000 52.2000 136.2000 ;
	    RECT 52.6000 136.1000 53.0000 136.6000 ;
	    RECT 51.8000 135.8000 53.0000 136.1000 ;
	    RECT 49.4000 134.8000 51.4000 135.1000 ;
	    RECT 47.0000 134.1000 47.4000 134.2000 ;
	    RECT 46.2000 133.8000 47.8000 134.1000 ;
	    RECT 48.5000 133.8000 49.8000 134.2000 ;
	    RECT 39.8000 133.0000 41.8000 133.1000 ;
	    RECT 39.8000 131.1000 40.2000 133.0000 ;
	    RECT 41.4000 131.1000 41.8000 133.0000 ;
	    RECT 42.2000 131.1000 42.6000 133.1000 ;
	    RECT 43.8000 132.8000 44.7000 133.1000 ;
	    RECT 44.3000 131.1000 44.7000 132.8000 ;
	    RECT 46.2000 131.1000 46.6000 133.8000 ;
	    RECT 47.4000 133.6000 47.8000 133.8000 ;
	    RECT 47.1000 133.1000 48.9000 133.3000 ;
	    RECT 49.4000 133.1000 49.7000 133.8000 ;
	    RECT 51.0000 133.1000 51.4000 134.8000 ;
	    RECT 51.8000 133.4000 52.2000 134.2000 ;
	    RECT 53.4000 133.1000 53.8000 139.9000 ;
	    RECT 56.1000 137.2000 56.5000 139.9000 ;
	    RECT 55.4000 136.8000 55.8000 137.2000 ;
	    RECT 56.1000 136.8000 57.0000 137.2000 ;
	    RECT 55.4000 136.2000 55.7000 136.8000 ;
	    RECT 56.1000 136.2000 56.5000 136.8000 ;
	    RECT 55.0000 135.9000 55.7000 136.2000 ;
	    RECT 56.0000 135.9000 56.5000 136.2000 ;
	    RECT 55.0000 135.8000 55.4000 135.9000 ;
	    RECT 56.0000 134.2000 56.3000 135.9000 ;
	    RECT 58.2000 135.8000 58.6000 136.6000 ;
	    RECT 56.6000 134.4000 57.0000 135.2000 ;
	    RECT 54.2000 133.4000 54.6000 134.2000 ;
	    RECT 55.0000 133.8000 56.3000 134.2000 ;
	    RECT 57.4000 134.1000 57.8000 134.2000 ;
	    RECT 57.0000 133.8000 57.8000 134.1000 ;
	    RECT 55.1000 133.1000 55.4000 133.8000 ;
	    RECT 57.0000 133.6000 57.4000 133.8000 ;
	    RECT 55.9000 133.1000 57.7000 133.3000 ;
	    RECT 59.0000 133.1000 59.4000 139.9000 ;
	    RECT 62.2000 135.8000 62.6000 136.6000 ;
	    RECT 63.0000 133.1000 63.4000 139.9000 ;
	    RECT 64.6000 135.6000 65.0000 139.9000 ;
	    RECT 66.7000 136.2000 67.1000 139.9000 ;
	    RECT 66.7000 135.9000 67.4000 136.2000 ;
	    RECT 64.6000 135.4000 66.6000 135.6000 ;
	    RECT 64.6000 135.3000 66.7000 135.4000 ;
	    RECT 66.3000 135.0000 66.7000 135.3000 ;
	    RECT 67.1000 135.2000 67.4000 135.9000 ;
	    RECT 67.8000 135.8000 68.2000 136.6000 ;
	    RECT 66.4000 133.5000 66.7000 135.0000 ;
	    RECT 67.0000 134.8000 67.4000 135.2000 ;
	    RECT 67.1000 134.1000 67.4000 134.8000 ;
	    RECT 67.8000 134.1000 68.2000 134.2000 ;
	    RECT 67.0000 133.8000 68.2000 134.1000 ;
	    RECT 65.5000 133.2000 66.7000 133.5000 ;
	    RECT 47.0000 133.0000 49.0000 133.1000 ;
	    RECT 47.0000 131.1000 47.4000 133.0000 ;
	    RECT 48.6000 131.1000 49.0000 133.0000 ;
	    RECT 49.4000 131.1000 49.8000 133.1000 ;
	    RECT 50.5000 132.8000 51.4000 133.1000 ;
	    RECT 52.9000 132.8000 53.8000 133.1000 ;
	    RECT 50.5000 131.1000 50.9000 132.8000 ;
	    RECT 52.9000 132.2000 53.3000 132.8000 ;
	    RECT 52.9000 131.8000 53.8000 132.2000 ;
	    RECT 52.9000 131.1000 53.3000 131.8000 ;
	    RECT 55.0000 131.1000 55.4000 133.1000 ;
	    RECT 55.8000 133.0000 57.8000 133.1000 ;
	    RECT 55.8000 131.1000 56.2000 133.0000 ;
	    RECT 57.4000 131.1000 57.8000 133.0000 ;
	    RECT 58.5000 132.8000 59.4000 133.1000 ;
	    RECT 62.5000 132.8000 63.4000 133.1000 ;
	    RECT 58.5000 132.2000 58.9000 132.8000 ;
	    RECT 62.5000 132.2000 62.9000 132.8000 ;
	    RECT 64.6000 132.4000 65.0000 133.2000 ;
	    RECT 58.5000 131.8000 59.4000 132.2000 ;
	    RECT 62.5000 131.8000 63.4000 132.2000 ;
	    RECT 65.5000 132.1000 65.8000 133.2000 ;
	    RECT 67.1000 133.1000 67.4000 133.8000 ;
	    RECT 68.6000 133.1000 69.0000 139.9000 ;
	    RECT 70.2000 133.4000 70.6000 134.2000 ;
	    RECT 58.5000 131.1000 58.9000 131.8000 ;
	    RECT 62.5000 131.1000 62.9000 131.8000 ;
	    RECT 65.4000 131.1000 65.8000 132.1000 ;
	    RECT 67.0000 131.1000 67.4000 133.1000 ;
	    RECT 68.1000 132.8000 69.0000 133.1000 ;
	    RECT 71.0000 133.1000 71.4000 139.9000 ;
	    RECT 71.8000 135.8000 72.2000 136.6000 ;
	    RECT 72.6000 135.6000 73.0000 139.9000 ;
	    RECT 74.7000 136.2000 75.1000 139.9000 ;
	    RECT 75.8000 137.9000 76.2000 139.9000 ;
	    RECT 75.9000 137.8000 76.2000 137.9000 ;
	    RECT 77.4000 137.9000 77.8000 139.9000 ;
	    RECT 77.4000 137.8000 77.7000 137.9000 ;
	    RECT 75.9000 137.5000 77.7000 137.8000 ;
	    RECT 75.9000 136.2000 76.2000 137.5000 ;
	    RECT 76.6000 136.4000 77.0000 137.2000 ;
	    RECT 74.7000 135.9000 75.4000 136.2000 ;
	    RECT 72.6000 135.4000 74.6000 135.6000 ;
	    RECT 72.6000 135.3000 74.7000 135.4000 ;
	    RECT 74.3000 135.0000 74.7000 135.3000 ;
	    RECT 75.1000 135.2000 75.4000 135.9000 ;
	    RECT 75.8000 135.8000 76.2000 136.2000 ;
	    RECT 74.4000 133.5000 74.7000 135.0000 ;
	    RECT 75.0000 134.8000 75.4000 135.2000 ;
	    RECT 75.1000 134.2000 75.4000 134.8000 ;
	    RECT 75.0000 133.8000 75.4000 134.2000 ;
	    RECT 75.9000 134.2000 76.2000 135.8000 ;
	    RECT 78.2000 135.4000 78.6000 136.2000 ;
	    RECT 79.0000 135.8000 79.4000 136.6000 ;
	    RECT 77.0000 134.8000 77.8000 135.2000 ;
	    RECT 75.9000 134.1000 76.7000 134.2000 ;
	    RECT 75.9000 133.9000 76.8000 134.1000 ;
	    RECT 73.5000 133.2000 74.7000 133.5000 ;
	    RECT 71.0000 132.8000 71.9000 133.1000 ;
	    RECT 68.1000 132.2000 68.5000 132.8000 ;
	    RECT 71.5000 132.2000 71.9000 132.8000 ;
	    RECT 72.6000 132.4000 73.0000 133.2000 ;
	    RECT 68.1000 131.8000 69.0000 132.2000 ;
	    RECT 71.5000 131.8000 72.2000 132.2000 ;
	    RECT 73.5000 132.1000 73.8000 133.2000 ;
	    RECT 75.1000 133.1000 75.4000 133.8000 ;
	    RECT 68.1000 131.1000 68.5000 131.8000 ;
	    RECT 71.5000 131.1000 71.9000 131.8000 ;
	    RECT 73.4000 131.1000 73.8000 132.1000 ;
	    RECT 75.0000 131.1000 75.4000 133.1000 ;
	    RECT 76.4000 132.1000 76.8000 133.9000 ;
	    RECT 79.8000 133.1000 80.2000 139.9000 ;
	    RECT 81.8000 136.8000 82.2000 137.2000 ;
	    RECT 81.8000 136.2000 82.1000 136.8000 ;
	    RECT 82.5000 136.2000 82.9000 139.9000 ;
	    RECT 85.9000 136.3000 86.3000 139.9000 ;
	    RECT 81.4000 135.9000 82.1000 136.2000 ;
	    RECT 82.4000 135.9000 82.9000 136.2000 ;
	    RECT 85.4000 135.9000 86.3000 136.3000 ;
	    RECT 88.3000 136.2000 88.7000 139.9000 ;
	    RECT 89.0000 136.8000 89.4000 137.2000 ;
	    RECT 89.1000 136.2000 89.4000 136.8000 ;
	    RECT 88.3000 135.9000 88.8000 136.2000 ;
	    RECT 89.1000 135.9000 89.8000 136.2000 ;
	    RECT 81.4000 135.8000 81.8000 135.9000 ;
	    RECT 82.4000 134.2000 82.7000 135.9000 ;
	    RECT 83.0000 134.4000 83.4000 135.2000 ;
	    RECT 85.5000 134.2000 85.8000 135.9000 ;
	    RECT 86.2000 134.8000 86.6000 135.6000 ;
	    RECT 87.8000 134.4000 88.2000 135.2000 ;
	    RECT 88.5000 135.1000 88.8000 135.9000 ;
	    RECT 89.4000 135.8000 89.8000 135.9000 ;
	    RECT 89.4000 135.1000 89.8000 135.2000 ;
	    RECT 88.5000 134.8000 89.8000 135.1000 ;
	    RECT 90.2000 134.8000 90.6000 135.2000 ;
	    RECT 88.5000 134.2000 88.8000 134.8000 ;
	    RECT 90.2000 134.2000 90.5000 134.8000 ;
	    RECT 81.4000 133.8000 82.7000 134.2000 ;
	    RECT 83.8000 134.1000 84.2000 134.2000 ;
	    RECT 83.4000 133.8000 84.2000 134.1000 ;
	    RECT 85.4000 134.1000 85.8000 134.2000 ;
	    RECT 87.0000 134.1000 87.4000 134.2000 ;
	    RECT 85.4000 133.8000 87.8000 134.1000 ;
	    RECT 88.5000 133.8000 89.8000 134.2000 ;
	    RECT 81.5000 133.1000 81.8000 133.8000 ;
	    RECT 83.4000 133.6000 83.8000 133.8000 ;
	    RECT 82.3000 133.1000 84.1000 133.3000 ;
	    RECT 79.3000 132.8000 80.2000 133.1000 ;
	    RECT 79.3000 132.2000 79.7000 132.8000 ;
	    RECT 77.4000 132.1000 77.8000 132.2000 ;
	    RECT 76.4000 131.8000 77.8000 132.1000 ;
	    RECT 79.0000 131.8000 79.7000 132.2000 ;
	    RECT 76.4000 131.1000 76.8000 131.8000 ;
	    RECT 79.3000 131.1000 79.7000 131.8000 ;
	    RECT 81.4000 131.1000 81.8000 133.1000 ;
	    RECT 82.2000 133.0000 84.2000 133.1000 ;
	    RECT 82.2000 131.1000 82.6000 133.0000 ;
	    RECT 83.8000 131.1000 84.2000 133.0000 ;
	    RECT 84.6000 132.4000 85.0000 133.2000 ;
	    RECT 85.5000 132.1000 85.8000 133.8000 ;
	    RECT 87.4000 133.6000 87.8000 133.8000 ;
	    RECT 87.1000 133.1000 88.9000 133.3000 ;
	    RECT 89.4000 133.1000 89.7000 133.8000 ;
	    RECT 90.2000 133.4000 90.6000 134.2000 ;
	    RECT 85.4000 131.1000 85.8000 132.1000 ;
	    RECT 87.0000 133.0000 89.0000 133.1000 ;
	    RECT 87.0000 131.1000 87.4000 133.0000 ;
	    RECT 88.6000 131.1000 89.0000 133.0000 ;
	    RECT 89.4000 131.1000 89.8000 133.1000 ;
	    RECT 91.0000 131.1000 91.4000 139.9000 ;
	    RECT 92.6000 137.9000 93.0000 139.9000 ;
	    RECT 92.7000 137.8000 93.0000 137.9000 ;
	    RECT 94.2000 137.9000 94.6000 139.9000 ;
	    RECT 95.8000 137.9000 96.2000 139.9000 ;
	    RECT 94.2000 137.8000 94.5000 137.9000 ;
	    RECT 92.7000 137.5000 94.5000 137.8000 ;
	    RECT 95.9000 137.8000 96.2000 137.9000 ;
	    RECT 97.4000 137.9000 97.8000 139.9000 ;
	    RECT 98.2000 137.9000 98.6000 139.9000 ;
	    RECT 97.4000 137.8000 97.7000 137.9000 ;
	    RECT 95.9000 137.5000 97.7000 137.8000 ;
	    RECT 93.4000 136.4000 93.8000 137.2000 ;
	    RECT 94.2000 136.2000 94.5000 137.5000 ;
	    RECT 96.6000 136.4000 97.0000 137.2000 ;
	    RECT 97.4000 136.2000 97.7000 137.5000 ;
	    RECT 98.3000 137.8000 98.6000 137.9000 ;
	    RECT 99.8000 137.9000 100.2000 139.9000 ;
	    RECT 101.4000 137.9000 101.8000 139.9000 ;
	    RECT 99.8000 137.8000 100.1000 137.9000 ;
	    RECT 98.3000 137.5000 100.1000 137.8000 ;
	    RECT 101.5000 137.8000 101.8000 137.9000 ;
	    RECT 103.0000 137.9000 103.4000 139.9000 ;
	    RECT 103.0000 137.8000 103.3000 137.9000 ;
	    RECT 101.5000 137.5000 103.3000 137.8000 ;
	    RECT 98.3000 136.2000 98.6000 137.5000 ;
	    RECT 99.0000 136.4000 99.4000 137.2000 ;
	    RECT 101.5000 136.2000 101.8000 137.5000 ;
	    RECT 102.2000 136.4000 102.6000 137.2000 ;
	    RECT 91.8000 135.4000 92.2000 136.2000 ;
	    RECT 94.2000 135.8000 94.6000 136.2000 ;
	    RECT 94.2000 135.2000 94.5000 135.8000 ;
	    RECT 95.0000 135.4000 95.4000 136.2000 ;
	    RECT 97.4000 135.8000 97.8000 136.2000 ;
	    RECT 98.2000 135.8000 98.6000 136.2000 ;
	    RECT 97.4000 135.2000 97.7000 135.8000 ;
	    RECT 92.6000 134.8000 93.4000 135.2000 ;
	    RECT 94.2000 134.8000 94.6000 135.2000 ;
	    RECT 95.8000 134.8000 96.6000 135.2000 ;
	    RECT 97.4000 134.8000 97.8000 135.2000 ;
	    RECT 94.2000 134.2000 94.5000 134.8000 ;
	    RECT 97.4000 134.2000 97.7000 134.8000 ;
	    RECT 93.7000 134.1000 94.5000 134.2000 ;
	    RECT 96.9000 134.1000 97.7000 134.2000 ;
	    RECT 93.6000 133.9000 94.5000 134.1000 ;
	    RECT 96.8000 133.9000 97.7000 134.1000 ;
	    RECT 98.3000 134.2000 98.6000 135.8000 ;
	    RECT 100.6000 135.4000 101.0000 136.2000 ;
	    RECT 101.4000 135.8000 101.8000 136.2000 ;
	    RECT 99.4000 134.8000 100.2000 135.2000 ;
	    RECT 101.5000 134.2000 101.8000 135.8000 ;
	    RECT 103.8000 135.4000 104.2000 136.2000 ;
	    RECT 102.2000 134.8000 103.4000 135.2000 ;
	    RECT 105.4000 135.1000 105.8000 139.9000 ;
	    RECT 106.5000 139.2000 106.9000 139.9000 ;
	    RECT 106.2000 138.8000 106.9000 139.2000 ;
	    RECT 106.5000 136.3000 106.9000 138.8000 ;
	    RECT 106.5000 135.9000 107.4000 136.3000 ;
	    RECT 108.6000 136.2000 109.0000 139.9000 ;
	    RECT 110.2000 136.2000 110.6000 139.9000 ;
	    RECT 108.6000 135.9000 110.6000 136.2000 ;
	    RECT 111.0000 139.1000 111.4000 139.9000 ;
	    RECT 112.6000 139.1000 113.0000 139.2000 ;
	    RECT 111.0000 138.8000 113.0000 139.1000 ;
	    RECT 111.0000 135.9000 111.4000 138.8000 ;
	    RECT 113.4000 135.9000 113.8000 139.9000 ;
	    RECT 114.2000 136.2000 114.6000 139.9000 ;
	    RECT 115.8000 136.2000 116.2000 139.9000 ;
	    RECT 117.9000 136.3000 118.3000 139.9000 ;
	    RECT 114.2000 135.9000 116.2000 136.2000 ;
	    RECT 117.4000 135.9000 118.3000 136.3000 ;
	    RECT 106.2000 135.1000 106.6000 135.6000 ;
	    RECT 105.4000 134.8000 106.6000 135.1000 ;
	    RECT 98.3000 134.1000 99.1000 134.2000 ;
	    RECT 101.5000 134.1000 102.3000 134.2000 ;
	    RECT 98.3000 133.9000 99.2000 134.1000 ;
	    RECT 101.5000 133.9000 102.4000 134.1000 ;
	    RECT 93.6000 131.1000 94.0000 133.9000 ;
	    RECT 96.8000 131.1000 97.2000 133.9000 ;
	    RECT 98.8000 131.1000 99.2000 133.9000 ;
	    RECT 102.0000 131.1000 102.4000 133.9000 ;
	    RECT 104.6000 132.4000 105.0000 133.2000 ;
	    RECT 105.4000 131.1000 105.8000 134.8000 ;
	    RECT 107.0000 134.2000 107.3000 135.9000 ;
	    RECT 109.0000 135.2000 109.4000 135.4000 ;
	    RECT 111.0000 135.2000 111.3000 135.9000 ;
	    RECT 113.5000 135.2000 113.8000 135.9000 ;
	    RECT 115.4000 135.2000 115.8000 135.4000 ;
	    RECT 108.6000 134.9000 109.4000 135.2000 ;
	    RECT 110.2000 134.9000 111.4000 135.2000 ;
	    RECT 108.6000 134.8000 109.0000 134.9000 ;
	    RECT 107.0000 133.8000 107.4000 134.2000 ;
	    RECT 107.8000 133.8000 108.2000 134.2000 ;
	    RECT 109.4000 133.8000 109.8000 134.6000 ;
	    RECT 107.0000 132.1000 107.3000 133.8000 ;
	    RECT 107.8000 133.2000 108.1000 133.8000 ;
	    RECT 107.8000 132.4000 108.2000 133.2000 ;
	    RECT 110.2000 133.1000 110.5000 134.9000 ;
	    RECT 111.0000 134.8000 111.4000 134.9000 ;
	    RECT 113.4000 134.9000 114.6000 135.2000 ;
	    RECT 115.4000 134.9000 116.2000 135.2000 ;
	    RECT 113.4000 134.8000 113.8000 134.9000 ;
	    RECT 111.0000 133.1000 111.4000 133.2000 ;
	    RECT 113.4000 133.1000 113.8000 133.2000 ;
	    RECT 114.3000 133.1000 114.6000 134.9000 ;
	    RECT 115.8000 134.8000 116.2000 134.9000 ;
	    RECT 115.0000 133.8000 115.4000 134.6000 ;
	    RECT 117.5000 134.2000 117.8000 135.9000 ;
	    RECT 118.2000 135.1000 118.6000 135.6000 ;
	    RECT 119.0000 135.1000 119.4000 139.9000 ;
	    RECT 118.2000 134.8000 119.4000 135.1000 ;
	    RECT 117.4000 133.8000 117.8000 134.2000 ;
	    RECT 107.0000 131.1000 107.4000 132.1000 ;
	    RECT 110.2000 131.1000 110.6000 133.1000 ;
	    RECT 111.0000 132.8000 113.8000 133.1000 ;
	    RECT 110.9000 132.4000 111.3000 132.8000 ;
	    RECT 113.5000 132.4000 113.9000 132.8000 ;
	    RECT 114.2000 131.1000 114.6000 133.1000 ;
	    RECT 116.6000 132.4000 117.0000 133.2000 ;
	    RECT 117.5000 133.1000 117.8000 133.8000 ;
	    RECT 118.2000 133.8000 118.6000 134.2000 ;
	    RECT 118.2000 133.1000 118.5000 133.8000 ;
	    RECT 117.4000 132.8000 118.5000 133.1000 ;
	    RECT 117.5000 132.1000 117.8000 132.8000 ;
	    RECT 117.4000 131.1000 117.8000 132.1000 ;
	    RECT 119.0000 131.1000 119.4000 134.8000 ;
	    RECT 120.6000 134.1000 121.0000 139.9000 ;
	    RECT 123.0000 135.1000 123.4000 139.9000 ;
	    RECT 125.4000 137.9000 125.8000 139.9000 ;
	    RECT 125.5000 137.8000 125.8000 137.9000 ;
	    RECT 127.0000 137.9000 127.4000 139.9000 ;
	    RECT 129.1000 139.2000 129.5000 139.9000 ;
	    RECT 128.6000 138.8000 129.5000 139.2000 ;
	    RECT 127.0000 137.8000 127.3000 137.9000 ;
	    RECT 125.5000 137.5000 127.3000 137.8000 ;
	    RECT 123.8000 135.8000 124.2000 136.6000 ;
	    RECT 126.2000 136.4000 126.6000 137.2000 ;
	    RECT 127.0000 136.2000 127.3000 137.5000 ;
	    RECT 129.1000 136.2000 129.5000 138.8000 ;
	    RECT 132.3000 139.2000 132.7000 139.9000 ;
	    RECT 134.7000 139.2000 135.7000 139.9000 ;
	    RECT 132.3000 138.8000 133.0000 139.2000 ;
	    RECT 134.7000 138.8000 136.2000 139.2000 ;
	    RECT 129.8000 136.8000 130.2000 137.2000 ;
	    RECT 129.9000 136.2000 130.2000 136.8000 ;
	    RECT 132.3000 136.3000 132.7000 138.8000 ;
	    RECT 124.6000 135.1000 125.0000 136.2000 ;
	    RECT 127.0000 135.8000 127.4000 136.2000 ;
	    RECT 129.1000 135.9000 129.6000 136.2000 ;
	    RECT 129.9000 135.9000 130.6000 136.2000 ;
	    RECT 131.8000 135.9000 132.7000 136.3000 ;
	    RECT 134.7000 135.9000 135.7000 138.8000 ;
	    RECT 138.5000 138.2000 138.9000 139.9000 ;
	    RECT 138.5000 137.8000 139.4000 138.2000 ;
	    RECT 137.8000 136.8000 138.2000 137.2000 ;
	    RECT 137.8000 136.2000 138.1000 136.8000 ;
	    RECT 138.5000 136.2000 138.9000 137.8000 ;
	    RECT 141.0000 136.8000 141.4000 137.2000 ;
	    RECT 141.0000 136.2000 141.3000 136.8000 ;
	    RECT 141.7000 136.2000 142.1000 139.9000 ;
	    RECT 137.4000 135.9000 138.1000 136.2000 ;
	    RECT 138.4000 135.9000 138.9000 136.2000 ;
	    RECT 140.6000 135.9000 141.3000 136.2000 ;
	    RECT 141.6000 135.9000 142.1000 136.2000 ;
	    RECT 144.1000 136.3000 144.5000 139.9000 ;
	    RECT 146.2000 137.9000 146.6000 139.9000 ;
	    RECT 146.3000 137.8000 146.6000 137.9000 ;
	    RECT 147.8000 137.9000 148.2000 139.9000 ;
	    RECT 147.8000 137.8000 148.1000 137.9000 ;
	    RECT 146.3000 137.5000 148.1000 137.8000 ;
	    RECT 144.1000 135.9000 145.0000 136.3000 ;
	    RECT 146.3000 136.2000 146.6000 137.5000 ;
	    RECT 147.0000 136.4000 147.4000 137.2000 ;
	    RECT 123.0000 134.8000 125.0000 135.1000 ;
	    RECT 125.4000 134.8000 126.2000 135.2000 ;
	    RECT 122.2000 134.1000 122.6000 134.2000 ;
	    RECT 120.6000 133.8000 122.6000 134.1000 ;
	    RECT 119.8000 132.4000 120.2000 133.2000 ;
	    RECT 120.6000 131.1000 121.0000 133.8000 ;
	    RECT 122.2000 133.4000 122.6000 133.8000 ;
	    RECT 121.4000 132.4000 121.8000 133.2000 ;
	    RECT 123.0000 133.1000 123.4000 134.8000 ;
	    RECT 127.0000 134.2000 127.3000 135.8000 ;
	    RECT 128.6000 134.4000 129.0000 135.2000 ;
	    RECT 129.3000 134.2000 129.6000 135.9000 ;
	    RECT 130.2000 135.8000 130.6000 135.9000 ;
	    RECT 131.9000 134.2000 132.2000 135.9000 ;
	    RECT 132.6000 134.8000 133.0000 135.6000 ;
	    RECT 134.2000 134.4000 134.6000 135.2000 ;
	    RECT 135.0000 134.2000 135.3000 135.9000 ;
	    RECT 137.4000 135.8000 137.8000 135.9000 ;
	    RECT 135.8000 134.4000 136.2000 135.2000 ;
	    RECT 126.5000 134.1000 127.3000 134.2000 ;
	    RECT 126.4000 133.9000 127.3000 134.1000 ;
	    RECT 127.8000 134.1000 128.2000 134.2000 ;
	    RECT 123.0000 132.8000 123.9000 133.1000 ;
	    RECT 123.5000 131.1000 123.9000 132.8000 ;
	    RECT 126.4000 131.1000 126.8000 133.9000 ;
	    RECT 127.8000 133.8000 128.6000 134.1000 ;
	    RECT 129.3000 133.8000 130.6000 134.2000 ;
	    RECT 131.8000 133.8000 132.2000 134.2000 ;
	    RECT 133.4000 134.1000 133.8000 134.2000 ;
	    RECT 135.0000 134.1000 135.4000 134.2000 ;
	    RECT 133.4000 133.8000 134.2000 134.1000 ;
	    RECT 135.0000 133.8000 136.2000 134.1000 ;
	    RECT 136.6000 133.8000 137.0000 134.6000 ;
	    RECT 138.4000 134.2000 138.7000 135.9000 ;
	    RECT 140.6000 135.8000 141.0000 135.9000 ;
	    RECT 139.0000 135.1000 139.4000 135.2000 ;
	    RECT 141.6000 135.1000 141.9000 135.9000 ;
	    RECT 139.0000 134.8000 141.9000 135.1000 ;
	    RECT 139.0000 134.4000 139.4000 134.8000 ;
	    RECT 141.6000 134.2000 141.9000 134.8000 ;
	    RECT 142.2000 134.4000 142.6000 135.2000 ;
	    RECT 143.8000 134.8000 144.2000 135.6000 ;
	    RECT 144.6000 134.2000 144.9000 135.9000 ;
	    RECT 146.2000 135.8000 146.6000 136.2000 ;
	    RECT 146.3000 134.2000 146.6000 135.8000 ;
	    RECT 147.4000 134.8000 148.2000 135.2000 ;
	    RECT 148.6000 135.1000 149.0000 136.2000 ;
	    RECT 149.4000 135.8000 149.8000 136.6000 ;
	    RECT 150.2000 135.1000 150.6000 139.9000 ;
	    RECT 152.9000 139.2000 153.3000 139.9000 ;
	    RECT 152.9000 138.8000 153.8000 139.2000 ;
	    RECT 152.2000 136.8000 152.6000 137.2000 ;
	    RECT 152.2000 136.2000 152.5000 136.8000 ;
	    RECT 152.9000 136.2000 153.3000 138.8000 ;
	    RECT 151.8000 135.9000 152.5000 136.2000 ;
	    RECT 152.8000 135.9000 153.3000 136.2000 ;
	    RECT 155.0000 135.9000 155.4000 139.9000 ;
	    RECT 156.6000 137.9000 157.0000 139.9000 ;
	    RECT 159.0000 137.9000 159.4000 139.9000 ;
	    RECT 151.8000 135.8000 152.2000 135.9000 ;
	    RECT 148.6000 134.8000 150.6000 135.1000 ;
	    RECT 137.4000 133.8000 138.7000 134.2000 ;
	    RECT 139.8000 134.1000 140.2000 134.2000 ;
	    RECT 139.4000 133.8000 140.2000 134.1000 ;
	    RECT 140.6000 133.8000 141.9000 134.2000 ;
	    RECT 143.0000 134.1000 143.4000 134.2000 ;
	    RECT 144.6000 134.1000 145.0000 134.2000 ;
	    RECT 142.6000 133.8000 143.4000 134.1000 ;
	    RECT 143.8000 133.8000 145.0000 134.1000 ;
	    RECT 146.3000 134.1000 147.1000 134.2000 ;
	    RECT 146.3000 133.9000 147.2000 134.1000 ;
	    RECT 128.2000 133.6000 128.6000 133.8000 ;
	    RECT 127.9000 133.1000 129.7000 133.3000 ;
	    RECT 130.2000 133.1000 130.5000 133.8000 ;
	    RECT 127.8000 133.0000 129.8000 133.1000 ;
	    RECT 127.8000 131.1000 128.2000 133.0000 ;
	    RECT 129.4000 131.1000 129.8000 133.0000 ;
	    RECT 130.2000 131.1000 130.6000 133.1000 ;
	    RECT 131.0000 132.4000 131.4000 133.2000 ;
	    RECT 131.9000 132.1000 132.2000 133.8000 ;
	    RECT 133.8000 133.6000 134.2000 133.8000 ;
	    RECT 133.5000 133.1000 135.3000 133.3000 ;
	    RECT 135.9000 133.1000 136.2000 133.8000 ;
	    RECT 137.5000 133.1000 137.8000 133.8000 ;
	    RECT 139.4000 133.6000 139.8000 133.8000 ;
	    RECT 138.3000 133.1000 140.1000 133.3000 ;
	    RECT 140.7000 133.1000 141.0000 133.8000 ;
	    RECT 142.6000 133.6000 143.0000 133.8000 ;
	    RECT 141.5000 133.1000 143.3000 133.3000 ;
	    RECT 143.8000 133.2000 144.1000 133.8000 ;
	    RECT 131.8000 131.1000 132.2000 132.1000 ;
	    RECT 133.4000 133.0000 135.4000 133.1000 ;
	    RECT 133.4000 131.1000 133.8000 133.0000 ;
	    RECT 135.0000 131.4000 135.4000 133.0000 ;
	    RECT 135.8000 131.7000 136.2000 133.1000 ;
	    RECT 136.6000 131.4000 137.0000 133.1000 ;
	    RECT 135.0000 131.1000 137.0000 131.4000 ;
	    RECT 137.4000 131.1000 137.8000 133.1000 ;
	    RECT 138.2000 133.0000 140.2000 133.1000 ;
	    RECT 138.2000 131.1000 138.6000 133.0000 ;
	    RECT 139.8000 131.1000 140.2000 133.0000 ;
	    RECT 140.6000 131.1000 141.0000 133.1000 ;
	    RECT 141.4000 133.0000 143.4000 133.1000 ;
	    RECT 141.4000 131.1000 141.8000 133.0000 ;
	    RECT 143.0000 131.1000 143.4000 133.0000 ;
	    RECT 143.8000 132.8000 144.2000 133.2000 ;
	    RECT 144.6000 132.1000 144.9000 133.8000 ;
	    RECT 145.4000 132.4000 145.8000 133.2000 ;
	    RECT 144.6000 131.1000 145.0000 132.1000 ;
	    RECT 146.8000 131.1000 147.2000 133.9000 ;
	    RECT 150.2000 133.1000 150.6000 134.8000 ;
	    RECT 152.8000 134.2000 153.1000 135.9000 ;
	    RECT 155.0000 135.2000 155.3000 135.9000 ;
	    RECT 156.6000 135.8000 156.9000 137.9000 ;
	    RECT 159.1000 137.8000 159.4000 137.9000 ;
	    RECT 160.6000 137.9000 161.0000 139.9000 ;
	    RECT 160.6000 137.8000 160.9000 137.9000 ;
	    RECT 159.1000 137.5000 160.9000 137.8000 ;
	    RECT 158.2000 137.1000 158.6000 137.2000 ;
	    RECT 159.8000 137.1000 160.2000 137.2000 ;
	    RECT 158.2000 136.8000 160.2000 137.1000 ;
	    RECT 159.8000 136.4000 160.2000 136.8000 ;
	    RECT 160.6000 136.2000 160.9000 137.5000 ;
	    RECT 155.7000 135.5000 156.9000 135.8000 ;
	    RECT 153.4000 134.4000 153.8000 135.2000 ;
	    RECT 155.0000 134.8000 155.4000 135.2000 ;
	    RECT 151.0000 133.4000 151.4000 134.2000 ;
	    RECT 151.8000 133.8000 153.1000 134.2000 ;
	    RECT 154.2000 134.1000 154.6000 134.2000 ;
	    RECT 153.8000 133.8000 154.6000 134.1000 ;
	    RECT 151.9000 133.1000 152.2000 133.8000 ;
	    RECT 153.8000 133.6000 154.2000 133.8000 ;
	    RECT 152.7000 133.1000 154.5000 133.3000 ;
	    RECT 155.0000 133.1000 155.3000 134.8000 ;
	    RECT 155.7000 133.8000 156.0000 135.5000 ;
	    RECT 158.2000 135.4000 158.6000 136.2000 ;
	    RECT 160.6000 135.8000 161.0000 136.2000 ;
	    RECT 156.6000 134.8000 157.0000 135.2000 ;
	    RECT 159.0000 134.8000 159.8000 135.2000 ;
	    RECT 156.6000 134.4000 156.9000 134.8000 ;
	    RECT 156.4000 134.0000 157.0000 134.4000 ;
	    RECT 157.4000 133.8000 157.8000 134.6000 ;
	    RECT 160.6000 134.2000 160.9000 135.8000 ;
	    RECT 160.1000 134.1000 160.9000 134.2000 ;
	    RECT 160.0000 133.9000 160.9000 134.1000 ;
	    RECT 162.2000 134.1000 162.6000 139.9000 ;
	    RECT 163.0000 135.8000 163.4000 139.9000 ;
	    RECT 163.8000 136.2000 164.2000 139.9000 ;
	    RECT 165.4000 136.2000 165.8000 139.9000 ;
	    RECT 167.5000 139.2000 167.9000 139.9000 ;
	    RECT 167.0000 138.8000 167.9000 139.2000 ;
	    RECT 163.8000 135.9000 165.8000 136.2000 ;
	    RECT 167.5000 136.2000 167.9000 138.8000 ;
	    RECT 168.2000 136.8000 168.6000 137.2000 ;
	    RECT 168.3000 136.2000 168.6000 136.8000 ;
	    RECT 170.7000 136.2000 171.1000 139.9000 ;
	    RECT 171.4000 136.8000 171.8000 137.2000 ;
	    RECT 171.5000 136.2000 171.8000 136.8000 ;
	    RECT 167.5000 135.9000 168.0000 136.2000 ;
	    RECT 168.3000 135.9000 169.0000 136.2000 ;
	    RECT 170.7000 135.9000 171.2000 136.2000 ;
	    RECT 171.5000 135.9000 172.2000 136.2000 ;
	    RECT 163.1000 135.2000 163.4000 135.8000 ;
	    RECT 165.0000 135.2000 165.4000 135.4000 ;
	    RECT 163.0000 134.9000 164.2000 135.2000 ;
	    RECT 165.0000 134.9000 165.8000 135.2000 ;
	    RECT 163.0000 134.8000 163.4000 134.9000 ;
	    RECT 163.0000 134.1000 163.4000 134.2000 ;
	    RECT 155.6000 133.7000 156.0000 133.8000 ;
	    RECT 155.6000 133.5000 157.1000 133.7000 ;
	    RECT 155.6000 133.4000 157.7000 133.5000 ;
	    RECT 156.8000 133.2000 157.7000 133.4000 ;
	    RECT 157.4000 133.1000 157.7000 133.2000 ;
	    RECT 149.7000 132.8000 150.6000 133.1000 ;
	    RECT 149.7000 131.1000 150.1000 132.8000 ;
	    RECT 151.8000 131.1000 152.2000 133.1000 ;
	    RECT 152.6000 133.0000 154.6000 133.1000 ;
	    RECT 152.6000 131.1000 153.0000 133.0000 ;
	    RECT 154.2000 131.1000 154.6000 133.0000 ;
	    RECT 155.0000 132.6000 155.7000 133.1000 ;
	    RECT 155.3000 131.1000 155.7000 132.6000 ;
	    RECT 157.4000 131.1000 157.8000 133.1000 ;
	    RECT 160.0000 131.1000 160.4000 133.9000 ;
	    RECT 162.2000 133.8000 163.4000 134.1000 ;
	    RECT 161.4000 132.4000 161.8000 133.2000 ;
	    RECT 162.2000 131.1000 162.6000 133.8000 ;
	    RECT 163.0000 132.8000 163.4000 133.2000 ;
	    RECT 163.9000 133.1000 164.2000 134.9000 ;
	    RECT 165.4000 134.8000 165.8000 134.9000 ;
	    RECT 164.6000 133.8000 165.0000 134.6000 ;
	    RECT 167.0000 134.4000 167.4000 135.2000 ;
	    RECT 167.7000 135.1000 168.0000 135.9000 ;
	    RECT 168.6000 135.8000 169.0000 135.9000 ;
	    RECT 170.2000 135.1000 170.6000 135.2000 ;
	    RECT 167.7000 134.8000 170.6000 135.1000 ;
	    RECT 167.7000 134.2000 168.0000 134.8000 ;
	    RECT 170.2000 134.4000 170.6000 134.8000 ;
	    RECT 170.9000 134.2000 171.2000 135.9000 ;
	    RECT 171.8000 135.8000 172.2000 135.9000 ;
	    RECT 166.2000 134.1000 166.6000 134.2000 ;
	    RECT 166.2000 133.8000 167.0000 134.1000 ;
	    RECT 167.7000 133.8000 169.0000 134.2000 ;
	    RECT 169.4000 134.1000 169.8000 134.2000 ;
	    RECT 169.4000 133.8000 170.2000 134.1000 ;
	    RECT 170.9000 133.8000 172.2000 134.2000 ;
	    RECT 166.6000 133.6000 167.0000 133.8000 ;
	    RECT 166.3000 133.1000 168.1000 133.3000 ;
	    RECT 168.6000 133.1000 168.9000 133.8000 ;
	    RECT 169.8000 133.6000 170.2000 133.8000 ;
	    RECT 169.5000 133.1000 171.3000 133.3000 ;
	    RECT 171.8000 133.1000 172.1000 133.8000 ;
	    RECT 163.1000 132.4000 163.5000 132.8000 ;
	    RECT 163.8000 131.1000 164.2000 133.1000 ;
	    RECT 166.2000 133.0000 168.2000 133.1000 ;
	    RECT 166.2000 131.1000 166.6000 133.0000 ;
	    RECT 167.8000 131.1000 168.2000 133.0000 ;
	    RECT 168.6000 131.1000 169.0000 133.1000 ;
	    RECT 169.4000 133.0000 171.4000 133.1000 ;
	    RECT 169.4000 131.1000 169.8000 133.0000 ;
	    RECT 171.0000 131.1000 171.4000 133.0000 ;
	    RECT 171.8000 131.1000 172.2000 133.1000 ;
	    RECT 1.4000 121.1000 1.8000 129.9000 ;
	    RECT 3.6000 127.1000 4.0000 129.9000 ;
	    RECT 3.1000 126.9000 4.0000 127.1000 ;
	    RECT 3.1000 126.8000 3.9000 126.9000 ;
	    RECT 3.1000 125.2000 3.4000 126.8000 ;
	    RECT 4.2000 125.8000 5.0000 126.2000 ;
	    RECT 3.0000 124.8000 3.4000 125.2000 ;
	    RECT 3.1000 123.5000 3.4000 124.8000 ;
	    RECT 3.8000 123.8000 4.2000 124.6000 ;
	    RECT 3.1000 123.2000 4.9000 123.5000 ;
	    RECT 3.1000 123.1000 3.4000 123.2000 ;
	    RECT 3.0000 121.1000 3.4000 123.1000 ;
	    RECT 4.6000 123.1000 4.9000 123.2000 ;
	    RECT 4.6000 121.1000 5.0000 123.1000 ;
	    RECT 7.0000 121.1000 7.4000 129.9000 ;
	    RECT 10.4000 127.1000 10.8000 129.9000 ;
	    RECT 13.6000 127.1000 14.0000 129.9000 ;
	    RECT 15.6000 127.1000 16.0000 129.9000 ;
	    RECT 18.8000 127.1000 19.2000 129.9000 ;
	    RECT 10.4000 126.9000 11.3000 127.1000 ;
	    RECT 13.6000 126.9000 14.5000 127.1000 ;
	    RECT 10.5000 126.8000 11.3000 126.9000 ;
	    RECT 13.7000 126.8000 14.5000 126.9000 ;
	    RECT 9.4000 125.8000 10.2000 126.2000 ;
	    RECT 11.0000 125.2000 11.3000 126.8000 ;
	    RECT 12.6000 125.8000 13.4000 126.2000 ;
	    RECT 14.2000 125.2000 14.5000 126.8000 ;
	    RECT 15.1000 126.9000 16.0000 127.1000 ;
	    RECT 18.3000 126.9000 19.2000 127.1000 ;
	    RECT 21.4000 127.9000 21.8000 129.9000 ;
	    RECT 23.0000 128.9000 23.4000 129.9000 ;
	    RECT 25.4000 128.9000 25.8000 129.9000 ;
	    RECT 15.1000 126.8000 15.9000 126.9000 ;
	    RECT 18.3000 126.8000 19.1000 126.9000 ;
	    RECT 15.1000 125.2000 15.4000 126.8000 ;
	    RECT 16.2000 125.8000 17.0000 126.2000 ;
	    RECT 11.0000 124.8000 11.4000 125.2000 ;
	    RECT 14.2000 124.8000 14.6000 125.2000 ;
	    RECT 15.0000 124.8000 15.4000 125.2000 ;
	    RECT 17.4000 124.8000 17.8000 125.6000 ;
	    RECT 18.3000 125.2000 18.6000 126.8000 ;
	    RECT 21.4000 126.2000 21.7000 127.9000 ;
	    RECT 23.0000 127.8000 23.3000 128.9000 ;
	    RECT 23.8000 128.1000 24.2000 128.6000 ;
	    RECT 24.6000 128.1000 25.0000 128.6000 ;
	    RECT 23.8000 127.8000 25.0000 128.1000 ;
	    RECT 25.5000 127.8000 25.8000 128.9000 ;
	    RECT 27.0000 127.9000 27.4000 129.9000 ;
	    RECT 22.1000 127.5000 23.3000 127.8000 ;
	    RECT 25.5000 127.5000 26.7000 127.8000 ;
	    RECT 19.4000 125.8000 20.2000 126.2000 ;
	    RECT 21.4000 125.8000 21.8000 126.2000 ;
	    RECT 22.1000 126.0000 22.4000 127.5000 ;
	    RECT 26.4000 126.0000 26.7000 127.5000 ;
	    RECT 27.1000 126.2000 27.4000 127.9000 ;
	    RECT 28.4000 127.2000 28.8000 129.9000 ;
	    RECT 29.4000 127.8000 29.8000 128.2000 ;
	    RECT 28.4000 127.1000 29.0000 127.2000 ;
	    RECT 29.4000 127.1000 29.7000 127.8000 ;
	    RECT 31.6000 127.1000 32.0000 129.9000 ;
	    RECT 18.2000 124.8000 18.6000 125.2000 ;
	    RECT 21.4000 125.1000 21.7000 125.8000 ;
	    RECT 22.1000 125.7000 22.5000 126.0000 ;
	    RECT 26.3000 125.7000 26.7000 126.0000 ;
	    RECT 27.0000 125.8000 27.4000 126.2000 ;
	    RECT 22.1000 125.6000 24.2000 125.7000 ;
	    RECT 22.2000 125.4000 24.2000 125.6000 ;
	    RECT 21.4000 124.8000 22.1000 125.1000 ;
	    RECT 10.2000 123.8000 10.6000 124.6000 ;
	    RECT 11.0000 123.5000 11.3000 124.8000 ;
	    RECT 13.4000 123.8000 13.8000 124.6000 ;
	    RECT 14.2000 123.5000 14.5000 124.8000 ;
	    RECT 9.5000 123.2000 11.3000 123.5000 ;
	    RECT 9.5000 123.1000 9.8000 123.2000 ;
	    RECT 9.4000 121.1000 9.8000 123.1000 ;
	    RECT 11.0000 123.1000 11.3000 123.2000 ;
	    RECT 12.7000 123.2000 14.5000 123.5000 ;
	    RECT 12.7000 123.1000 13.0000 123.2000 ;
	    RECT 11.0000 121.1000 11.4000 123.1000 ;
	    RECT 12.6000 121.1000 13.0000 123.1000 ;
	    RECT 14.2000 123.1000 14.5000 123.2000 ;
	    RECT 15.1000 123.5000 15.4000 124.8000 ;
	    RECT 15.8000 123.8000 16.2000 124.6000 ;
	    RECT 18.3000 123.5000 18.6000 124.8000 ;
	    RECT 19.0000 123.8000 19.4000 124.6000 ;
	    RECT 15.1000 123.2000 16.9000 123.5000 ;
	    RECT 18.3000 123.2000 20.1000 123.5000 ;
	    RECT 15.1000 123.1000 15.4000 123.2000 ;
	    RECT 14.2000 121.1000 14.6000 123.1000 ;
	    RECT 15.0000 121.1000 15.4000 123.1000 ;
	    RECT 16.6000 121.1000 17.0000 123.2000 ;
	    RECT 18.3000 123.1000 18.6000 123.2000 ;
	    RECT 18.2000 121.1000 18.6000 123.1000 ;
	    RECT 19.8000 123.1000 20.1000 123.2000 ;
	    RECT 19.8000 121.1000 20.2000 123.1000 ;
	    RECT 21.7000 121.1000 22.1000 124.8000 ;
	    RECT 23.8000 121.1000 24.2000 125.4000 ;
	    RECT 24.6000 125.6000 26.7000 125.7000 ;
	    RECT 24.6000 125.4000 26.6000 125.6000 ;
	    RECT 24.6000 121.1000 25.0000 125.4000 ;
	    RECT 27.1000 125.1000 27.4000 125.8000 ;
	    RECT 27.9000 126.8000 29.7000 127.1000 ;
	    RECT 31.1000 126.9000 32.0000 127.1000 ;
	    RECT 36.0000 127.1000 36.4000 129.9000 ;
	    RECT 37.7000 128.2000 38.1000 129.9000 ;
	    RECT 37.7000 127.9000 38.6000 128.2000 ;
	    RECT 36.0000 126.9000 36.9000 127.1000 ;
	    RECT 31.1000 126.8000 31.9000 126.9000 ;
	    RECT 36.1000 126.8000 36.9000 126.9000 ;
	    RECT 27.9000 125.2000 28.2000 126.8000 ;
	    RECT 29.0000 125.8000 29.8000 126.2000 ;
	    RECT 26.7000 124.8000 27.4000 125.1000 ;
	    RECT 27.8000 124.8000 28.2000 125.2000 ;
	    RECT 30.2000 124.8000 30.6000 125.6000 ;
	    RECT 31.1000 125.2000 31.4000 126.8000 ;
	    RECT 32.2000 125.8000 33.0000 126.2000 ;
	    RECT 35.0000 125.8000 35.8000 126.2000 ;
	    RECT 31.0000 124.8000 31.4000 125.2000 ;
	    RECT 34.2000 124.8000 34.6000 125.6000 ;
	    RECT 36.6000 125.2000 36.9000 126.8000 ;
	    RECT 36.6000 124.8000 37.0000 125.2000 ;
	    RECT 26.7000 121.1000 27.1000 124.8000 ;
	    RECT 27.9000 123.5000 28.2000 124.8000 ;
	    RECT 28.6000 123.8000 29.0000 124.6000 ;
	    RECT 31.1000 123.5000 31.4000 124.8000 ;
	    RECT 31.8000 123.8000 32.2000 124.6000 ;
	    RECT 35.8000 123.8000 36.2000 124.6000 ;
	    RECT 36.6000 123.5000 36.9000 124.8000 ;
	    RECT 37.4000 124.4000 37.8000 125.2000 ;
	    RECT 27.9000 123.2000 29.7000 123.5000 ;
	    RECT 27.9000 123.1000 28.2000 123.2000 ;
	    RECT 27.8000 121.1000 28.2000 123.1000 ;
	    RECT 29.4000 123.1000 29.7000 123.2000 ;
	    RECT 31.1000 123.2000 32.9000 123.5000 ;
	    RECT 31.1000 123.1000 31.4000 123.2000 ;
	    RECT 29.4000 121.1000 29.8000 123.1000 ;
	    RECT 31.0000 121.1000 31.4000 123.1000 ;
	    RECT 32.6000 123.1000 32.9000 123.2000 ;
	    RECT 35.1000 123.2000 36.9000 123.5000 ;
	    RECT 35.1000 123.1000 35.4000 123.2000 ;
	    RECT 32.6000 121.1000 33.0000 123.1000 ;
	    RECT 35.0000 121.1000 35.4000 123.1000 ;
	    RECT 36.6000 123.1000 36.9000 123.2000 ;
	    RECT 38.2000 124.1000 38.6000 127.9000 ;
	    RECT 39.0000 126.8000 39.4000 127.6000 ;
	    RECT 39.0000 125.8000 39.4000 126.2000 ;
	    RECT 39.0000 125.1000 39.3000 125.8000 ;
	    RECT 39.8000 125.1000 40.2000 129.9000 ;
	    RECT 41.7000 128.2000 42.1000 129.9000 ;
	    RECT 44.6000 128.9000 45.0000 129.9000 ;
	    RECT 41.7000 127.9000 42.6000 128.2000 ;
	    RECT 39.0000 124.8000 40.2000 125.1000 ;
	    RECT 39.0000 124.1000 39.4000 124.2000 ;
	    RECT 38.2000 123.8000 39.4000 124.1000 ;
	    RECT 36.6000 121.1000 37.0000 123.1000 ;
	    RECT 38.2000 121.1000 38.6000 123.8000 ;
	    RECT 39.8000 121.1000 40.2000 124.8000 ;
	    RECT 41.4000 124.4000 41.8000 125.2000 ;
	    RECT 42.2000 124.1000 42.6000 127.9000 ;
	    RECT 43.8000 127.8000 44.2000 128.6000 ;
	    RECT 44.7000 127.8000 45.0000 128.9000 ;
	    RECT 46.2000 127.9000 46.6000 129.9000 ;
	    RECT 43.0000 127.1000 43.4000 127.6000 ;
	    RECT 43.8000 127.1000 44.1000 127.8000 ;
	    RECT 44.7000 127.5000 45.9000 127.8000 ;
	    RECT 43.0000 126.8000 44.1000 127.1000 ;
	    RECT 45.6000 126.0000 45.9000 127.5000 ;
	    RECT 46.3000 126.2000 46.6000 127.9000 ;
	    RECT 47.6000 127.1000 48.0000 129.9000 ;
	    RECT 51.0000 128.9000 51.4000 129.9000 ;
	    RECT 50.2000 127.8000 50.6000 128.6000 ;
	    RECT 51.1000 127.8000 51.4000 128.9000 ;
	    RECT 52.6000 127.9000 53.0000 129.9000 ;
	    RECT 51.1000 127.5000 52.3000 127.8000 ;
	    RECT 45.5000 125.7000 45.9000 126.0000 ;
	    RECT 46.2000 125.8000 46.6000 126.2000 ;
	    RECT 43.8000 125.6000 45.9000 125.7000 ;
	    RECT 43.8000 125.4000 45.8000 125.6000 ;
	    RECT 43.0000 124.8000 43.4000 125.2000 ;
	    RECT 43.0000 124.1000 43.3000 124.8000 ;
	    RECT 42.2000 123.8000 43.3000 124.1000 ;
	    RECT 42.2000 121.1000 42.6000 123.8000 ;
	    RECT 43.8000 121.1000 44.2000 125.4000 ;
	    RECT 46.3000 125.1000 46.6000 125.8000 ;
	    RECT 47.1000 126.9000 48.0000 127.1000 ;
	    RECT 47.1000 126.8000 47.9000 126.9000 ;
	    RECT 47.1000 125.2000 47.4000 126.8000 ;
	    RECT 48.2000 125.8000 49.0000 126.2000 ;
	    RECT 52.0000 126.0000 52.3000 127.5000 ;
	    RECT 52.7000 126.2000 53.0000 127.9000 ;
	    RECT 54.0000 127.1000 54.4000 129.9000 ;
	    RECT 51.9000 125.7000 52.3000 126.0000 ;
	    RECT 52.6000 125.8000 53.0000 126.2000 ;
	    RECT 50.2000 125.6000 52.3000 125.7000 ;
	    RECT 45.9000 124.8000 46.6000 125.1000 ;
	    RECT 47.0000 124.8000 47.4000 125.2000 ;
	    RECT 49.4000 124.8000 49.8000 125.6000 ;
	    RECT 50.2000 125.4000 52.2000 125.6000 ;
	    RECT 45.9000 121.1000 46.3000 124.8000 ;
	    RECT 47.1000 123.5000 47.4000 124.8000 ;
	    RECT 47.8000 123.8000 48.2000 124.6000 ;
	    RECT 47.1000 123.2000 48.9000 123.5000 ;
	    RECT 47.1000 123.1000 47.4000 123.2000 ;
	    RECT 47.0000 121.1000 47.4000 123.1000 ;
	    RECT 48.6000 123.1000 48.9000 123.2000 ;
	    RECT 48.6000 121.1000 49.0000 123.1000 ;
	    RECT 50.2000 121.1000 50.6000 125.4000 ;
	    RECT 52.7000 125.1000 53.0000 125.8000 ;
	    RECT 53.5000 126.9000 54.4000 127.1000 ;
	    RECT 53.5000 126.8000 54.3000 126.9000 ;
	    RECT 53.5000 125.2000 53.8000 126.8000 ;
	    RECT 56.6000 126.2000 57.0000 129.9000 ;
	    RECT 58.2000 127.6000 58.6000 129.9000 ;
	    RECT 57.5000 127.3000 58.6000 127.6000 ;
	    RECT 54.6000 125.8000 55.4000 126.2000 ;
	    RECT 52.3000 124.8000 53.0000 125.1000 ;
	    RECT 53.4000 124.8000 53.8000 125.2000 ;
	    RECT 55.8000 124.8000 56.2000 125.6000 ;
	    RECT 56.6000 125.1000 56.9000 126.2000 ;
	    RECT 57.5000 125.8000 57.8000 127.3000 ;
	    RECT 61.2000 127.1000 61.6000 129.9000 ;
	    RECT 64.6000 128.9000 65.0000 129.9000 ;
	    RECT 63.8000 127.8000 64.2000 128.6000 ;
	    RECT 64.7000 127.8000 65.0000 128.9000 ;
	    RECT 66.2000 127.9000 66.6000 129.9000 ;
	    RECT 64.7000 127.5000 65.9000 127.8000 ;
	    RECT 57.2000 125.4000 57.8000 125.8000 ;
	    RECT 57.5000 125.1000 57.8000 125.4000 ;
	    RECT 60.7000 126.9000 61.6000 127.1000 ;
	    RECT 60.7000 126.8000 61.5000 126.9000 ;
	    RECT 60.7000 125.2000 61.0000 126.8000 ;
	    RECT 61.8000 125.8000 62.6000 126.2000 ;
	    RECT 65.6000 126.0000 65.9000 127.5000 ;
	    RECT 66.3000 127.2000 66.6000 127.9000 ;
	    RECT 66.2000 126.8000 66.6000 127.2000 ;
	    RECT 68.8000 127.1000 69.2000 129.9000 ;
	    RECT 72.0000 127.1000 72.4000 129.9000 ;
	    RECT 74.7000 128.2000 75.1000 129.9000 ;
	    RECT 74.2000 127.9000 75.1000 128.2000 ;
	    RECT 68.8000 126.9000 69.7000 127.1000 ;
	    RECT 72.0000 126.9000 72.9000 127.1000 ;
	    RECT 68.9000 126.8000 69.7000 126.9000 ;
	    RECT 72.1000 126.8000 72.9000 126.9000 ;
	    RECT 73.4000 126.8000 73.8000 127.6000 ;
	    RECT 66.3000 126.2000 66.6000 126.8000 ;
	    RECT 65.5000 125.7000 65.9000 126.0000 ;
	    RECT 66.2000 125.8000 66.6000 126.2000 ;
	    RECT 67.8000 125.8000 68.6000 126.2000 ;
	    RECT 52.3000 121.1000 52.7000 124.8000 ;
	    RECT 53.5000 123.5000 53.8000 124.8000 ;
	    RECT 54.2000 123.8000 54.6000 124.6000 ;
	    RECT 55.0000 123.8000 55.4000 124.2000 ;
	    RECT 55.0000 123.5000 55.3000 123.8000 ;
	    RECT 53.5000 123.2000 55.3000 123.5000 ;
	    RECT 53.5000 123.1000 53.8000 123.2000 ;
	    RECT 53.4000 121.1000 53.8000 123.1000 ;
	    RECT 55.0000 123.1000 55.3000 123.2000 ;
	    RECT 55.0000 121.1000 55.4000 123.1000 ;
	    RECT 56.6000 121.1000 57.0000 125.1000 ;
	    RECT 57.5000 124.8000 58.6000 125.1000 ;
	    RECT 60.6000 124.8000 61.0000 125.2000 ;
	    RECT 58.2000 121.1000 58.6000 124.8000 ;
	    RECT 60.7000 123.5000 61.0000 124.8000 ;
	    RECT 63.8000 125.6000 65.9000 125.7000 ;
	    RECT 63.8000 125.4000 65.8000 125.6000 ;
	    RECT 61.4000 123.8000 61.8000 124.6000 ;
	    RECT 60.7000 123.2000 62.5000 123.5000 ;
	    RECT 60.7000 123.1000 61.0000 123.2000 ;
	    RECT 60.6000 121.1000 61.0000 123.1000 ;
	    RECT 62.2000 123.1000 62.5000 123.2000 ;
	    RECT 62.2000 121.1000 62.6000 123.1000 ;
	    RECT 63.8000 121.1000 64.2000 125.4000 ;
	    RECT 66.3000 125.1000 66.6000 125.8000 ;
	    RECT 65.9000 124.8000 66.6000 125.1000 ;
	    RECT 67.0000 124.8000 67.4000 125.6000 ;
	    RECT 69.4000 125.2000 69.7000 126.8000 ;
	    RECT 71.0000 125.8000 71.8000 126.2000 ;
	    RECT 69.4000 124.8000 69.8000 125.2000 ;
	    RECT 70.2000 125.1000 70.6000 125.6000 ;
	    RECT 72.6000 125.2000 72.9000 126.8000 ;
	    RECT 74.2000 126.1000 74.6000 127.9000 ;
	    RECT 73.4000 125.8000 74.6000 126.1000 ;
	    RECT 73.4000 125.2000 73.7000 125.8000 ;
	    RECT 71.0000 125.1000 71.4000 125.2000 ;
	    RECT 70.2000 124.8000 71.4000 125.1000 ;
	    RECT 72.6000 124.8000 73.0000 125.2000 ;
	    RECT 73.4000 124.8000 73.8000 125.2000 ;
	    RECT 65.9000 121.1000 66.3000 124.8000 ;
	    RECT 68.6000 123.8000 69.0000 124.6000 ;
	    RECT 69.4000 123.5000 69.7000 124.8000 ;
	    RECT 71.8000 123.8000 72.2000 124.6000 ;
	    RECT 72.6000 123.5000 72.9000 124.8000 ;
	    RECT 67.9000 123.2000 69.7000 123.5000 ;
	    RECT 67.9000 123.1000 68.2000 123.2000 ;
	    RECT 67.8000 121.1000 68.2000 123.1000 ;
	    RECT 69.4000 123.1000 69.7000 123.2000 ;
	    RECT 71.1000 123.2000 72.9000 123.5000 ;
	    RECT 71.1000 123.1000 71.4000 123.2000 ;
	    RECT 69.4000 121.1000 69.8000 123.1000 ;
	    RECT 71.0000 121.1000 71.4000 123.1000 ;
	    RECT 72.6000 123.1000 72.9000 123.2000 ;
	    RECT 72.6000 121.1000 73.0000 123.1000 ;
	    RECT 74.2000 121.1000 74.6000 125.8000 ;
	    RECT 75.0000 125.1000 75.4000 125.2000 ;
	    RECT 75.8000 125.1000 76.2000 129.9000 ;
	    RECT 79.2000 127.1000 79.6000 129.9000 ;
	    RECT 79.2000 126.9000 80.1000 127.1000 ;
	    RECT 79.3000 126.8000 80.1000 126.9000 ;
	    RECT 78.2000 125.8000 79.0000 126.2000 ;
	    RECT 75.0000 124.8000 76.2000 125.1000 ;
	    RECT 75.0000 124.4000 75.4000 124.8000 ;
	    RECT 75.8000 121.1000 76.2000 124.8000 ;
	    RECT 79.8000 125.2000 80.1000 126.8000 ;
	    RECT 79.8000 124.8000 80.2000 125.2000 ;
	    RECT 79.0000 123.8000 79.4000 124.6000 ;
	    RECT 79.8000 123.5000 80.1000 124.8000 ;
	    RECT 78.3000 123.2000 80.1000 123.5000 ;
	    RECT 78.3000 123.1000 78.6000 123.2000 ;
	    RECT 78.2000 121.1000 78.6000 123.1000 ;
	    RECT 79.8000 123.1000 80.1000 123.2000 ;
	    RECT 79.8000 121.1000 80.2000 123.1000 ;
	    RECT 81.4000 121.1000 81.8000 129.9000 ;
	    RECT 83.3000 129.2000 83.7000 129.9000 ;
	    RECT 83.0000 128.8000 83.7000 129.2000 ;
	    RECT 83.3000 128.2000 83.7000 128.8000 ;
	    RECT 83.3000 127.9000 84.2000 128.2000 ;
	    RECT 83.0000 124.4000 83.4000 125.2000 ;
	    RECT 83.8000 121.1000 84.2000 127.9000 ;
	    RECT 85.4000 127.7000 85.8000 129.9000 ;
	    RECT 87.5000 129.2000 88.1000 129.9000 ;
	    RECT 87.5000 128.9000 88.2000 129.2000 ;
	    RECT 89.8000 128.9000 90.2000 129.9000 ;
	    RECT 92.0000 129.2000 92.4000 129.9000 ;
	    RECT 92.0000 128.9000 93.0000 129.2000 ;
	    RECT 87.8000 128.5000 88.2000 128.9000 ;
	    RECT 89.9000 128.6000 90.2000 128.9000 ;
	    RECT 89.9000 128.3000 91.3000 128.6000 ;
	    RECT 90.9000 128.2000 91.3000 128.3000 ;
	    RECT 91.8000 128.2000 92.2000 128.6000 ;
	    RECT 92.6000 128.5000 93.0000 128.9000 ;
	    RECT 86.9000 127.7000 87.3000 127.8000 ;
	    RECT 84.6000 126.8000 85.0000 127.6000 ;
	    RECT 85.4000 127.4000 87.3000 127.7000 ;
	    RECT 85.4000 125.7000 85.8000 127.4000 ;
	    RECT 88.9000 127.1000 89.3000 127.2000 ;
	    RECT 91.8000 127.1000 92.1000 128.2000 ;
	    RECT 94.2000 127.5000 94.6000 129.9000 ;
	    RECT 95.0000 127.8000 95.4000 128.6000 ;
	    RECT 93.4000 127.1000 94.2000 127.2000 ;
	    RECT 88.7000 126.8000 94.2000 127.1000 ;
	    RECT 95.8000 127.1000 96.2000 129.9000 ;
	    RECT 97.9000 129.2000 98.3000 129.9000 ;
	    RECT 99.3000 129.2000 99.7000 129.9000 ;
	    RECT 97.4000 128.8000 98.3000 129.2000 ;
	    RECT 99.0000 128.8000 99.7000 129.2000 ;
	    RECT 97.9000 128.2000 98.3000 128.8000 ;
	    RECT 97.4000 127.9000 98.3000 128.2000 ;
	    RECT 99.3000 128.2000 99.7000 128.8000 ;
	    RECT 102.7000 129.2000 103.1000 129.9000 ;
	    RECT 102.7000 128.8000 103.4000 129.2000 ;
	    RECT 102.7000 128.2000 103.1000 128.8000 ;
	    RECT 99.3000 127.9000 100.2000 128.2000 ;
	    RECT 96.6000 127.1000 97.0000 127.6000 ;
	    RECT 95.8000 126.8000 97.0000 127.1000 ;
	    RECT 87.8000 126.4000 88.2000 126.5000 ;
	    RECT 86.3000 126.1000 88.2000 126.4000 ;
	    RECT 88.7000 126.2000 89.0000 126.8000 ;
	    RECT 92.3000 126.7000 92.7000 126.8000 ;
	    RECT 91.8000 126.2000 92.2000 126.3000 ;
	    RECT 93.1000 126.2000 93.5000 126.3000 ;
	    RECT 86.3000 126.0000 86.7000 126.1000 ;
	    RECT 88.6000 125.8000 89.0000 126.2000 ;
	    RECT 91.0000 125.9000 93.5000 126.2000 ;
	    RECT 91.0000 125.8000 91.4000 125.9000 ;
	    RECT 87.1000 125.7000 87.5000 125.8000 ;
	    RECT 85.4000 125.4000 87.5000 125.7000 ;
	    RECT 85.4000 121.1000 85.8000 125.4000 ;
	    RECT 88.7000 125.2000 89.0000 125.8000 ;
	    RECT 91.8000 125.5000 94.6000 125.6000 ;
	    RECT 91.7000 125.4000 94.6000 125.5000 ;
	    RECT 87.8000 124.9000 89.0000 125.2000 ;
	    RECT 89.7000 125.3000 94.6000 125.4000 ;
	    RECT 89.7000 125.1000 92.1000 125.3000 ;
	    RECT 87.8000 124.4000 88.1000 124.9000 ;
	    RECT 87.4000 124.0000 88.1000 124.4000 ;
	    RECT 88.9000 124.5000 89.3000 124.6000 ;
	    RECT 89.7000 124.5000 90.0000 125.1000 ;
	    RECT 88.9000 124.2000 90.0000 124.5000 ;
	    RECT 90.3000 124.5000 93.0000 124.8000 ;
	    RECT 90.3000 124.4000 90.7000 124.5000 ;
	    RECT 92.6000 124.4000 93.0000 124.5000 ;
	    RECT 89.5000 123.7000 89.9000 123.8000 ;
	    RECT 90.9000 123.7000 91.3000 123.8000 ;
	    RECT 87.8000 123.1000 88.2000 123.5000 ;
	    RECT 89.5000 123.4000 91.3000 123.7000 ;
	    RECT 89.9000 123.1000 90.2000 123.4000 ;
	    RECT 92.6000 123.1000 93.0000 123.5000 ;
	    RECT 87.5000 121.1000 88.1000 123.1000 ;
	    RECT 89.8000 121.1000 90.2000 123.1000 ;
	    RECT 92.0000 122.8000 93.0000 123.1000 ;
	    RECT 92.0000 121.1000 92.4000 122.8000 ;
	    RECT 94.2000 121.1000 94.6000 125.3000 ;
	    RECT 95.8000 125.1000 96.2000 126.8000 ;
	    RECT 96.6000 125.1000 97.0000 125.2000 ;
	    RECT 95.8000 124.8000 97.0000 125.1000 ;
	    RECT 95.8000 121.1000 96.2000 124.8000 ;
	    RECT 97.4000 121.1000 97.8000 127.9000 ;
	    RECT 98.2000 124.4000 98.6000 125.2000 ;
	    RECT 99.0000 124.4000 99.4000 125.2000 ;
	    RECT 99.8000 121.1000 100.2000 127.9000 ;
	    RECT 102.2000 127.9000 103.1000 128.2000 ;
	    RECT 100.6000 126.8000 101.0000 127.6000 ;
	    RECT 101.4000 126.8000 101.8000 127.6000 ;
	    RECT 102.2000 121.1000 102.6000 127.9000 ;
	    RECT 103.8000 127.7000 104.2000 129.9000 ;
	    RECT 105.9000 129.2000 106.5000 129.9000 ;
	    RECT 105.9000 128.9000 106.6000 129.2000 ;
	    RECT 108.2000 128.9000 108.6000 129.9000 ;
	    RECT 110.4000 129.2000 110.8000 129.9000 ;
	    RECT 110.4000 128.9000 111.4000 129.2000 ;
	    RECT 106.2000 128.5000 106.6000 128.9000 ;
	    RECT 108.3000 128.6000 108.6000 128.9000 ;
	    RECT 108.3000 128.3000 109.7000 128.6000 ;
	    RECT 109.3000 128.2000 109.7000 128.3000 ;
	    RECT 110.2000 128.2000 110.6000 128.6000 ;
	    RECT 111.0000 128.5000 111.4000 128.9000 ;
	    RECT 105.3000 127.7000 105.7000 127.8000 ;
	    RECT 103.8000 127.4000 105.7000 127.7000 ;
	    RECT 103.8000 125.7000 104.2000 127.4000 ;
	    RECT 107.3000 127.1000 107.7000 127.2000 ;
	    RECT 110.2000 127.1000 110.5000 128.2000 ;
	    RECT 112.6000 127.5000 113.0000 129.9000 ;
	    RECT 116.3000 129.2000 116.7000 129.9000 ;
	    RECT 115.8000 128.8000 116.7000 129.2000 ;
	    RECT 116.3000 128.2000 116.7000 128.8000 ;
	    RECT 115.8000 127.9000 116.7000 128.2000 ;
	    RECT 111.8000 127.1000 112.6000 127.2000 ;
	    RECT 107.1000 126.8000 112.6000 127.1000 ;
	    RECT 115.0000 126.8000 115.4000 127.6000 ;
	    RECT 106.2000 126.4000 106.6000 126.5000 ;
	    RECT 104.7000 126.1000 106.6000 126.4000 ;
	    RECT 104.7000 126.0000 105.1000 126.1000 ;
	    RECT 105.5000 125.7000 105.9000 125.8000 ;
	    RECT 103.8000 125.4000 105.9000 125.7000 ;
	    RECT 103.0000 124.4000 103.4000 125.2000 ;
	    RECT 103.8000 121.1000 104.2000 125.4000 ;
	    RECT 107.1000 125.2000 107.4000 126.8000 ;
	    RECT 110.7000 126.7000 111.1000 126.8000 ;
	    RECT 110.2000 126.2000 110.6000 126.3000 ;
	    RECT 111.5000 126.2000 111.9000 126.3000 ;
	    RECT 109.4000 125.9000 111.9000 126.2000 ;
	    RECT 109.4000 125.8000 109.8000 125.9000 ;
	    RECT 110.2000 125.5000 113.0000 125.6000 ;
	    RECT 110.1000 125.4000 113.0000 125.5000 ;
	    RECT 106.2000 124.9000 107.4000 125.2000 ;
	    RECT 108.1000 125.3000 113.0000 125.4000 ;
	    RECT 108.1000 125.1000 110.5000 125.3000 ;
	    RECT 106.2000 124.4000 106.5000 124.9000 ;
	    RECT 105.8000 124.2000 106.5000 124.4000 ;
	    RECT 107.3000 124.5000 107.7000 124.6000 ;
	    RECT 108.1000 124.5000 108.4000 125.1000 ;
	    RECT 107.3000 124.2000 108.4000 124.5000 ;
	    RECT 108.7000 124.5000 111.4000 124.8000 ;
	    RECT 108.7000 124.4000 109.1000 124.5000 ;
	    RECT 111.0000 124.4000 111.4000 124.5000 ;
	    RECT 105.4000 124.0000 106.5000 124.2000 ;
	    RECT 105.4000 123.8000 106.1000 124.0000 ;
	    RECT 107.9000 123.7000 108.3000 123.8000 ;
	    RECT 109.3000 123.7000 109.7000 123.8000 ;
	    RECT 106.2000 123.1000 106.6000 123.5000 ;
	    RECT 107.9000 123.4000 109.7000 123.7000 ;
	    RECT 108.3000 123.1000 108.6000 123.4000 ;
	    RECT 111.0000 123.1000 111.4000 123.5000 ;
	    RECT 105.9000 121.1000 106.5000 123.1000 ;
	    RECT 108.2000 121.1000 108.6000 123.1000 ;
	    RECT 110.4000 122.8000 111.4000 123.1000 ;
	    RECT 110.4000 121.1000 110.8000 122.8000 ;
	    RECT 112.6000 121.1000 113.0000 125.3000 ;
	    RECT 115.8000 121.1000 116.2000 127.9000 ;
	    RECT 117.4000 127.8000 117.8000 128.6000 ;
	    RECT 116.6000 124.4000 117.0000 125.2000 ;
	    RECT 118.2000 121.1000 118.6000 129.9000 ;
	    RECT 119.3000 128.4000 119.7000 129.9000 ;
	    RECT 119.0000 127.9000 119.7000 128.4000 ;
	    RECT 121.4000 127.9000 121.8000 129.9000 ;
	    RECT 119.0000 126.2000 119.3000 127.9000 ;
	    RECT 121.4000 127.8000 121.7000 127.9000 ;
	    RECT 120.8000 127.6000 121.7000 127.8000 ;
	    RECT 119.6000 127.5000 121.7000 127.6000 ;
	    RECT 119.6000 127.3000 121.1000 127.5000 ;
	    RECT 119.6000 127.2000 120.0000 127.3000 ;
	    RECT 119.0000 125.8000 119.4000 126.2000 ;
	    RECT 119.0000 125.1000 119.3000 125.8000 ;
	    RECT 119.7000 125.5000 120.0000 127.2000 ;
	    RECT 121.4000 127.1000 121.8000 127.2000 ;
	    RECT 122.2000 127.1000 122.6000 129.9000 ;
	    RECT 123.8000 127.6000 124.2000 129.9000 ;
	    RECT 124.6000 127.9000 125.0000 129.9000 ;
	    RECT 125.4000 128.0000 125.8000 129.9000 ;
	    RECT 127.0000 128.0000 127.4000 129.9000 ;
	    RECT 125.4000 127.9000 127.4000 128.0000 ;
	    RECT 129.4000 127.9000 129.8000 129.9000 ;
	    RECT 130.1000 128.2000 130.5000 128.6000 ;
	    RECT 131.1000 128.2000 131.5000 128.6000 ;
	    RECT 120.4000 126.9000 120.8000 127.0000 ;
	    RECT 120.4000 126.6000 120.9000 126.9000 ;
	    RECT 120.6000 126.2000 120.9000 126.6000 ;
	    RECT 121.4000 126.8000 122.6000 127.1000 ;
	    RECT 121.4000 126.4000 121.8000 126.8000 ;
	    RECT 122.2000 126.2000 122.6000 126.8000 ;
	    RECT 123.1000 127.3000 124.2000 127.6000 ;
	    RECT 120.6000 125.8000 121.0000 126.2000 ;
	    RECT 119.7000 125.2000 120.9000 125.5000 ;
	    RECT 119.0000 121.1000 119.4000 125.1000 ;
	    RECT 120.6000 123.1000 120.9000 125.2000 ;
	    RECT 122.2000 125.1000 122.5000 126.2000 ;
	    RECT 123.1000 125.8000 123.4000 127.3000 ;
	    RECT 124.7000 127.2000 125.0000 127.9000 ;
	    RECT 125.5000 127.7000 127.3000 127.9000 ;
	    RECT 126.6000 127.2000 127.0000 127.4000 ;
	    RECT 124.6000 126.8000 125.9000 127.2000 ;
	    RECT 126.6000 127.1000 127.4000 127.2000 ;
	    RECT 128.6000 127.1000 129.0000 127.2000 ;
	    RECT 126.6000 126.9000 129.0000 127.1000 ;
	    RECT 127.0000 126.8000 129.0000 126.9000 ;
	    RECT 122.8000 125.4000 123.4000 125.8000 ;
	    RECT 123.1000 125.1000 123.4000 125.4000 ;
	    RECT 124.6000 125.1000 125.0000 125.2000 ;
	    RECT 125.6000 125.1000 125.9000 126.8000 ;
	    RECT 126.2000 125.8000 126.6000 126.6000 ;
	    RECT 128.6000 126.4000 129.0000 126.8000 ;
	    RECT 127.8000 126.1000 128.2000 126.2000 ;
	    RECT 129.4000 126.1000 129.7000 127.9000 ;
	    RECT 130.2000 127.8000 130.6000 128.2000 ;
	    RECT 131.0000 127.8000 131.4000 128.2000 ;
	    RECT 131.8000 127.9000 132.2000 129.9000 ;
	    RECT 131.0000 126.8000 131.4000 127.2000 ;
	    RECT 131.0000 126.2000 131.3000 126.8000 ;
	    RECT 130.2000 126.1000 130.6000 126.2000 ;
	    RECT 127.8000 125.8000 128.6000 126.1000 ;
	    RECT 129.4000 125.8000 130.6000 126.1000 ;
	    RECT 131.0000 126.1000 131.4000 126.2000 ;
	    RECT 131.9000 126.1000 132.2000 127.9000 ;
	    RECT 135.0000 128.9000 135.4000 129.9000 ;
	    RECT 135.0000 127.2000 135.3000 128.9000 ;
	    RECT 135.8000 127.8000 136.2000 128.6000 ;
	    RECT 132.6000 126.4000 133.0000 127.2000 ;
	    RECT 135.0000 126.8000 135.4000 127.2000 ;
	    RECT 135.8000 126.8000 136.2000 127.2000 ;
	    RECT 133.4000 126.1000 133.8000 126.2000 ;
	    RECT 134.2000 126.1000 134.6000 126.2000 ;
	    RECT 131.0000 125.8000 132.2000 126.1000 ;
	    RECT 133.0000 125.8000 134.6000 126.1000 ;
	    RECT 128.2000 125.6000 128.6000 125.8000 ;
	    RECT 130.2000 125.1000 130.5000 125.8000 ;
	    RECT 131.1000 125.1000 131.4000 125.8000 ;
	    RECT 133.0000 125.6000 133.4000 125.8000 ;
	    RECT 134.2000 125.4000 134.6000 125.8000 ;
	    RECT 135.0000 125.1000 135.3000 126.8000 ;
	    RECT 135.8000 126.1000 136.1000 126.8000 ;
	    RECT 136.6000 126.1000 137.0000 129.9000 ;
	    RECT 137.4000 127.8000 137.8000 128.6000 ;
	    RECT 139.5000 128.2000 139.9000 129.9000 ;
	    RECT 139.0000 127.9000 139.9000 128.2000 ;
	    RECT 142.1000 128.2000 142.9000 129.9000 ;
	    RECT 144.9000 128.2000 145.3000 129.9000 ;
	    RECT 147.1000 128.2000 147.5000 128.6000 ;
	    RECT 142.1000 127.9000 143.4000 128.2000 ;
	    RECT 144.9000 127.9000 145.8000 128.2000 ;
	    RECT 138.2000 126.8000 138.6000 127.6000 ;
	    RECT 135.8000 125.8000 137.0000 126.1000 ;
	    RECT 121.4000 124.1000 121.8000 124.2000 ;
	    RECT 122.2000 124.1000 122.6000 125.1000 ;
	    RECT 123.1000 124.8000 124.2000 125.1000 ;
	    RECT 124.6000 124.8000 125.3000 125.1000 ;
	    RECT 125.6000 124.8000 126.1000 125.1000 ;
	    RECT 121.4000 123.8000 122.6000 124.1000 ;
	    RECT 120.6000 121.1000 121.0000 123.1000 ;
	    RECT 122.2000 121.1000 122.6000 123.8000 ;
	    RECT 123.8000 121.1000 124.2000 124.8000 ;
	    RECT 125.0000 124.2000 125.3000 124.8000 ;
	    RECT 125.0000 123.8000 125.4000 124.2000 ;
	    RECT 125.7000 121.1000 126.1000 124.8000 ;
	    RECT 127.8000 124.8000 129.8000 125.1000 ;
	    RECT 127.8000 121.1000 128.2000 124.8000 ;
	    RECT 129.4000 121.1000 129.8000 124.8000 ;
	    RECT 130.2000 121.1000 130.6000 125.1000 ;
	    RECT 131.0000 121.1000 131.4000 125.1000 ;
	    RECT 131.8000 124.8000 133.8000 125.1000 ;
	    RECT 131.8000 121.1000 132.2000 124.8000 ;
	    RECT 133.4000 121.1000 133.8000 124.8000 ;
	    RECT 134.5000 124.7000 135.4000 125.1000 ;
	    RECT 134.5000 122.2000 134.9000 124.7000 ;
	    RECT 134.5000 121.8000 135.4000 122.2000 ;
	    RECT 134.5000 121.1000 134.9000 121.8000 ;
	    RECT 136.6000 121.1000 137.0000 125.8000 ;
	    RECT 139.0000 121.1000 139.4000 127.9000 ;
	    RECT 142.3000 127.8000 143.4000 127.9000 ;
	    RECT 141.4000 126.4000 141.8000 127.2000 ;
	    RECT 142.3000 126.2000 142.6000 127.8000 ;
	    RECT 143.0000 127.1000 143.4000 127.2000 ;
	    RECT 143.8000 127.1000 144.2000 127.2000 ;
	    RECT 143.0000 126.8000 144.2000 127.1000 ;
	    RECT 143.0000 126.6000 143.3000 126.8000 ;
	    RECT 142.9000 126.2000 143.3000 126.6000 ;
	    RECT 140.6000 126.1000 141.0000 126.2000 ;
	    RECT 139.8000 125.8000 141.4000 126.1000 ;
	    RECT 142.2000 125.8000 142.6000 126.2000 ;
	    RECT 139.8000 125.2000 140.1000 125.8000 ;
	    RECT 141.0000 125.6000 141.4000 125.8000 ;
	    RECT 142.3000 125.7000 142.6000 125.8000 ;
	    RECT 143.8000 126.1000 144.2000 126.2000 ;
	    RECT 145.4000 126.1000 145.8000 127.9000 ;
	    RECT 147.0000 127.8000 147.4000 128.2000 ;
	    RECT 147.8000 127.9000 148.2000 129.9000 ;
	    RECT 151.5000 128.2000 151.9000 129.9000 ;
	    RECT 146.2000 126.8000 146.6000 127.6000 ;
	    RECT 143.8000 125.8000 145.8000 126.1000 ;
	    RECT 147.0000 126.1000 147.4000 126.2000 ;
	    RECT 147.9000 126.1000 148.2000 127.9000 ;
	    RECT 151.0000 127.9000 151.9000 128.2000 ;
	    RECT 154.1000 127.9000 154.9000 129.9000 ;
	    RECT 156.9000 128.2000 157.3000 129.9000 ;
	    RECT 159.3000 129.2000 159.7000 129.9000 ;
	    RECT 159.3000 128.8000 160.2000 129.2000 ;
	    RECT 159.3000 128.2000 159.7000 128.8000 ;
	    RECT 161.7000 128.2000 162.1000 129.9000 ;
	    RECT 156.9000 127.9000 157.8000 128.2000 ;
	    RECT 159.3000 127.9000 160.2000 128.2000 ;
	    RECT 148.6000 126.4000 149.0000 127.2000 ;
	    RECT 150.2000 126.8000 150.6000 127.6000 ;
	    RECT 149.4000 126.1000 149.8000 126.2000 ;
	    RECT 147.0000 125.8000 148.2000 126.1000 ;
	    RECT 149.0000 125.8000 149.8000 126.1000 ;
	    RECT 151.0000 126.1000 151.4000 127.9000 ;
	    RECT 153.4000 126.4000 153.8000 127.2000 ;
	    RECT 154.3000 126.2000 154.6000 127.9000 ;
	    RECT 155.0000 126.8000 155.4000 127.2000 ;
	    RECT 155.0000 126.6000 155.3000 126.8000 ;
	    RECT 154.9000 126.2000 155.3000 126.6000 ;
	    RECT 152.6000 126.1000 153.0000 126.2000 ;
	    RECT 151.0000 125.8000 153.4000 126.1000 ;
	    RECT 154.2000 125.8000 154.6000 126.2000 ;
	    RECT 142.3000 125.4000 143.3000 125.7000 ;
	    RECT 143.8000 125.4000 144.2000 125.8000 ;
	    RECT 139.8000 124.4000 140.2000 125.2000 ;
	    RECT 143.0000 125.1000 143.3000 125.4000 ;
	    RECT 140.6000 124.8000 142.6000 125.1000 ;
	    RECT 140.6000 121.1000 141.0000 124.8000 ;
	    RECT 142.2000 121.4000 142.6000 124.8000 ;
	    RECT 143.0000 121.7000 143.4000 125.1000 ;
	    RECT 143.8000 121.4000 144.2000 125.1000 ;
	    RECT 144.6000 124.4000 145.0000 125.2000 ;
	    RECT 142.2000 121.1000 144.2000 121.4000 ;
	    RECT 145.4000 121.1000 145.8000 125.8000 ;
	    RECT 147.1000 125.1000 147.4000 125.8000 ;
	    RECT 149.0000 125.6000 149.4000 125.8000 ;
	    RECT 147.0000 121.1000 147.4000 125.1000 ;
	    RECT 147.8000 124.8000 149.8000 125.1000 ;
	    RECT 147.8000 121.1000 148.2000 124.8000 ;
	    RECT 149.4000 121.1000 149.8000 124.8000 ;
	    RECT 151.0000 121.1000 151.4000 125.8000 ;
	    RECT 153.0000 125.6000 153.4000 125.8000 ;
	    RECT 154.3000 125.7000 154.6000 125.8000 ;
	    RECT 155.8000 126.1000 156.2000 126.2000 ;
	    RECT 157.4000 126.1000 157.8000 127.9000 ;
	    RECT 158.2000 126.8000 158.6000 127.6000 ;
	    RECT 155.8000 125.8000 157.8000 126.1000 ;
	    RECT 154.3000 125.4000 155.3000 125.7000 ;
	    RECT 155.8000 125.4000 156.2000 125.8000 ;
	    RECT 151.8000 124.4000 152.2000 125.2000 ;
	    RECT 155.0000 125.1000 155.3000 125.4000 ;
	    RECT 152.6000 124.8000 154.6000 125.1000 ;
	    RECT 152.6000 121.1000 153.0000 124.8000 ;
	    RECT 154.2000 121.4000 154.6000 124.8000 ;
	    RECT 155.0000 121.7000 155.4000 125.1000 ;
	    RECT 155.8000 121.4000 156.2000 125.1000 ;
	    RECT 156.6000 124.4000 157.0000 125.2000 ;
	    RECT 154.2000 121.1000 156.2000 121.4000 ;
	    RECT 157.4000 121.1000 157.8000 125.8000 ;
	    RECT 159.0000 124.4000 159.4000 125.2000 ;
	    RECT 159.8000 121.1000 160.2000 127.9000 ;
	    RECT 161.4000 127.8000 162.6000 128.2000 ;
	    RECT 160.6000 126.8000 161.0000 127.6000 ;
	    RECT 161.4000 127.2000 161.7000 127.8000 ;
	    RECT 161.4000 126.8000 161.8000 127.2000 ;
	    RECT 161.4000 124.4000 161.8000 125.2000 ;
	    RECT 162.2000 121.1000 162.6000 127.8000 ;
	    RECT 163.0000 126.8000 163.4000 127.6000 ;
	    RECT 163.8000 127.5000 164.2000 129.9000 ;
	    RECT 166.0000 129.2000 166.4000 129.9000 ;
	    RECT 165.4000 128.9000 166.4000 129.2000 ;
	    RECT 168.2000 128.9000 168.6000 129.9000 ;
	    RECT 170.3000 129.2000 170.9000 129.9000 ;
	    RECT 170.2000 128.9000 170.9000 129.2000 ;
	    RECT 165.4000 128.5000 165.8000 128.9000 ;
	    RECT 168.2000 128.6000 168.5000 128.9000 ;
	    RECT 166.2000 128.2000 166.6000 128.6000 ;
	    RECT 167.1000 128.3000 168.5000 128.6000 ;
	    RECT 170.2000 128.5000 170.6000 128.9000 ;
	    RECT 167.1000 128.2000 167.5000 128.3000 ;
	    RECT 166.3000 127.2000 166.6000 128.2000 ;
	    RECT 171.1000 127.7000 171.5000 127.8000 ;
	    RECT 172.6000 127.7000 173.0000 129.9000 ;
	    RECT 171.1000 127.4000 173.0000 127.7000 ;
	    RECT 164.2000 127.1000 165.0000 127.2000 ;
	    RECT 166.2000 127.1000 166.6000 127.2000 ;
	    RECT 169.1000 127.1000 169.5000 127.2000 ;
	    RECT 164.2000 126.8000 169.7000 127.1000 ;
	    RECT 165.7000 126.7000 166.1000 126.8000 ;
	    RECT 164.9000 126.2000 165.3000 126.3000 ;
	    RECT 164.9000 125.9000 167.4000 126.2000 ;
	    RECT 167.0000 125.8000 167.4000 125.9000 ;
	    RECT 163.8000 125.5000 166.6000 125.6000 ;
	    RECT 163.8000 125.4000 166.7000 125.5000 ;
	    RECT 163.8000 125.3000 168.7000 125.4000 ;
	    RECT 163.8000 121.1000 164.2000 125.3000 ;
	    RECT 166.3000 125.1000 168.7000 125.3000 ;
	    RECT 165.4000 124.5000 168.1000 124.8000 ;
	    RECT 165.4000 124.4000 165.8000 124.5000 ;
	    RECT 167.7000 124.4000 168.1000 124.5000 ;
	    RECT 168.4000 124.5000 168.7000 125.1000 ;
	    RECT 169.4000 125.2000 169.7000 126.8000 ;
	    RECT 170.2000 126.4000 170.6000 126.5000 ;
	    RECT 170.2000 126.1000 172.1000 126.4000 ;
	    RECT 171.7000 126.0000 172.1000 126.1000 ;
	    RECT 170.9000 125.7000 171.3000 125.8000 ;
	    RECT 172.6000 125.7000 173.0000 127.4000 ;
	    RECT 170.9000 125.4000 173.0000 125.7000 ;
	    RECT 169.4000 124.9000 170.6000 125.2000 ;
	    RECT 169.1000 124.5000 169.5000 124.6000 ;
	    RECT 168.4000 124.2000 169.5000 124.5000 ;
	    RECT 170.3000 124.4000 170.6000 124.9000 ;
	    RECT 170.3000 124.0000 171.0000 124.4000 ;
	    RECT 167.1000 123.7000 167.5000 123.8000 ;
	    RECT 168.5000 123.7000 168.9000 123.8000 ;
	    RECT 165.4000 123.1000 165.8000 123.5000 ;
	    RECT 167.1000 123.4000 168.9000 123.7000 ;
	    RECT 168.2000 123.1000 168.5000 123.4000 ;
	    RECT 170.2000 123.1000 170.6000 123.5000 ;
	    RECT 165.4000 122.8000 166.4000 123.1000 ;
	    RECT 166.0000 121.1000 166.4000 122.8000 ;
	    RECT 168.2000 121.1000 168.6000 123.1000 ;
	    RECT 170.3000 121.1000 170.9000 123.1000 ;
	    RECT 172.6000 121.1000 173.0000 125.4000 ;
	    RECT 0.6000 115.6000 1.0000 119.9000 ;
	    RECT 2.7000 116.2000 3.1000 119.9000 ;
	    RECT 2.7000 115.9000 3.4000 116.2000 ;
	    RECT 0.6000 115.4000 2.6000 115.6000 ;
	    RECT 0.6000 115.3000 2.7000 115.4000 ;
	    RECT 2.3000 115.0000 2.7000 115.3000 ;
	    RECT 3.1000 115.2000 3.4000 115.9000 ;
	    RECT 2.4000 113.5000 2.7000 115.0000 ;
	    RECT 3.0000 114.8000 3.4000 115.2000 ;
	    RECT 1.5000 113.2000 2.7000 113.5000 ;
	    RECT 0.6000 112.4000 1.0000 113.2000 ;
	    RECT 1.5000 112.1000 1.8000 113.2000 ;
	    RECT 3.1000 113.1000 3.4000 114.8000 ;
	    RECT 3.8000 113.4000 4.2000 114.2000 ;
	    RECT 1.4000 111.1000 1.8000 112.1000 ;
	    RECT 3.0000 111.1000 3.4000 113.1000 ;
	    RECT 4.6000 113.1000 5.0000 119.9000 ;
	    RECT 5.4000 116.1000 5.8000 116.6000 ;
	    RECT 6.2000 116.1000 6.6000 119.9000 ;
	    RECT 5.4000 115.8000 6.6000 116.1000 ;
	    RECT 4.6000 112.8000 5.5000 113.1000 ;
	    RECT 5.1000 112.2000 5.5000 112.8000 ;
	    RECT 5.1000 111.8000 5.8000 112.2000 ;
	    RECT 5.1000 111.1000 5.5000 111.8000 ;
	    RECT 6.2000 111.1000 6.6000 115.8000 ;
	    RECT 8.6000 116.1000 9.0000 119.9000 ;
	    RECT 10.2000 117.1000 10.6000 119.9000 ;
	    RECT 11.8000 117.9000 12.2000 119.9000 ;
	    RECT 11.9000 117.8000 12.2000 117.9000 ;
	    RECT 13.4000 117.9000 13.8000 119.9000 ;
	    RECT 13.4000 117.8000 13.7000 117.9000 ;
	    RECT 11.9000 117.5000 13.7000 117.8000 ;
	    RECT 10.2000 116.8000 11.3000 117.1000 ;
	    RECT 9.4000 116.1000 9.8000 116.6000 ;
	    RECT 8.6000 115.8000 9.8000 116.1000 ;
	    RECT 8.6000 111.1000 9.0000 115.8000 ;
	    RECT 10.2000 113.1000 10.6000 116.8000 ;
	    RECT 11.0000 116.2000 11.3000 116.8000 ;
	    RECT 11.9000 116.2000 12.2000 117.5000 ;
	    RECT 12.6000 116.4000 13.0000 117.2000 ;
	    RECT 15.3000 116.2000 15.7000 119.9000 ;
	    RECT 11.0000 115.8000 11.4000 116.2000 ;
	    RECT 11.8000 115.8000 12.2000 116.2000 ;
	    RECT 13.4000 116.1000 13.8000 116.2000 ;
	    RECT 14.2000 116.1000 14.6000 116.2000 ;
	    RECT 13.4000 115.8000 14.6000 116.1000 ;
	    RECT 11.9000 114.2000 12.2000 115.8000 ;
	    RECT 14.2000 115.4000 14.6000 115.8000 ;
	    RECT 15.0000 115.9000 15.7000 116.2000 ;
	    RECT 15.0000 115.2000 15.3000 115.9000 ;
	    RECT 17.4000 115.6000 17.8000 119.9000 ;
	    RECT 18.2000 116.2000 18.6000 119.9000 ;
	    RECT 18.2000 115.9000 19.3000 116.2000 ;
	    RECT 19.8000 115.9000 20.2000 119.9000 ;
	    RECT 15.8000 115.4000 17.8000 115.6000 ;
	    RECT 15.7000 115.3000 17.8000 115.4000 ;
	    RECT 19.0000 115.6000 19.3000 115.9000 ;
	    RECT 13.0000 114.8000 13.8000 115.2000 ;
	    RECT 15.0000 114.8000 15.4000 115.2000 ;
	    RECT 15.7000 115.0000 16.1000 115.3000 ;
	    RECT 19.0000 115.2000 19.6000 115.6000 ;
	    RECT 11.0000 113.4000 11.4000 114.2000 ;
	    RECT 11.9000 114.1000 12.7000 114.2000 ;
	    RECT 11.9000 113.9000 12.8000 114.1000 ;
	    RECT 9.7000 112.8000 10.6000 113.1000 ;
	    RECT 9.7000 111.1000 10.1000 112.8000 ;
	    RECT 12.4000 112.2000 12.8000 113.9000 ;
	    RECT 11.8000 111.8000 12.8000 112.2000 ;
	    RECT 12.4000 111.1000 12.8000 111.8000 ;
	    RECT 15.0000 113.1000 15.3000 114.8000 ;
	    RECT 15.7000 113.5000 16.0000 115.0000 ;
	    RECT 19.0000 113.7000 19.3000 115.2000 ;
	    RECT 19.9000 114.8000 20.2000 115.9000 ;
	    RECT 15.7000 113.2000 16.9000 113.5000 ;
	    RECT 18.2000 113.4000 19.3000 113.7000 ;
	    RECT 15.0000 111.1000 15.4000 113.1000 ;
	    RECT 16.6000 112.1000 16.9000 113.2000 ;
	    RECT 17.4000 112.4000 17.8000 113.2000 ;
	    RECT 16.6000 111.1000 17.0000 112.1000 ;
	    RECT 18.2000 111.1000 18.6000 113.4000 ;
	    RECT 19.8000 111.1000 20.2000 114.8000 ;
	    RECT 21.4000 116.1000 21.8000 119.9000 ;
	    RECT 22.2000 116.1000 22.6000 116.6000 ;
	    RECT 21.4000 115.8000 22.6000 116.1000 ;
	    RECT 21.4000 111.1000 21.8000 115.8000 ;
	    RECT 23.0000 113.1000 23.4000 119.9000 ;
	    RECT 24.6000 115.6000 25.0000 119.9000 ;
	    RECT 26.7000 117.1000 27.1000 119.9000 ;
	    RECT 28.6000 117.9000 29.0000 119.9000 ;
	    RECT 28.7000 117.8000 29.0000 117.9000 ;
	    RECT 30.2000 117.9000 30.6000 119.9000 ;
	    RECT 30.2000 117.8000 30.5000 117.9000 ;
	    RECT 28.7000 117.5000 30.5000 117.8000 ;
	    RECT 28.6000 117.1000 29.0000 117.2000 ;
	    RECT 26.7000 116.8000 29.0000 117.1000 ;
	    RECT 26.7000 116.2000 27.1000 116.8000 ;
	    RECT 29.4000 116.4000 29.8000 117.2000 ;
	    RECT 30.2000 116.2000 30.5000 117.5000 ;
	    RECT 26.7000 115.9000 27.4000 116.2000 ;
	    RECT 24.6000 115.4000 26.6000 115.6000 ;
	    RECT 24.6000 115.3000 26.7000 115.4000 ;
	    RECT 26.3000 115.0000 26.7000 115.3000 ;
	    RECT 27.1000 115.2000 27.4000 115.9000 ;
	    RECT 30.2000 115.8000 30.6000 116.2000 ;
	    RECT 23.8000 113.4000 24.2000 114.2000 ;
	    RECT 26.4000 113.5000 26.7000 115.0000 ;
	    RECT 27.0000 114.8000 27.4000 115.2000 ;
	    RECT 28.6000 114.8000 29.4000 115.2000 ;
	    RECT 25.5000 113.2000 26.7000 113.5000 ;
	    RECT 22.5000 112.8000 23.4000 113.1000 ;
	    RECT 22.5000 112.2000 22.9000 112.8000 ;
	    RECT 24.6000 112.4000 25.0000 113.2000 ;
	    RECT 22.5000 111.8000 23.4000 112.2000 ;
	    RECT 25.5000 112.1000 25.8000 113.2000 ;
	    RECT 27.1000 113.1000 27.4000 114.8000 ;
	    RECT 30.2000 114.2000 30.5000 115.8000 ;
	    RECT 29.7000 114.1000 30.5000 114.2000 ;
	    RECT 22.5000 111.1000 22.9000 111.8000 ;
	    RECT 25.4000 111.1000 25.8000 112.1000 ;
	    RECT 27.0000 111.1000 27.4000 113.1000 ;
	    RECT 29.6000 113.9000 30.5000 114.1000 ;
	    RECT 29.6000 112.2000 30.0000 113.9000 ;
	    RECT 29.4000 111.8000 30.0000 112.2000 ;
	    RECT 29.6000 111.1000 30.0000 111.8000 ;
	    RECT 31.8000 111.1000 32.2000 119.9000 ;
	    RECT 33.4000 117.1000 33.8000 119.9000 ;
	    RECT 35.0000 117.9000 35.4000 119.9000 ;
	    RECT 35.1000 117.8000 35.4000 117.9000 ;
	    RECT 36.6000 117.9000 37.0000 119.9000 ;
	    RECT 36.6000 117.8000 36.9000 117.9000 ;
	    RECT 35.1000 117.5000 36.9000 117.8000 ;
	    RECT 34.2000 117.1000 34.6000 117.2000 ;
	    RECT 33.4000 116.8000 34.6000 117.1000 ;
	    RECT 33.4000 111.1000 33.8000 116.8000 ;
	    RECT 35.8000 116.4000 36.2000 117.2000 ;
	    RECT 36.6000 116.2000 36.9000 117.5000 ;
	    RECT 38.2000 117.1000 38.6000 119.9000 ;
	    RECT 38.2000 116.8000 39.3000 117.1000 ;
	    RECT 36.6000 115.8000 37.0000 116.2000 ;
	    RECT 37.4000 115.8000 37.8000 116.6000 ;
	    RECT 35.0000 114.8000 35.8000 115.2000 ;
	    RECT 36.6000 114.2000 36.9000 115.8000 ;
	    RECT 36.1000 114.1000 36.9000 114.2000 ;
	    RECT 36.0000 113.9000 36.9000 114.1000 ;
	    RECT 35.0000 112.1000 35.4000 112.2000 ;
	    RECT 36.0000 112.1000 36.4000 113.9000 ;
	    RECT 38.2000 113.1000 38.6000 116.8000 ;
	    RECT 39.0000 116.2000 39.3000 116.8000 ;
	    RECT 39.8000 116.2000 40.2000 119.9000 ;
	    RECT 39.0000 115.8000 39.4000 116.2000 ;
	    RECT 39.8000 115.9000 40.9000 116.2000 ;
	    RECT 41.4000 115.9000 41.8000 119.9000 ;
	    RECT 40.6000 115.6000 40.9000 115.9000 ;
	    RECT 40.6000 115.2000 41.2000 115.6000 ;
	    RECT 39.0000 113.4000 39.4000 114.2000 ;
	    RECT 40.6000 113.7000 40.9000 115.2000 ;
	    RECT 41.5000 114.8000 41.8000 115.9000 ;
	    RECT 42.2000 115.6000 42.6000 119.9000 ;
	    RECT 44.3000 116.2000 44.7000 119.9000 ;
	    RECT 45.4000 117.9000 45.8000 119.9000 ;
	    RECT 45.5000 117.8000 45.8000 117.9000 ;
	    RECT 47.0000 117.9000 47.4000 119.9000 ;
	    RECT 47.0000 117.8000 47.3000 117.9000 ;
	    RECT 45.5000 117.5000 47.3000 117.8000 ;
	    RECT 45.5000 116.2000 45.8000 117.5000 ;
	    RECT 46.2000 116.4000 46.6000 117.2000 ;
	    RECT 44.3000 115.9000 45.0000 116.2000 ;
	    RECT 42.2000 115.4000 44.2000 115.6000 ;
	    RECT 42.2000 115.3000 44.3000 115.4000 ;
	    RECT 43.9000 115.0000 44.3000 115.3000 ;
	    RECT 44.7000 115.2000 45.0000 115.9000 ;
	    RECT 45.4000 115.8000 45.8000 116.2000 ;
	    RECT 39.8000 113.4000 40.9000 113.7000 ;
	    RECT 35.0000 111.8000 36.4000 112.1000 ;
	    RECT 36.0000 111.1000 36.4000 111.8000 ;
	    RECT 37.7000 112.8000 38.6000 113.1000 ;
	    RECT 37.7000 111.1000 38.1000 112.8000 ;
	    RECT 39.8000 111.1000 40.2000 113.4000 ;
	    RECT 41.4000 113.1000 41.8000 114.8000 ;
	    RECT 44.0000 113.5000 44.3000 115.0000 ;
	    RECT 44.6000 114.8000 45.0000 115.2000 ;
	    RECT 44.7000 114.2000 45.0000 114.8000 ;
	    RECT 44.6000 113.8000 45.0000 114.2000 ;
	    RECT 45.5000 114.2000 45.8000 115.8000 ;
	    RECT 47.8000 115.4000 48.2000 116.2000 ;
	    RECT 48.6000 115.6000 49.0000 119.9000 ;
	    RECT 50.7000 116.2000 51.1000 119.9000 ;
	    RECT 50.7000 115.9000 51.4000 116.2000 ;
	    RECT 48.6000 115.4000 50.6000 115.6000 ;
	    RECT 48.6000 115.3000 50.7000 115.4000 ;
	    RECT 46.6000 114.8000 47.4000 115.2000 ;
	    RECT 50.3000 115.0000 50.7000 115.3000 ;
	    RECT 51.1000 115.2000 51.4000 115.9000 ;
	    RECT 45.5000 114.1000 46.3000 114.2000 ;
	    RECT 45.5000 113.9000 46.4000 114.1000 ;
	    RECT 43.1000 113.2000 44.3000 113.5000 ;
	    RECT 42.2000 113.1000 42.6000 113.2000 ;
	    RECT 41.4000 112.8000 42.6000 113.1000 ;
	    RECT 41.4000 111.1000 41.8000 112.8000 ;
	    RECT 42.2000 112.4000 42.6000 112.8000 ;
	    RECT 43.1000 112.1000 43.4000 113.2000 ;
	    RECT 44.7000 113.1000 45.0000 113.8000 ;
	    RECT 43.0000 111.1000 43.4000 112.1000 ;
	    RECT 44.6000 111.1000 45.0000 113.1000 ;
	    RECT 46.0000 112.1000 46.4000 113.9000 ;
	    RECT 50.4000 113.5000 50.7000 115.0000 ;
	    RECT 51.0000 114.8000 51.4000 115.2000 ;
	    RECT 51.1000 114.2000 51.4000 114.8000 ;
	    RECT 51.0000 113.8000 51.4000 114.2000 ;
	    RECT 49.5000 113.2000 50.7000 113.5000 ;
	    RECT 48.6000 112.4000 49.0000 113.2000 ;
	    RECT 47.0000 112.1000 47.4000 112.2000 ;
	    RECT 49.5000 112.1000 49.8000 113.2000 ;
	    RECT 51.1000 113.1000 51.4000 113.8000 ;
	    RECT 51.8000 113.4000 52.2000 114.2000 ;
	    RECT 46.0000 111.8000 47.4000 112.1000 ;
	    RECT 46.0000 111.1000 46.4000 111.8000 ;
	    RECT 49.4000 111.1000 49.8000 112.1000 ;
	    RECT 51.0000 111.1000 51.4000 113.1000 ;
	    RECT 52.6000 113.1000 53.0000 119.9000 ;
	    RECT 53.4000 116.1000 53.8000 116.6000 ;
	    RECT 54.2000 116.1000 54.6000 119.9000 ;
	    RECT 56.6000 117.9000 57.0000 119.9000 ;
	    RECT 56.7000 117.8000 57.0000 117.9000 ;
	    RECT 58.2000 117.9000 58.6000 119.9000 ;
	    RECT 58.2000 117.8000 58.5000 117.9000 ;
	    RECT 56.7000 117.5000 58.5000 117.8000 ;
	    RECT 57.4000 116.4000 57.8000 117.2000 ;
	    RECT 53.4000 115.8000 54.6000 116.1000 ;
	    RECT 52.6000 112.8000 53.5000 113.1000 ;
	    RECT 53.1000 111.1000 53.5000 112.8000 ;
	    RECT 54.2000 111.1000 54.6000 115.8000 ;
	    RECT 58.2000 116.2000 58.5000 117.5000 ;
	    RECT 58.2000 115.8000 58.6000 116.2000 ;
	    RECT 59.0000 115.9000 59.4000 119.9000 ;
	    RECT 60.6000 116.2000 61.0000 119.9000 ;
	    RECT 59.9000 115.9000 61.0000 116.2000 ;
	    RECT 63.0000 116.2000 63.4000 119.9000 ;
	    RECT 63.0000 115.9000 64.1000 116.2000 ;
	    RECT 64.6000 115.9000 65.0000 119.9000 ;
	    RECT 65.4000 117.9000 65.8000 119.9000 ;
	    RECT 65.5000 117.8000 65.8000 117.9000 ;
	    RECT 67.0000 117.9000 67.4000 119.9000 ;
	    RECT 68.6000 117.9000 69.0000 119.9000 ;
	    RECT 67.0000 117.8000 67.3000 117.9000 ;
	    RECT 65.5000 117.5000 67.3000 117.8000 ;
	    RECT 68.7000 117.8000 69.0000 117.9000 ;
	    RECT 70.2000 117.9000 70.6000 119.9000 ;
	    RECT 70.2000 117.8000 70.5000 117.9000 ;
	    RECT 68.7000 117.5000 70.5000 117.8000 ;
	    RECT 65.5000 116.2000 65.8000 117.5000 ;
	    RECT 66.2000 116.4000 66.6000 117.2000 ;
	    RECT 68.7000 116.2000 69.0000 117.5000 ;
	    RECT 69.4000 116.4000 69.8000 117.2000 ;
	    RECT 56.6000 114.8000 57.4000 115.2000 ;
	    RECT 58.2000 114.2000 58.5000 115.8000 ;
	    RECT 57.7000 114.1000 58.5000 114.2000 ;
	    RECT 57.6000 113.9000 58.5000 114.1000 ;
	    RECT 59.0000 114.8000 59.3000 115.9000 ;
	    RECT 59.9000 115.6000 60.2000 115.9000 ;
	    RECT 59.6000 115.2000 60.2000 115.6000 ;
	    RECT 57.6000 112.2000 58.0000 113.9000 ;
	    RECT 57.4000 111.8000 58.0000 112.2000 ;
	    RECT 57.6000 111.1000 58.0000 111.8000 ;
	    RECT 59.0000 111.1000 59.4000 114.8000 ;
	    RECT 59.9000 113.7000 60.2000 115.2000 ;
	    RECT 63.8000 115.6000 64.1000 115.9000 ;
	    RECT 63.8000 115.2000 64.4000 115.6000 ;
	    RECT 63.8000 113.7000 64.1000 115.2000 ;
	    RECT 64.7000 114.8000 65.0000 115.9000 ;
	    RECT 65.4000 115.8000 65.8000 116.2000 ;
	    RECT 68.6000 115.8000 69.0000 116.2000 ;
	    RECT 59.9000 113.4000 61.0000 113.7000 ;
	    RECT 60.6000 111.1000 61.0000 113.4000 ;
	    RECT 63.0000 113.4000 64.1000 113.7000 ;
	    RECT 63.0000 111.1000 63.4000 113.4000 ;
	    RECT 64.6000 111.1000 65.0000 114.8000 ;
	    RECT 65.5000 114.2000 65.8000 115.8000 ;
	    RECT 66.6000 114.8000 67.4000 115.2000 ;
	    RECT 68.7000 114.2000 69.0000 115.8000 ;
	    RECT 71.8000 115.6000 72.2000 119.9000 ;
	    RECT 73.9000 117.9000 74.5000 119.9000 ;
	    RECT 76.2000 117.9000 76.6000 119.9000 ;
	    RECT 78.4000 118.2000 78.8000 119.9000 ;
	    RECT 78.4000 117.9000 79.4000 118.2000 ;
	    RECT 74.2000 117.5000 74.6000 117.9000 ;
	    RECT 76.3000 117.6000 76.6000 117.9000 ;
	    RECT 75.9000 117.3000 77.7000 117.6000 ;
	    RECT 79.0000 117.5000 79.4000 117.9000 ;
	    RECT 75.9000 117.2000 76.3000 117.3000 ;
	    RECT 77.3000 117.2000 77.7000 117.3000 ;
	    RECT 73.8000 116.6000 74.5000 117.0000 ;
	    RECT 74.2000 116.1000 74.5000 116.6000 ;
	    RECT 75.3000 116.5000 76.4000 116.8000 ;
	    RECT 75.3000 116.4000 75.7000 116.5000 ;
	    RECT 74.2000 115.8000 75.4000 116.1000 ;
	    RECT 71.8000 115.3000 73.9000 115.6000 ;
	    RECT 69.8000 114.8000 70.6000 115.2000 ;
	    RECT 65.5000 114.1000 66.3000 114.2000 ;
	    RECT 68.7000 114.1000 69.5000 114.2000 ;
	    RECT 65.5000 113.9000 66.4000 114.1000 ;
	    RECT 68.7000 113.9000 69.6000 114.1000 ;
	    RECT 66.0000 112.1000 66.4000 113.9000 ;
	    RECT 67.0000 112.1000 67.4000 112.2000 ;
	    RECT 66.0000 111.8000 67.4000 112.1000 ;
	    RECT 69.2000 112.1000 69.6000 113.9000 ;
	    RECT 71.8000 113.6000 72.2000 115.3000 ;
	    RECT 73.5000 115.2000 73.9000 115.3000 ;
	    RECT 72.7000 114.9000 73.1000 115.0000 ;
	    RECT 72.7000 114.6000 74.6000 114.9000 ;
	    RECT 74.2000 114.5000 74.6000 114.6000 ;
	    RECT 75.1000 114.2000 75.4000 115.8000 ;
	    RECT 76.1000 115.9000 76.4000 116.5000 ;
	    RECT 76.7000 116.5000 77.1000 116.6000 ;
	    RECT 79.0000 116.5000 79.4000 116.6000 ;
	    RECT 76.7000 116.2000 79.4000 116.5000 ;
	    RECT 76.1000 115.7000 78.5000 115.9000 ;
	    RECT 80.6000 115.7000 81.0000 119.9000 ;
	    RECT 76.1000 115.6000 81.0000 115.7000 ;
	    RECT 78.1000 115.5000 81.0000 115.6000 ;
	    RECT 78.2000 115.4000 81.0000 115.5000 ;
	    RECT 81.4000 115.7000 81.8000 119.9000 ;
	    RECT 83.6000 118.2000 84.0000 119.9000 ;
	    RECT 83.0000 117.9000 84.0000 118.2000 ;
	    RECT 85.8000 117.9000 86.2000 119.9000 ;
	    RECT 87.9000 117.9000 88.5000 119.9000 ;
	    RECT 83.0000 117.5000 83.4000 117.9000 ;
	    RECT 85.8000 117.6000 86.1000 117.9000 ;
	    RECT 84.7000 117.3000 86.5000 117.6000 ;
	    RECT 87.8000 117.5000 88.2000 117.9000 ;
	    RECT 84.7000 117.2000 85.1000 117.3000 ;
	    RECT 86.1000 117.2000 86.5000 117.3000 ;
	    RECT 88.3000 117.0000 89.0000 117.2000 ;
	    RECT 87.9000 116.8000 89.0000 117.0000 ;
	    RECT 83.0000 116.5000 83.4000 116.6000 ;
	    RECT 85.3000 116.5000 85.7000 116.6000 ;
	    RECT 83.0000 116.2000 85.7000 116.5000 ;
	    RECT 86.0000 116.5000 87.1000 116.8000 ;
	    RECT 86.0000 115.9000 86.3000 116.5000 ;
	    RECT 86.7000 116.4000 87.1000 116.5000 ;
	    RECT 87.9000 116.6000 88.6000 116.8000 ;
	    RECT 87.9000 116.1000 88.2000 116.6000 ;
	    RECT 83.9000 115.7000 86.3000 115.9000 ;
	    RECT 81.4000 115.6000 86.3000 115.7000 ;
	    RECT 87.0000 115.8000 88.2000 116.1000 ;
	    RECT 81.4000 115.5000 84.3000 115.6000 ;
	    RECT 81.4000 115.4000 84.2000 115.5000 ;
	    RECT 87.0000 115.2000 87.3000 115.8000 ;
	    RECT 90.2000 115.6000 90.6000 119.9000 ;
	    RECT 88.5000 115.3000 90.6000 115.6000 ;
	    RECT 88.5000 115.2000 88.9000 115.3000 ;
	    RECT 77.4000 115.1000 77.8000 115.2000 ;
	    RECT 84.6000 115.1000 85.0000 115.2000 ;
	    RECT 77.4000 114.8000 79.9000 115.1000 ;
	    RECT 78.2000 114.7000 78.6000 114.8000 ;
	    RECT 79.5000 114.7000 79.9000 114.8000 ;
	    RECT 82.5000 114.8000 85.0000 115.1000 ;
	    RECT 87.0000 114.8000 87.4000 115.2000 ;
	    RECT 89.3000 114.9000 89.7000 115.0000 ;
	    RECT 82.5000 114.7000 82.9000 114.8000 ;
	    RECT 83.8000 114.7000 84.2000 114.8000 ;
	    RECT 78.7000 114.2000 79.1000 114.3000 ;
	    RECT 83.3000 114.2000 83.7000 114.3000 ;
	    RECT 87.0000 114.2000 87.3000 114.8000 ;
	    RECT 87.8000 114.6000 89.7000 114.9000 ;
	    RECT 87.8000 114.5000 88.2000 114.6000 ;
	    RECT 75.1000 114.1000 80.6000 114.2000 ;
	    RECT 81.8000 114.1000 87.3000 114.2000 ;
	    RECT 75.1000 113.9000 87.3000 114.1000 ;
	    RECT 75.3000 113.8000 75.7000 113.9000 ;
	    RECT 71.8000 113.3000 73.7000 113.6000 ;
	    RECT 70.2000 112.1000 70.6000 112.2000 ;
	    RECT 69.2000 111.8000 70.6000 112.1000 ;
	    RECT 66.0000 111.1000 66.4000 111.8000 ;
	    RECT 69.2000 111.1000 69.6000 111.8000 ;
	    RECT 71.8000 111.1000 72.2000 113.3000 ;
	    RECT 73.3000 113.2000 73.7000 113.3000 ;
	    RECT 78.2000 112.8000 78.5000 113.9000 ;
	    RECT 79.8000 113.8000 82.6000 113.9000 ;
	    RECT 77.3000 112.7000 77.7000 112.8000 ;
	    RECT 74.2000 112.1000 74.6000 112.5000 ;
	    RECT 76.3000 112.4000 77.7000 112.7000 ;
	    RECT 78.2000 112.4000 78.6000 112.8000 ;
	    RECT 76.3000 112.1000 76.6000 112.4000 ;
	    RECT 79.0000 112.1000 79.4000 112.5000 ;
	    RECT 73.9000 111.8000 74.6000 112.1000 ;
	    RECT 73.9000 111.1000 74.5000 111.8000 ;
	    RECT 76.2000 111.1000 76.6000 112.1000 ;
	    RECT 78.4000 111.8000 79.4000 112.1000 ;
	    RECT 78.4000 111.1000 78.8000 111.8000 ;
	    RECT 80.6000 111.1000 81.0000 113.5000 ;
	    RECT 81.4000 111.1000 81.8000 113.5000 ;
	    RECT 83.9000 112.8000 84.2000 113.9000 ;
	    RECT 86.7000 113.8000 87.1000 113.9000 ;
	    RECT 90.2000 113.6000 90.6000 115.3000 ;
	    RECT 88.7000 113.3000 90.6000 113.6000 ;
	    RECT 88.7000 113.2000 89.1000 113.3000 ;
	    RECT 83.0000 112.1000 83.4000 112.5000 ;
	    RECT 83.8000 112.4000 84.2000 112.8000 ;
	    RECT 84.7000 112.7000 85.1000 112.8000 ;
	    RECT 84.7000 112.4000 86.1000 112.7000 ;
	    RECT 85.8000 112.1000 86.1000 112.4000 ;
	    RECT 87.8000 112.1000 88.2000 112.5000 ;
	    RECT 83.0000 111.8000 84.0000 112.1000 ;
	    RECT 83.6000 111.1000 84.0000 111.8000 ;
	    RECT 85.8000 111.1000 86.2000 112.1000 ;
	    RECT 87.8000 111.8000 88.5000 112.1000 ;
	    RECT 87.9000 111.1000 88.5000 111.8000 ;
	    RECT 90.2000 111.1000 90.6000 113.3000 ;
	    RECT 91.0000 115.6000 91.4000 119.9000 ;
	    RECT 93.1000 117.9000 93.7000 119.9000 ;
	    RECT 95.4000 117.9000 95.8000 119.9000 ;
	    RECT 97.6000 118.2000 98.0000 119.9000 ;
	    RECT 97.6000 117.9000 98.6000 118.2000 ;
	    RECT 93.4000 117.5000 93.8000 117.9000 ;
	    RECT 95.5000 117.6000 95.8000 117.9000 ;
	    RECT 95.1000 117.3000 96.9000 117.6000 ;
	    RECT 98.2000 117.5000 98.6000 117.9000 ;
	    RECT 95.1000 117.2000 95.5000 117.3000 ;
	    RECT 96.5000 117.2000 96.9000 117.3000 ;
	    RECT 92.6000 117.0000 93.3000 117.2000 ;
	    RECT 92.6000 116.8000 93.7000 117.0000 ;
	    RECT 93.0000 116.6000 93.7000 116.8000 ;
	    RECT 93.4000 116.1000 93.7000 116.6000 ;
	    RECT 94.5000 116.5000 95.6000 116.8000 ;
	    RECT 94.5000 116.4000 94.9000 116.5000 ;
	    RECT 93.4000 115.8000 94.6000 116.1000 ;
	    RECT 91.0000 115.3000 93.1000 115.6000 ;
	    RECT 91.0000 113.6000 91.4000 115.3000 ;
	    RECT 92.7000 115.2000 93.1000 115.3000 ;
	    RECT 91.9000 114.9000 92.3000 115.0000 ;
	    RECT 91.9000 114.6000 93.8000 114.9000 ;
	    RECT 93.4000 114.5000 93.8000 114.6000 ;
	    RECT 94.3000 114.2000 94.6000 115.8000 ;
	    RECT 95.3000 115.9000 95.6000 116.5000 ;
	    RECT 95.9000 116.5000 96.3000 116.6000 ;
	    RECT 98.2000 116.5000 98.6000 116.6000 ;
	    RECT 95.9000 116.2000 98.6000 116.5000 ;
	    RECT 95.3000 115.7000 97.7000 115.9000 ;
	    RECT 99.8000 115.7000 100.2000 119.9000 ;
	    RECT 95.3000 115.6000 100.2000 115.7000 ;
	    RECT 97.3000 115.5000 100.2000 115.6000 ;
	    RECT 97.4000 115.4000 100.2000 115.5000 ;
	    RECT 100.6000 115.6000 101.0000 119.9000 ;
	    RECT 102.7000 117.9000 103.3000 119.9000 ;
	    RECT 105.0000 117.9000 105.4000 119.9000 ;
	    RECT 107.2000 118.2000 107.6000 119.9000 ;
	    RECT 107.2000 117.9000 108.2000 118.2000 ;
	    RECT 103.0000 117.5000 103.4000 117.9000 ;
	    RECT 105.1000 117.6000 105.4000 117.9000 ;
	    RECT 104.7000 117.3000 106.5000 117.6000 ;
	    RECT 107.8000 117.5000 108.2000 117.9000 ;
	    RECT 104.7000 117.2000 105.1000 117.3000 ;
	    RECT 106.1000 117.2000 106.5000 117.3000 ;
	    RECT 102.6000 116.6000 103.3000 117.0000 ;
	    RECT 103.0000 116.1000 103.3000 116.6000 ;
	    RECT 104.1000 116.5000 105.2000 116.8000 ;
	    RECT 104.1000 116.4000 104.5000 116.5000 ;
	    RECT 103.0000 115.8000 104.2000 116.1000 ;
	    RECT 100.6000 115.3000 102.7000 115.6000 ;
	    RECT 96.6000 115.1000 97.0000 115.2000 ;
	    RECT 96.6000 114.8000 99.1000 115.1000 ;
	    RECT 97.4000 114.7000 97.8000 114.8000 ;
	    RECT 98.7000 114.7000 99.1000 114.8000 ;
	    RECT 97.9000 114.2000 98.3000 114.3000 ;
	    RECT 94.3000 113.9000 99.8000 114.2000 ;
	    RECT 94.5000 113.8000 94.9000 113.9000 ;
	    RECT 91.0000 113.3000 92.9000 113.6000 ;
	    RECT 91.0000 111.1000 91.4000 113.3000 ;
	    RECT 92.5000 113.2000 92.9000 113.3000 ;
	    RECT 97.4000 112.8000 97.7000 113.9000 ;
	    RECT 99.0000 113.8000 99.8000 113.9000 ;
	    RECT 100.6000 113.6000 101.0000 115.3000 ;
	    RECT 102.3000 115.2000 102.7000 115.3000 ;
	    RECT 101.5000 114.9000 101.9000 115.0000 ;
	    RECT 101.5000 114.6000 103.4000 114.9000 ;
	    RECT 103.0000 114.5000 103.4000 114.6000 ;
	    RECT 103.9000 114.2000 104.2000 115.8000 ;
	    RECT 104.9000 115.9000 105.2000 116.5000 ;
	    RECT 105.5000 116.5000 105.9000 116.6000 ;
	    RECT 107.8000 116.5000 108.2000 116.6000 ;
	    RECT 105.5000 116.2000 108.2000 116.5000 ;
	    RECT 104.9000 115.7000 107.3000 115.9000 ;
	    RECT 109.4000 115.7000 109.8000 119.9000 ;
	    RECT 104.9000 115.6000 109.8000 115.7000 ;
	    RECT 106.9000 115.5000 109.8000 115.6000 ;
	    RECT 107.0000 115.4000 109.8000 115.5000 ;
	    RECT 111.8000 115.7000 112.2000 119.9000 ;
	    RECT 114.0000 118.2000 114.4000 119.9000 ;
	    RECT 113.4000 117.9000 114.4000 118.2000 ;
	    RECT 116.2000 117.9000 116.6000 119.9000 ;
	    RECT 118.3000 117.9000 118.9000 119.9000 ;
	    RECT 113.4000 117.5000 113.8000 117.9000 ;
	    RECT 116.2000 117.6000 116.5000 117.9000 ;
	    RECT 115.1000 117.3000 116.9000 117.6000 ;
	    RECT 118.2000 117.5000 118.6000 117.9000 ;
	    RECT 115.1000 117.2000 115.5000 117.3000 ;
	    RECT 116.5000 117.2000 116.9000 117.3000 ;
	    RECT 113.4000 116.5000 113.8000 116.6000 ;
	    RECT 115.7000 116.5000 116.1000 116.6000 ;
	    RECT 113.4000 116.2000 116.1000 116.5000 ;
	    RECT 116.4000 116.5000 117.5000 116.8000 ;
	    RECT 116.4000 115.9000 116.7000 116.5000 ;
	    RECT 117.1000 116.4000 117.5000 116.5000 ;
	    RECT 118.3000 116.6000 119.0000 117.0000 ;
	    RECT 118.3000 116.1000 118.6000 116.6000 ;
	    RECT 114.3000 115.7000 116.7000 115.9000 ;
	    RECT 111.8000 115.6000 116.7000 115.7000 ;
	    RECT 117.4000 115.8000 118.6000 116.1000 ;
	    RECT 111.8000 115.5000 114.7000 115.6000 ;
	    RECT 111.8000 115.4000 114.6000 115.5000 ;
	    RECT 106.2000 115.1000 106.6000 115.2000 ;
	    RECT 115.0000 115.1000 115.4000 115.2000 ;
	    RECT 115.8000 115.1000 116.2000 115.2000 ;
	    RECT 106.2000 114.8000 108.7000 115.1000 ;
	    RECT 107.0000 114.7000 107.4000 114.8000 ;
	    RECT 108.3000 114.7000 108.7000 114.8000 ;
	    RECT 112.9000 114.8000 116.2000 115.1000 ;
	    RECT 112.9000 114.7000 113.3000 114.8000 ;
	    RECT 107.5000 114.2000 107.9000 114.3000 ;
	    RECT 113.7000 114.2000 114.1000 114.3000 ;
	    RECT 117.4000 114.2000 117.7000 115.8000 ;
	    RECT 120.6000 115.6000 121.0000 119.9000 ;
	    RECT 121.8000 116.8000 122.2000 117.2000 ;
	    RECT 121.8000 116.2000 122.1000 116.8000 ;
	    RECT 122.5000 116.2000 122.9000 119.9000 ;
	    RECT 121.4000 115.9000 122.1000 116.2000 ;
	    RECT 122.4000 115.9000 122.9000 116.2000 ;
	    RECT 124.9000 116.3000 125.3000 119.9000 ;
	    RECT 127.8000 117.9000 128.2000 119.9000 ;
	    RECT 124.9000 115.9000 125.8000 116.3000 ;
	    RECT 121.4000 115.8000 121.8000 115.9000 ;
	    RECT 118.9000 115.3000 121.0000 115.6000 ;
	    RECT 118.9000 115.2000 119.3000 115.3000 ;
	    RECT 119.7000 114.9000 120.1000 115.0000 ;
	    RECT 118.2000 114.6000 120.1000 114.9000 ;
	    RECT 118.2000 114.5000 118.6000 114.6000 ;
	    RECT 103.9000 114.1000 109.4000 114.2000 ;
	    RECT 112.2000 114.1000 117.7000 114.2000 ;
	    RECT 103.9000 113.9000 117.7000 114.1000 ;
	    RECT 104.1000 113.8000 104.5000 113.9000 ;
	    RECT 96.5000 112.7000 96.9000 112.8000 ;
	    RECT 93.4000 112.1000 93.8000 112.5000 ;
	    RECT 95.5000 112.4000 96.9000 112.7000 ;
	    RECT 97.4000 112.4000 97.8000 112.8000 ;
	    RECT 95.5000 112.1000 95.8000 112.4000 ;
	    RECT 98.2000 112.1000 98.6000 112.5000 ;
	    RECT 93.1000 111.8000 93.8000 112.1000 ;
	    RECT 93.1000 111.1000 93.7000 111.8000 ;
	    RECT 95.4000 111.1000 95.8000 112.1000 ;
	    RECT 97.6000 111.8000 98.6000 112.1000 ;
	    RECT 97.6000 111.1000 98.0000 111.8000 ;
	    RECT 99.8000 111.1000 100.2000 113.5000 ;
	    RECT 100.6000 113.3000 102.5000 113.6000 ;
	    RECT 100.6000 111.1000 101.0000 113.3000 ;
	    RECT 102.1000 113.2000 102.5000 113.3000 ;
	    RECT 107.0000 112.8000 107.3000 113.9000 ;
	    RECT 108.6000 113.8000 113.0000 113.9000 ;
	    RECT 106.1000 112.7000 106.5000 112.8000 ;
	    RECT 103.0000 112.1000 103.4000 112.5000 ;
	    RECT 105.1000 112.4000 106.5000 112.7000 ;
	    RECT 107.0000 112.4000 107.4000 112.8000 ;
	    RECT 105.1000 112.1000 105.4000 112.4000 ;
	    RECT 107.8000 112.1000 108.2000 112.5000 ;
	    RECT 102.7000 111.8000 103.4000 112.1000 ;
	    RECT 102.7000 111.1000 103.3000 111.8000 ;
	    RECT 105.0000 111.1000 105.4000 112.1000 ;
	    RECT 107.2000 111.8000 108.2000 112.1000 ;
	    RECT 107.2000 111.1000 107.6000 111.8000 ;
	    RECT 109.4000 111.1000 109.8000 113.5000 ;
	    RECT 111.8000 111.1000 112.2000 113.5000 ;
	    RECT 114.3000 113.2000 114.6000 113.9000 ;
	    RECT 117.1000 113.8000 117.5000 113.9000 ;
	    RECT 120.6000 113.6000 121.0000 115.3000 ;
	    RECT 122.4000 115.2000 122.7000 115.9000 ;
	    RECT 122.2000 114.8000 122.7000 115.2000 ;
	    RECT 122.4000 114.2000 122.7000 114.8000 ;
	    RECT 123.0000 115.1000 123.4000 115.2000 ;
	    RECT 123.8000 115.1000 124.2000 115.2000 ;
	    RECT 123.0000 114.8000 124.2000 115.1000 ;
	    RECT 124.6000 114.8000 125.0000 115.6000 ;
	    RECT 123.0000 114.4000 123.4000 114.8000 ;
	    RECT 125.4000 114.2000 125.7000 115.9000 ;
	    RECT 127.9000 115.8000 128.2000 117.9000 ;
	    RECT 129.4000 115.9000 129.8000 119.9000 ;
	    RECT 130.5000 116.3000 130.9000 119.9000 ;
	    RECT 130.5000 115.9000 131.4000 116.3000 ;
	    RECT 133.9000 116.2000 134.3000 119.9000 ;
	    RECT 134.6000 116.8000 135.0000 117.2000 ;
	    RECT 134.7000 116.2000 135.0000 116.8000 ;
	    RECT 133.9000 115.9000 134.4000 116.2000 ;
	    RECT 134.7000 115.9000 135.4000 116.2000 ;
	    RECT 127.9000 115.5000 129.1000 115.8000 ;
	    RECT 127.8000 114.8000 128.2000 115.2000 ;
	    RECT 121.4000 113.8000 122.7000 114.2000 ;
	    RECT 123.8000 114.1000 124.2000 114.2000 ;
	    RECT 123.4000 113.8000 124.2000 114.1000 ;
	    RECT 125.4000 113.8000 125.8000 114.2000 ;
	    RECT 127.0000 113.8000 127.4000 114.6000 ;
	    RECT 127.9000 114.4000 128.2000 114.8000 ;
	    RECT 127.9000 114.1000 128.4000 114.4000 ;
	    RECT 128.0000 114.0000 128.4000 114.1000 ;
	    RECT 128.8000 113.8000 129.1000 115.5000 ;
	    RECT 129.5000 115.2000 129.8000 115.9000 ;
	    RECT 129.4000 114.8000 129.8000 115.2000 ;
	    RECT 130.2000 114.8000 130.6000 115.6000 ;
	    RECT 119.1000 113.3000 121.0000 113.6000 ;
	    RECT 119.1000 113.2000 119.5000 113.3000 ;
	    RECT 113.4000 112.1000 113.8000 112.5000 ;
	    RECT 114.2000 112.4000 114.6000 113.2000 ;
	    RECT 115.1000 112.7000 115.5000 112.8000 ;
	    RECT 115.1000 112.4000 116.5000 112.7000 ;
	    RECT 116.2000 112.1000 116.5000 112.4000 ;
	    RECT 118.2000 112.1000 118.6000 112.5000 ;
	    RECT 113.4000 111.8000 114.4000 112.1000 ;
	    RECT 114.0000 111.1000 114.4000 111.8000 ;
	    RECT 116.2000 111.1000 116.6000 112.1000 ;
	    RECT 118.2000 111.8000 118.9000 112.1000 ;
	    RECT 118.3000 111.1000 118.9000 111.8000 ;
	    RECT 120.6000 111.1000 121.0000 113.3000 ;
	    RECT 121.5000 113.1000 121.8000 113.8000 ;
	    RECT 123.4000 113.6000 123.8000 113.8000 ;
	    RECT 122.3000 113.1000 124.1000 113.3000 ;
	    RECT 121.4000 111.1000 121.8000 113.1000 ;
	    RECT 122.2000 113.0000 124.2000 113.1000 ;
	    RECT 122.2000 111.1000 122.6000 113.0000 ;
	    RECT 123.8000 111.1000 124.2000 113.0000 ;
	    RECT 125.4000 112.2000 125.7000 113.8000 ;
	    RECT 128.8000 113.7000 129.2000 113.8000 ;
	    RECT 127.7000 113.5000 129.2000 113.7000 ;
	    RECT 127.1000 113.4000 129.2000 113.5000 ;
	    RECT 127.1000 113.2000 128.0000 113.4000 ;
	    RECT 126.2000 112.4000 126.6000 113.2000 ;
	    RECT 127.1000 113.1000 127.4000 113.2000 ;
	    RECT 129.5000 113.1000 129.8000 114.8000 ;
	    RECT 125.4000 111.1000 125.8000 112.2000 ;
	    RECT 127.0000 111.1000 127.4000 113.1000 ;
	    RECT 129.1000 112.6000 129.8000 113.1000 ;
	    RECT 131.0000 114.2000 131.3000 115.9000 ;
	    RECT 133.4000 114.4000 133.8000 115.2000 ;
	    RECT 134.1000 115.1000 134.4000 115.9000 ;
	    RECT 135.0000 115.8000 135.4000 115.9000 ;
	    RECT 135.8000 115.8000 136.2000 116.6000 ;
	    RECT 135.0000 115.1000 135.4000 115.2000 ;
	    RECT 134.1000 114.8000 135.4000 115.1000 ;
	    RECT 134.1000 114.2000 134.4000 114.8000 ;
	    RECT 131.0000 114.1000 131.4000 114.2000 ;
	    RECT 132.6000 114.1000 133.0000 114.2000 ;
	    RECT 131.0000 113.8000 133.4000 114.1000 ;
	    RECT 134.1000 113.8000 135.4000 114.2000 ;
	    RECT 129.1000 112.2000 129.5000 112.6000 ;
	    RECT 129.1000 111.8000 129.8000 112.2000 ;
	    RECT 131.0000 112.1000 131.3000 113.8000 ;
	    RECT 133.0000 113.6000 133.4000 113.8000 ;
	    RECT 131.8000 112.4000 132.2000 113.2000 ;
	    RECT 132.7000 113.1000 134.5000 113.3000 ;
	    RECT 135.0000 113.1000 135.3000 113.8000 ;
	    RECT 136.6000 113.1000 137.0000 119.9000 ;
	    RECT 139.5000 116.2000 139.9000 119.9000 ;
	    RECT 142.2000 117.9000 142.6000 119.9000 ;
	    RECT 140.2000 116.8000 140.6000 117.2000 ;
	    RECT 140.3000 116.2000 140.6000 116.8000 ;
	    RECT 139.5000 115.9000 140.0000 116.2000 ;
	    RECT 140.3000 115.9000 141.0000 116.2000 ;
	    RECT 137.4000 115.1000 137.8000 115.2000 ;
	    RECT 139.0000 115.1000 139.4000 115.2000 ;
	    RECT 137.4000 114.8000 139.4000 115.1000 ;
	    RECT 139.0000 114.4000 139.4000 114.8000 ;
	    RECT 139.7000 114.2000 140.0000 115.9000 ;
	    RECT 140.6000 115.8000 141.0000 115.9000 ;
	    RECT 142.3000 115.8000 142.6000 117.9000 ;
	    RECT 143.8000 115.9000 144.2000 119.9000 ;
	    RECT 145.9000 119.2000 146.3000 119.9000 ;
	    RECT 145.4000 118.8000 146.3000 119.2000 ;
	    RECT 145.9000 116.2000 146.3000 118.8000 ;
	    RECT 146.6000 116.8000 147.0000 117.2000 ;
	    RECT 146.7000 116.2000 147.0000 116.8000 ;
	    RECT 148.2000 116.8000 148.6000 117.2000 ;
	    RECT 148.2000 116.2000 148.5000 116.8000 ;
	    RECT 148.9000 116.2000 149.3000 119.9000 ;
	    RECT 145.9000 115.9000 146.4000 116.2000 ;
	    RECT 146.7000 115.9000 147.4000 116.2000 ;
	    RECT 142.3000 115.5000 143.5000 115.8000 ;
	    RECT 142.2000 114.8000 142.6000 115.2000 ;
	    RECT 137.4000 114.1000 137.8000 114.2000 ;
	    RECT 138.2000 114.1000 138.6000 114.2000 ;
	    RECT 137.4000 113.8000 139.0000 114.1000 ;
	    RECT 139.7000 113.8000 141.0000 114.2000 ;
	    RECT 141.4000 113.8000 141.8000 114.6000 ;
	    RECT 142.3000 114.4000 142.6000 114.8000 ;
	    RECT 142.2000 114.0000 142.8000 114.4000 ;
	    RECT 143.2000 113.8000 143.5000 115.5000 ;
	    RECT 143.9000 115.2000 144.2000 115.9000 ;
	    RECT 143.8000 114.8000 144.2000 115.2000 ;
	    RECT 144.6000 115.1000 145.0000 115.2000 ;
	    RECT 145.4000 115.1000 145.8000 115.2000 ;
	    RECT 144.6000 114.8000 145.8000 115.1000 ;
	    RECT 137.4000 113.4000 137.8000 113.8000 ;
	    RECT 138.6000 113.6000 139.0000 113.8000 ;
	    RECT 138.3000 113.1000 140.1000 113.3000 ;
	    RECT 140.6000 113.1000 140.9000 113.8000 ;
	    RECT 143.2000 113.7000 143.6000 113.8000 ;
	    RECT 142.1000 113.5000 143.6000 113.7000 ;
	    RECT 141.5000 113.4000 143.6000 113.5000 ;
	    RECT 141.5000 113.2000 142.4000 113.4000 ;
	    RECT 141.5000 113.1000 141.8000 113.2000 ;
	    RECT 143.9000 113.1000 144.2000 114.8000 ;
	    RECT 145.4000 114.4000 145.8000 114.8000 ;
	    RECT 146.1000 114.2000 146.4000 115.9000 ;
	    RECT 147.0000 115.8000 147.4000 115.9000 ;
	    RECT 147.8000 115.9000 148.5000 116.2000 ;
	    RECT 148.8000 115.9000 149.3000 116.2000 ;
	    RECT 147.8000 115.8000 148.2000 115.9000 ;
	    RECT 147.0000 115.1000 147.4000 115.2000 ;
	    RECT 148.8000 115.1000 149.1000 115.9000 ;
	    RECT 151.0000 115.8000 151.4000 116.6000 ;
	    RECT 147.0000 114.8000 149.1000 115.1000 ;
	    RECT 148.8000 114.2000 149.1000 114.8000 ;
	    RECT 149.4000 114.4000 149.8000 115.2000 ;
	    RECT 144.6000 114.1000 145.0000 114.2000 ;
	    RECT 144.6000 113.8000 145.4000 114.1000 ;
	    RECT 146.1000 113.8000 147.4000 114.2000 ;
	    RECT 147.8000 113.8000 149.1000 114.2000 ;
	    RECT 150.2000 114.1000 150.6000 114.2000 ;
	    RECT 149.8000 113.8000 150.6000 114.1000 ;
	    RECT 145.0000 113.6000 145.4000 113.8000 ;
	    RECT 144.7000 113.1000 146.5000 113.3000 ;
	    RECT 147.0000 113.1000 147.3000 113.8000 ;
	    RECT 147.9000 113.1000 148.2000 113.8000 ;
	    RECT 149.8000 113.6000 150.2000 113.8000 ;
	    RECT 148.7000 113.1000 150.5000 113.3000 ;
	    RECT 151.8000 113.1000 152.2000 119.9000 ;
	    RECT 153.4000 117.1000 153.8000 119.9000 ;
	    RECT 152.6000 116.8000 153.8000 117.1000 ;
	    RECT 152.6000 116.2000 152.9000 116.8000 ;
	    RECT 152.6000 115.8000 153.0000 116.2000 ;
	    RECT 152.6000 113.4000 153.0000 114.2000 ;
	    RECT 132.6000 113.0000 134.6000 113.1000 ;
	    RECT 129.1000 111.1000 129.5000 111.8000 ;
	    RECT 131.0000 111.1000 131.4000 112.1000 ;
	    RECT 132.6000 111.1000 133.0000 113.0000 ;
	    RECT 134.2000 111.1000 134.6000 113.0000 ;
	    RECT 135.0000 111.1000 135.4000 113.1000 ;
	    RECT 136.1000 112.8000 137.0000 113.1000 ;
	    RECT 138.2000 113.0000 140.2000 113.1000 ;
	    RECT 136.1000 112.2000 136.5000 112.8000 ;
	    RECT 135.8000 111.8000 136.5000 112.2000 ;
	    RECT 136.1000 111.1000 136.5000 111.8000 ;
	    RECT 138.2000 111.1000 138.6000 113.0000 ;
	    RECT 139.8000 111.1000 140.2000 113.0000 ;
	    RECT 140.6000 111.1000 141.0000 113.1000 ;
	    RECT 141.4000 111.1000 141.8000 113.1000 ;
	    RECT 143.5000 112.6000 144.2000 113.1000 ;
	    RECT 144.6000 113.0000 146.6000 113.1000 ;
	    RECT 143.5000 111.1000 143.9000 112.6000 ;
	    RECT 144.6000 111.1000 145.0000 113.0000 ;
	    RECT 146.2000 111.1000 146.6000 113.0000 ;
	    RECT 147.0000 111.1000 147.4000 113.1000 ;
	    RECT 147.8000 111.1000 148.2000 113.1000 ;
	    RECT 148.6000 113.0000 150.6000 113.1000 ;
	    RECT 148.6000 111.1000 149.0000 113.0000 ;
	    RECT 150.2000 111.1000 150.6000 113.0000 ;
	    RECT 151.3000 112.8000 152.2000 113.1000 ;
	    RECT 151.3000 112.2000 151.7000 112.8000 ;
	    RECT 151.0000 111.8000 151.7000 112.2000 ;
	    RECT 151.3000 111.1000 151.7000 111.8000 ;
	    RECT 153.4000 111.1000 153.8000 116.8000 ;
	    RECT 154.2000 114.8000 154.6000 115.2000 ;
	    RECT 154.2000 114.2000 154.5000 114.8000 ;
	    RECT 154.2000 113.4000 154.6000 114.2000 ;
	    RECT 155.0000 113.4000 155.4000 114.2000 ;
	    RECT 155.8000 113.1000 156.2000 119.9000 ;
	    RECT 156.6000 115.8000 157.0000 116.6000 ;
	    RECT 157.4000 113.4000 157.8000 114.2000 ;
	    RECT 158.2000 114.1000 158.6000 119.9000 ;
	    RECT 160.3000 115.9000 161.3000 119.9000 ;
	    RECT 160.6000 115.2000 160.9000 115.9000 ;
	    RECT 163.0000 115.7000 163.4000 119.9000 ;
	    RECT 165.2000 118.2000 165.6000 119.9000 ;
	    RECT 164.6000 117.9000 165.6000 118.2000 ;
	    RECT 167.4000 117.9000 167.8000 119.9000 ;
	    RECT 169.5000 117.9000 170.1000 119.9000 ;
	    RECT 164.6000 117.5000 165.0000 117.9000 ;
	    RECT 167.4000 117.6000 167.7000 117.9000 ;
	    RECT 166.3000 117.3000 168.1000 117.6000 ;
	    RECT 169.4000 117.5000 169.8000 117.9000 ;
	    RECT 166.3000 117.2000 166.7000 117.3000 ;
	    RECT 167.7000 117.2000 168.1000 117.3000 ;
	    RECT 164.6000 116.5000 165.0000 116.6000 ;
	    RECT 166.9000 116.5000 167.3000 116.6000 ;
	    RECT 164.6000 116.2000 167.3000 116.5000 ;
	    RECT 167.6000 116.5000 168.7000 116.8000 ;
	    RECT 167.6000 115.9000 167.9000 116.5000 ;
	    RECT 168.3000 116.4000 168.7000 116.5000 ;
	    RECT 169.5000 116.6000 170.2000 117.0000 ;
	    RECT 169.5000 116.1000 169.8000 116.6000 ;
	    RECT 165.5000 115.7000 167.9000 115.9000 ;
	    RECT 163.0000 115.6000 167.9000 115.7000 ;
	    RECT 168.6000 115.8000 169.8000 116.1000 ;
	    RECT 163.0000 115.5000 165.9000 115.6000 ;
	    RECT 163.0000 115.4000 165.8000 115.5000 ;
	    RECT 159.8000 114.4000 160.2000 115.2000 ;
	    RECT 160.6000 114.8000 161.0000 115.2000 ;
	    RECT 160.6000 114.2000 160.9000 114.8000 ;
	    RECT 161.4000 114.4000 161.8000 115.2000 ;
	    RECT 166.2000 115.1000 166.6000 115.2000 ;
	    RECT 167.0000 115.1000 167.4000 115.2000 ;
	    RECT 164.1000 114.8000 167.4000 115.1000 ;
	    RECT 164.1000 114.7000 164.5000 114.8000 ;
	    RECT 159.0000 114.1000 159.4000 114.2000 ;
	    RECT 160.6000 114.1000 161.0000 114.2000 ;
	    RECT 158.2000 113.8000 159.8000 114.1000 ;
	    RECT 160.6000 113.8000 161.8000 114.1000 ;
	    RECT 162.2000 113.8000 162.6000 114.6000 ;
	    RECT 164.9000 114.2000 165.3000 114.3000 ;
	    RECT 168.6000 114.2000 168.9000 115.8000 ;
	    RECT 171.8000 115.6000 172.2000 119.9000 ;
	    RECT 170.1000 115.3000 172.2000 115.6000 ;
	    RECT 170.1000 115.2000 170.5000 115.3000 ;
	    RECT 170.9000 114.9000 171.3000 115.0000 ;
	    RECT 169.4000 114.6000 171.3000 114.9000 ;
	    RECT 169.4000 114.5000 169.8000 114.6000 ;
	    RECT 163.4000 113.9000 168.9000 114.2000 ;
	    RECT 163.4000 113.8000 164.2000 113.9000 ;
	    RECT 155.8000 112.8000 156.7000 113.1000 ;
	    RECT 156.3000 111.1000 156.7000 112.8000 ;
	    RECT 158.2000 111.1000 158.6000 113.8000 ;
	    RECT 159.4000 113.6000 159.8000 113.8000 ;
	    RECT 159.1000 113.1000 160.9000 113.3000 ;
	    RECT 161.5000 113.1000 161.8000 113.8000 ;
	    RECT 159.0000 113.0000 161.0000 113.1000 ;
	    RECT 159.0000 111.1000 159.4000 113.0000 ;
	    RECT 160.6000 111.4000 161.0000 113.0000 ;
	    RECT 161.4000 111.7000 161.8000 113.1000 ;
	    RECT 162.2000 111.4000 162.6000 113.1000 ;
	    RECT 160.6000 111.1000 162.6000 111.4000 ;
	    RECT 163.0000 111.1000 163.4000 113.5000 ;
	    RECT 165.5000 113.2000 165.8000 113.9000 ;
	    RECT 166.2000 113.8000 166.6000 113.9000 ;
	    RECT 168.3000 113.8000 168.7000 113.9000 ;
	    RECT 171.8000 113.6000 172.2000 115.3000 ;
	    RECT 170.3000 113.3000 172.2000 113.6000 ;
	    RECT 170.3000 113.2000 170.7000 113.3000 ;
	    RECT 164.6000 112.1000 165.0000 112.5000 ;
	    RECT 165.4000 112.4000 165.8000 113.2000 ;
	    RECT 166.3000 112.7000 166.7000 112.8000 ;
	    RECT 166.3000 112.4000 167.7000 112.7000 ;
	    RECT 167.4000 112.1000 167.7000 112.4000 ;
	    RECT 169.4000 112.1000 169.8000 112.5000 ;
	    RECT 164.6000 111.8000 165.6000 112.1000 ;
	    RECT 165.2000 111.1000 165.6000 111.8000 ;
	    RECT 167.4000 111.1000 167.8000 112.1000 ;
	    RECT 169.4000 111.8000 170.1000 112.1000 ;
	    RECT 169.5000 111.1000 170.1000 111.8000 ;
	    RECT 171.8000 111.1000 172.2000 113.3000 ;
	    RECT 0.6000 105.1000 1.0000 105.2000 ;
	    RECT 1.4000 105.1000 1.8000 109.9000 ;
	    RECT 4.0000 107.1000 4.4000 109.9000 ;
	    RECT 5.7000 108.2000 6.1000 109.9000 ;
	    RECT 5.7000 107.9000 6.6000 108.2000 ;
	    RECT 4.0000 106.9000 4.9000 107.1000 ;
	    RECT 4.1000 106.8000 4.9000 106.9000 ;
	    RECT 3.0000 105.8000 3.8000 106.2000 ;
	    RECT 0.6000 104.8000 1.8000 105.1000 ;
	    RECT 2.2000 105.1000 2.6000 105.6000 ;
	    RECT 4.6000 105.2000 4.9000 106.8000 ;
	    RECT 3.0000 105.1000 3.4000 105.2000 ;
	    RECT 2.2000 104.8000 3.4000 105.1000 ;
	    RECT 4.6000 104.8000 5.0000 105.2000 ;
	    RECT 1.4000 101.1000 1.8000 104.8000 ;
	    RECT 3.8000 103.8000 4.2000 104.6000 ;
	    RECT 4.6000 103.5000 4.9000 104.8000 ;
	    RECT 5.4000 104.4000 5.8000 105.2000 ;
	    RECT 3.1000 103.2000 4.9000 103.5000 ;
	    RECT 3.1000 103.1000 3.4000 103.2000 ;
	    RECT 3.0000 101.1000 3.4000 103.1000 ;
	    RECT 4.6000 103.1000 4.9000 103.2000 ;
	    RECT 6.2000 104.1000 6.6000 107.9000 ;
	    RECT 7.0000 106.8000 7.4000 107.6000 ;
	    RECT 8.4000 107.1000 8.8000 109.9000 ;
	    RECT 7.9000 106.9000 8.8000 107.1000 ;
	    RECT 11.0000 107.9000 11.4000 109.9000 ;
	    RECT 12.6000 108.9000 13.0000 109.9000 ;
	    RECT 7.9000 106.8000 8.7000 106.9000 ;
	    RECT 7.9000 105.2000 8.2000 106.8000 ;
	    RECT 11.0000 106.2000 11.3000 107.9000 ;
	    RECT 12.6000 107.8000 12.9000 108.9000 ;
	    RECT 13.4000 107.8000 13.8000 108.6000 ;
	    RECT 11.7000 107.5000 12.9000 107.8000 ;
	    RECT 9.0000 105.8000 9.8000 106.2000 ;
	    RECT 11.0000 105.8000 11.4000 106.2000 ;
	    RECT 11.7000 106.0000 12.0000 107.5000 ;
	    RECT 14.8000 107.2000 15.2000 109.9000 ;
	    RECT 15.8000 107.8000 16.2000 108.2000 ;
	    RECT 14.8000 107.1000 15.4000 107.2000 ;
	    RECT 15.8000 107.1000 16.1000 107.8000 ;
	    RECT 14.3000 106.8000 16.1000 107.1000 ;
	    RECT 7.0000 104.8000 7.4000 105.2000 ;
	    RECT 7.8000 104.8000 8.2000 105.2000 ;
	    RECT 11.0000 105.1000 11.3000 105.8000 ;
	    RECT 11.7000 105.7000 12.1000 106.0000 ;
	    RECT 11.7000 105.6000 13.8000 105.7000 ;
	    RECT 11.8000 105.4000 13.8000 105.6000 ;
	    RECT 11.0000 104.8000 11.7000 105.1000 ;
	    RECT 7.0000 104.1000 7.3000 104.8000 ;
	    RECT 6.2000 103.8000 7.3000 104.1000 ;
	    RECT 4.6000 101.1000 5.0000 103.1000 ;
	    RECT 6.2000 101.1000 6.6000 103.8000 ;
	    RECT 7.9000 103.5000 8.2000 104.8000 ;
	    RECT 8.6000 103.8000 9.0000 104.6000 ;
	    RECT 7.9000 103.2000 9.7000 103.5000 ;
	    RECT 7.9000 103.1000 8.2000 103.2000 ;
	    RECT 7.8000 101.1000 8.2000 103.1000 ;
	    RECT 9.4000 101.1000 9.8000 103.2000 ;
	    RECT 11.3000 101.1000 11.7000 104.8000 ;
	    RECT 13.4000 101.1000 13.8000 105.4000 ;
	    RECT 14.3000 105.2000 14.6000 106.8000 ;
	    RECT 17.4000 106.2000 17.8000 109.9000 ;
	    RECT 19.0000 107.6000 19.4000 109.9000 ;
	    RECT 20.6000 108.9000 21.0000 109.9000 ;
	    RECT 19.8000 107.8000 20.2000 108.6000 ;
	    RECT 20.7000 107.8000 21.0000 108.9000 ;
	    RECT 22.2000 107.9000 22.6000 109.9000 ;
	    RECT 18.3000 107.3000 19.4000 107.6000 ;
	    RECT 20.7000 107.5000 21.9000 107.8000 ;
	    RECT 15.4000 105.8000 16.2000 106.2000 ;
	    RECT 14.2000 104.8000 14.6000 105.2000 ;
	    RECT 16.6000 104.8000 17.0000 105.6000 ;
	    RECT 17.4000 105.1000 17.7000 106.2000 ;
	    RECT 18.3000 105.8000 18.6000 107.3000 ;
	    RECT 21.6000 106.0000 21.9000 107.5000 ;
	    RECT 22.3000 107.2000 22.6000 107.9000 ;
	    RECT 22.2000 106.8000 22.6000 107.2000 ;
	    RECT 23.6000 107.1000 24.0000 109.9000 ;
	    RECT 22.3000 106.2000 22.6000 106.8000 ;
	    RECT 18.0000 105.4000 18.6000 105.8000 ;
	    RECT 21.5000 105.7000 21.9000 106.0000 ;
	    RECT 22.2000 105.8000 22.6000 106.2000 ;
	    RECT 18.3000 105.1000 18.6000 105.4000 ;
	    RECT 19.8000 105.6000 21.9000 105.7000 ;
	    RECT 19.8000 105.4000 21.8000 105.6000 ;
	    RECT 14.3000 103.5000 14.6000 104.8000 ;
	    RECT 15.0000 103.8000 15.4000 104.6000 ;
	    RECT 15.8000 104.1000 16.2000 104.2000 ;
	    RECT 17.4000 104.1000 17.8000 105.1000 ;
	    RECT 18.3000 104.8000 19.4000 105.1000 ;
	    RECT 15.8000 103.8000 17.8000 104.1000 ;
	    RECT 14.3000 103.2000 16.1000 103.5000 ;
	    RECT 14.3000 103.1000 14.6000 103.2000 ;
	    RECT 14.2000 101.1000 14.6000 103.1000 ;
	    RECT 15.8000 103.1000 16.1000 103.2000 ;
	    RECT 15.8000 101.1000 16.2000 103.1000 ;
	    RECT 17.4000 101.1000 17.8000 103.8000 ;
	    RECT 19.0000 101.1000 19.4000 104.8000 ;
	    RECT 19.8000 101.1000 20.2000 105.4000 ;
	    RECT 22.3000 105.1000 22.6000 105.8000 ;
	    RECT 23.1000 106.9000 24.0000 107.1000 ;
	    RECT 23.1000 106.8000 23.9000 106.9000 ;
	    RECT 23.1000 105.2000 23.4000 106.8000 ;
	    RECT 24.2000 105.8000 25.0000 106.2000 ;
	    RECT 21.9000 104.8000 22.6000 105.1000 ;
	    RECT 23.0000 104.8000 23.4000 105.2000 ;
	    RECT 25.4000 104.8000 25.8000 105.6000 ;
	    RECT 21.9000 101.1000 22.3000 104.8000 ;
	    RECT 23.1000 103.5000 23.4000 104.8000 ;
	    RECT 23.8000 103.8000 24.2000 104.6000 ;
	    RECT 23.1000 103.2000 24.9000 103.5000 ;
	    RECT 23.1000 103.1000 23.4000 103.2000 ;
	    RECT 23.0000 101.1000 23.4000 103.1000 ;
	    RECT 24.6000 103.1000 24.9000 103.2000 ;
	    RECT 24.6000 101.1000 25.0000 103.1000 ;
	    RECT 26.2000 101.1000 26.6000 109.9000 ;
	    RECT 29.6000 107.1000 30.0000 109.9000 ;
	    RECT 32.3000 109.2000 32.7000 109.9000 ;
	    RECT 31.8000 108.8000 32.7000 109.2000 ;
	    RECT 32.3000 108.2000 32.7000 108.8000 ;
	    RECT 31.8000 107.9000 32.7000 108.2000 ;
	    RECT 29.6000 106.9000 30.5000 107.1000 ;
	    RECT 29.7000 106.8000 30.5000 106.9000 ;
	    RECT 31.0000 106.8000 31.4000 107.6000 ;
	    RECT 28.6000 105.8000 29.4000 106.2000 ;
	    RECT 30.2000 106.1000 30.5000 106.8000 ;
	    RECT 30.2000 105.8000 31.3000 106.1000 ;
	    RECT 27.8000 104.8000 28.2000 105.6000 ;
	    RECT 30.2000 105.2000 30.5000 105.8000 ;
	    RECT 31.0000 105.2000 31.3000 105.8000 ;
	    RECT 30.2000 104.8000 30.6000 105.2000 ;
	    RECT 31.0000 104.8000 31.4000 105.2000 ;
	    RECT 29.4000 103.8000 29.8000 104.6000 ;
	    RECT 30.2000 103.5000 30.5000 104.8000 ;
	    RECT 28.7000 103.2000 30.5000 103.5000 ;
	    RECT 28.7000 103.1000 29.0000 103.2000 ;
	    RECT 28.6000 101.1000 29.0000 103.1000 ;
	    RECT 30.2000 103.1000 30.5000 103.2000 ;
	    RECT 30.2000 101.1000 30.6000 103.1000 ;
	    RECT 31.8000 101.1000 32.2000 107.9000 ;
	    RECT 32.6000 105.1000 33.0000 105.2000 ;
	    RECT 33.4000 105.1000 33.8000 109.9000 ;
	    RECT 35.6000 107.1000 36.0000 109.9000 ;
	    RECT 38.8000 107.1000 39.2000 109.9000 ;
	    RECT 42.2000 108.9000 42.6000 109.9000 ;
	    RECT 41.4000 107.8000 41.8000 108.6000 ;
	    RECT 42.3000 107.8000 42.6000 108.9000 ;
	    RECT 43.8000 107.9000 44.2000 109.9000 ;
	    RECT 42.3000 107.5000 43.5000 107.8000 ;
	    RECT 35.1000 106.9000 36.0000 107.1000 ;
	    RECT 38.3000 106.9000 39.2000 107.1000 ;
	    RECT 35.1000 106.8000 35.9000 106.9000 ;
	    RECT 38.3000 106.8000 39.1000 106.9000 ;
	    RECT 35.1000 105.2000 35.4000 106.8000 ;
	    RECT 36.2000 105.8000 37.0000 106.2000 ;
	    RECT 32.6000 104.8000 33.8000 105.1000 ;
	    RECT 35.0000 104.8000 35.4000 105.2000 ;
	    RECT 37.4000 104.8000 37.8000 105.6000 ;
	    RECT 38.3000 105.2000 38.6000 106.8000 ;
	    RECT 39.4000 105.8000 40.2000 106.2000 ;
	    RECT 43.2000 106.0000 43.5000 107.5000 ;
	    RECT 43.9000 106.2000 44.2000 107.9000 ;
	    RECT 43.1000 105.7000 43.5000 106.0000 ;
	    RECT 43.8000 105.8000 44.2000 106.2000 ;
	    RECT 41.4000 105.6000 43.5000 105.7000 ;
	    RECT 38.2000 104.8000 38.6000 105.2000 ;
	    RECT 40.6000 104.8000 41.0000 105.6000 ;
	    RECT 41.4000 105.4000 43.4000 105.6000 ;
	    RECT 32.6000 104.4000 33.0000 104.8000 ;
	    RECT 33.4000 101.1000 33.8000 104.8000 ;
	    RECT 35.1000 103.5000 35.4000 104.8000 ;
	    RECT 35.8000 103.8000 36.2000 104.6000 ;
	    RECT 38.3000 103.5000 38.6000 104.8000 ;
	    RECT 39.0000 103.8000 39.4000 104.6000 ;
	    RECT 35.1000 103.2000 36.9000 103.5000 ;
	    RECT 35.1000 103.1000 35.4000 103.2000 ;
	    RECT 35.0000 101.1000 35.4000 103.1000 ;
	    RECT 36.6000 103.1000 36.9000 103.2000 ;
	    RECT 38.3000 103.2000 40.1000 103.5000 ;
	    RECT 38.3000 103.1000 38.6000 103.2000 ;
	    RECT 36.6000 101.1000 37.0000 103.1000 ;
	    RECT 38.2000 101.1000 38.6000 103.1000 ;
	    RECT 39.8000 103.1000 40.1000 103.2000 ;
	    RECT 39.8000 101.1000 40.2000 103.1000 ;
	    RECT 41.4000 101.1000 41.8000 105.4000 ;
	    RECT 43.9000 105.1000 44.2000 105.8000 ;
	    RECT 43.5000 104.8000 44.2000 105.1000 ;
	    RECT 44.6000 105.1000 45.0000 109.9000 ;
	    RECT 46.5000 108.2000 46.9000 109.9000 ;
	    RECT 46.5000 107.9000 47.4000 108.2000 ;
	    RECT 46.2000 105.1000 46.6000 105.2000 ;
	    RECT 44.6000 104.8000 46.6000 105.1000 ;
	    RECT 43.5000 101.1000 43.9000 104.8000 ;
	    RECT 44.6000 101.1000 45.0000 104.8000 ;
	    RECT 46.2000 104.4000 46.6000 104.8000 ;
	    RECT 47.0000 104.1000 47.4000 107.9000 ;
	    RECT 47.8000 106.8000 48.2000 107.6000 ;
	    RECT 49.2000 107.1000 49.6000 109.9000 ;
	    RECT 52.6000 108.9000 53.0000 109.9000 ;
	    RECT 51.8000 107.8000 52.2000 108.6000 ;
	    RECT 52.7000 107.8000 53.0000 108.9000 ;
	    RECT 54.2000 107.9000 54.6000 109.9000 ;
	    RECT 52.7000 107.5000 53.9000 107.8000 ;
	    RECT 48.7000 106.9000 49.6000 107.1000 ;
	    RECT 48.7000 106.8000 49.5000 106.9000 ;
	    RECT 48.7000 105.2000 49.0000 106.8000 ;
	    RECT 49.8000 105.8000 50.6000 106.2000 ;
	    RECT 53.6000 106.0000 53.9000 107.5000 ;
	    RECT 54.3000 106.2000 54.6000 107.9000 ;
	    RECT 56.8000 107.1000 57.2000 109.9000 ;
	    RECT 59.5000 108.2000 59.9000 109.9000 ;
	    RECT 59.0000 107.9000 59.9000 108.2000 ;
	    RECT 56.8000 106.9000 57.7000 107.1000 ;
	    RECT 56.9000 106.8000 57.7000 106.9000 ;
	    RECT 58.2000 106.8000 58.6000 107.6000 ;
	    RECT 53.5000 105.7000 53.9000 106.0000 ;
	    RECT 54.2000 105.8000 54.6000 106.2000 ;
	    RECT 55.8000 105.8000 56.6000 106.2000 ;
	    RECT 57.4000 106.1000 57.7000 106.8000 ;
	    RECT 58.2000 106.1000 58.6000 106.2000 ;
	    RECT 57.4000 105.8000 58.6000 106.1000 ;
	    RECT 47.8000 104.8000 48.2000 105.2000 ;
	    RECT 48.6000 104.8000 49.0000 105.2000 ;
	    RECT 47.8000 104.1000 48.1000 104.8000 ;
	    RECT 47.0000 103.8000 48.1000 104.1000 ;
	    RECT 47.0000 101.1000 47.4000 103.8000 ;
	    RECT 48.7000 103.5000 49.0000 104.8000 ;
	    RECT 51.8000 105.6000 53.9000 105.7000 ;
	    RECT 51.8000 105.4000 53.8000 105.6000 ;
	    RECT 49.4000 103.8000 49.8000 104.6000 ;
	    RECT 50.2000 103.8000 50.6000 104.2000 ;
	    RECT 50.2000 103.5000 50.5000 103.8000 ;
	    RECT 48.7000 103.2000 50.5000 103.5000 ;
	    RECT 48.7000 103.1000 49.0000 103.2000 ;
	    RECT 48.6000 101.1000 49.0000 103.1000 ;
	    RECT 50.2000 103.1000 50.5000 103.2000 ;
	    RECT 50.2000 101.1000 50.6000 103.1000 ;
	    RECT 51.8000 101.1000 52.2000 105.4000 ;
	    RECT 54.3000 105.1000 54.6000 105.8000 ;
	    RECT 53.9000 104.8000 54.6000 105.1000 ;
	    RECT 55.0000 105.1000 55.4000 105.6000 ;
	    RECT 57.4000 105.2000 57.7000 105.8000 ;
	    RECT 55.8000 105.1000 56.2000 105.2000 ;
	    RECT 55.0000 104.8000 56.2000 105.1000 ;
	    RECT 57.4000 104.8000 57.8000 105.2000 ;
	    RECT 58.2000 104.8000 58.6000 105.2000 ;
	    RECT 53.9000 101.1000 54.3000 104.8000 ;
	    RECT 56.6000 103.8000 57.0000 104.6000 ;
	    RECT 57.4000 103.5000 57.7000 104.8000 ;
	    RECT 58.2000 104.1000 58.5000 104.8000 ;
	    RECT 59.0000 104.1000 59.4000 107.9000 ;
	    RECT 62.8000 107.1000 63.2000 109.9000 ;
	    RECT 66.0000 107.1000 66.4000 109.9000 ;
	    RECT 69.2000 107.1000 69.6000 109.9000 ;
	    RECT 62.3000 106.9000 63.2000 107.1000 ;
	    RECT 65.5000 106.9000 66.4000 107.1000 ;
	    RECT 68.7000 106.9000 69.6000 107.1000 ;
	    RECT 62.3000 106.8000 63.1000 106.9000 ;
	    RECT 65.5000 106.8000 66.3000 106.9000 ;
	    RECT 68.7000 106.8000 69.5000 106.9000 ;
	    RECT 62.3000 105.2000 62.6000 106.8000 ;
	    RECT 63.4000 105.8000 64.2000 106.2000 ;
	    RECT 59.8000 104.4000 60.2000 105.2000 ;
	    RECT 62.2000 104.8000 62.6000 105.2000 ;
	    RECT 64.6000 104.8000 65.0000 105.6000 ;
	    RECT 65.5000 105.2000 65.8000 106.8000 ;
	    RECT 66.6000 105.8000 67.4000 106.2000 ;
	    RECT 65.4000 104.8000 65.8000 105.2000 ;
	    RECT 67.8000 104.8000 68.2000 105.6000 ;
	    RECT 68.7000 105.2000 69.0000 106.8000 ;
	    RECT 69.8000 105.8000 70.6000 106.2000 ;
	    RECT 72.6000 106.1000 73.0000 109.9000 ;
	    RECT 73.4000 106.1000 73.8000 106.2000 ;
	    RECT 72.6000 105.8000 73.8000 106.1000 ;
	    RECT 68.6000 104.8000 69.0000 105.2000 ;
	    RECT 58.2000 103.8000 59.4000 104.1000 ;
	    RECT 55.9000 103.2000 57.7000 103.5000 ;
	    RECT 55.9000 103.1000 56.2000 103.2000 ;
	    RECT 55.8000 101.1000 56.2000 103.1000 ;
	    RECT 57.4000 103.1000 57.7000 103.2000 ;
	    RECT 57.4000 101.1000 57.8000 103.1000 ;
	    RECT 59.0000 101.1000 59.4000 103.8000 ;
	    RECT 62.3000 103.5000 62.6000 104.8000 ;
	    RECT 63.0000 103.8000 63.4000 104.6000 ;
	    RECT 65.5000 103.5000 65.8000 104.8000 ;
	    RECT 66.2000 103.8000 66.6000 104.6000 ;
	    RECT 67.0000 103.8000 67.4000 104.2000 ;
	    RECT 67.0000 103.5000 67.3000 103.8000 ;
	    RECT 62.3000 103.2000 64.1000 103.5000 ;
	    RECT 65.5000 103.2000 67.3000 103.5000 ;
	    RECT 62.3000 103.1000 62.6000 103.2000 ;
	    RECT 62.2000 101.1000 62.6000 103.1000 ;
	    RECT 63.8000 101.1000 64.2000 103.2000 ;
	    RECT 65.5000 103.1000 65.8000 103.2000 ;
	    RECT 65.4000 101.1000 65.8000 103.1000 ;
	    RECT 67.0000 103.1000 67.3000 103.2000 ;
	    RECT 68.7000 103.5000 69.0000 104.8000 ;
	    RECT 69.4000 103.8000 69.8000 104.6000 ;
	    RECT 68.7000 103.2000 70.5000 103.5000 ;
	    RECT 68.7000 103.1000 69.0000 103.2000 ;
	    RECT 67.0000 101.1000 67.4000 103.1000 ;
	    RECT 68.6000 101.1000 69.0000 103.1000 ;
	    RECT 70.2000 103.1000 70.5000 103.2000 ;
	    RECT 70.2000 101.1000 70.6000 103.1000 ;
	    RECT 72.6000 101.1000 73.0000 105.8000 ;
	    RECT 75.0000 101.1000 75.4000 109.9000 ;
	    RECT 75.8000 101.1000 76.2000 109.9000 ;
	    RECT 78.0000 107.1000 78.4000 109.9000 ;
	    RECT 81.2000 107.1000 81.6000 109.9000 ;
	    RECT 77.5000 106.9000 78.4000 107.1000 ;
	    RECT 80.7000 106.9000 81.6000 107.1000 ;
	    RECT 85.6000 107.1000 86.0000 109.9000 ;
	    RECT 88.8000 107.1000 89.2000 109.9000 ;
	    RECT 90.8000 107.1000 91.2000 109.9000 ;
	    RECT 93.4000 107.5000 93.8000 109.9000 ;
	    RECT 95.6000 109.2000 96.0000 109.9000 ;
	    RECT 95.0000 108.9000 96.0000 109.2000 ;
	    RECT 97.8000 108.9000 98.2000 109.9000 ;
	    RECT 99.9000 109.2000 100.5000 109.9000 ;
	    RECT 99.8000 108.9000 100.5000 109.2000 ;
	    RECT 95.0000 108.5000 95.4000 108.9000 ;
	    RECT 97.8000 108.6000 98.1000 108.9000 ;
	    RECT 95.8000 108.2000 96.2000 108.6000 ;
	    RECT 96.7000 108.3000 98.1000 108.6000 ;
	    RECT 99.8000 108.5000 100.2000 108.9000 ;
	    RECT 96.7000 108.2000 97.1000 108.3000 ;
	    RECT 85.6000 106.9000 86.5000 107.1000 ;
	    RECT 88.8000 106.9000 89.7000 107.1000 ;
	    RECT 77.5000 106.8000 78.3000 106.9000 ;
	    RECT 80.7000 106.8000 81.5000 106.9000 ;
	    RECT 85.7000 106.8000 86.5000 106.9000 ;
	    RECT 88.9000 106.8000 89.7000 106.9000 ;
	    RECT 77.5000 105.2000 77.8000 106.8000 ;
	    RECT 78.6000 105.8000 79.4000 106.2000 ;
	    RECT 77.4000 104.8000 77.8000 105.2000 ;
	    RECT 79.8000 104.8000 80.2000 105.6000 ;
	    RECT 80.7000 105.2000 81.0000 106.8000 ;
	    RECT 81.8000 105.8000 82.6000 106.2000 ;
	    RECT 84.6000 105.8000 85.4000 106.2000 ;
	    RECT 80.6000 104.8000 81.0000 105.2000 ;
	    RECT 83.0000 104.8000 83.4000 105.6000 ;
	    RECT 83.8000 104.8000 84.2000 105.6000 ;
	    RECT 86.2000 105.2000 86.5000 106.8000 ;
	    RECT 89.4000 106.2000 89.7000 106.8000 ;
	    RECT 90.3000 106.9000 91.2000 107.1000 ;
	    RECT 93.8000 107.1000 94.6000 107.2000 ;
	    RECT 95.9000 107.1000 96.2000 108.2000 ;
	    RECT 100.7000 107.7000 101.1000 107.8000 ;
	    RECT 102.2000 107.7000 102.6000 109.9000 ;
	    RECT 103.3000 109.2000 103.7000 109.9000 ;
	    RECT 103.0000 108.8000 103.7000 109.2000 ;
	    RECT 103.3000 108.4000 103.7000 108.8000 ;
	    RECT 100.7000 107.4000 102.6000 107.7000 ;
	    RECT 98.7000 107.1000 99.1000 107.2000 ;
	    RECT 90.3000 106.8000 91.1000 106.9000 ;
	    RECT 93.8000 106.8000 99.3000 107.1000 ;
	    RECT 87.8000 105.8000 88.6000 106.2000 ;
	    RECT 89.4000 105.8000 89.8000 106.2000 ;
	    RECT 86.2000 104.8000 86.6000 105.2000 ;
	    RECT 87.0000 104.8000 87.4000 105.6000 ;
	    RECT 89.4000 105.2000 89.7000 105.8000 ;
	    RECT 90.3000 105.2000 90.6000 106.8000 ;
	    RECT 95.3000 106.7000 95.7000 106.8000 ;
	    RECT 94.5000 106.2000 94.9000 106.3000 ;
	    RECT 99.0000 106.2000 99.3000 106.8000 ;
	    RECT 99.8000 106.4000 100.2000 106.5000 ;
	    RECT 91.4000 105.8000 92.2000 106.2000 ;
	    RECT 94.5000 105.9000 97.0000 106.2000 ;
	    RECT 96.6000 105.8000 97.0000 105.9000 ;
	    RECT 99.0000 105.8000 99.4000 106.2000 ;
	    RECT 99.8000 106.1000 101.7000 106.4000 ;
	    RECT 101.3000 106.0000 101.7000 106.1000 ;
	    RECT 89.4000 104.8000 89.8000 105.2000 ;
	    RECT 90.2000 104.8000 90.6000 105.2000 ;
	    RECT 92.6000 104.8000 93.0000 105.6000 ;
	    RECT 93.4000 105.5000 96.2000 105.6000 ;
	    RECT 93.4000 105.4000 96.3000 105.5000 ;
	    RECT 93.4000 105.3000 98.3000 105.4000 ;
	    RECT 77.5000 103.5000 77.8000 104.8000 ;
	    RECT 78.2000 103.8000 78.6000 104.6000 ;
	    RECT 80.7000 103.5000 81.0000 104.8000 ;
	    RECT 81.4000 103.8000 81.8000 104.6000 ;
	    RECT 85.4000 103.8000 85.8000 104.6000 ;
	    RECT 86.2000 103.5000 86.5000 104.8000 ;
	    RECT 88.6000 103.8000 89.0000 104.6000 ;
	    RECT 89.4000 103.5000 89.7000 104.8000 ;
	    RECT 77.5000 103.2000 79.3000 103.5000 ;
	    RECT 77.5000 103.1000 77.8000 103.2000 ;
	    RECT 77.4000 101.1000 77.8000 103.1000 ;
	    RECT 79.0000 103.1000 79.3000 103.2000 ;
	    RECT 80.7000 103.2000 82.5000 103.5000 ;
	    RECT 80.7000 103.1000 81.0000 103.2000 ;
	    RECT 79.0000 101.1000 79.4000 103.1000 ;
	    RECT 80.6000 101.1000 81.0000 103.1000 ;
	    RECT 82.2000 103.1000 82.5000 103.2000 ;
	    RECT 84.7000 103.2000 86.5000 103.5000 ;
	    RECT 84.7000 103.1000 85.0000 103.2000 ;
	    RECT 82.2000 101.1000 82.6000 103.1000 ;
	    RECT 84.6000 101.1000 85.0000 103.1000 ;
	    RECT 86.2000 103.1000 86.5000 103.2000 ;
	    RECT 87.9000 103.2000 89.7000 103.5000 ;
	    RECT 87.9000 103.1000 88.2000 103.2000 ;
	    RECT 86.2000 101.1000 86.6000 103.1000 ;
	    RECT 87.8000 101.1000 88.2000 103.1000 ;
	    RECT 89.4000 103.1000 89.7000 103.2000 ;
	    RECT 90.3000 103.5000 90.6000 104.8000 ;
	    RECT 91.0000 103.8000 91.4000 104.6000 ;
	    RECT 90.3000 103.2000 92.1000 103.5000 ;
	    RECT 90.3000 103.1000 90.6000 103.2000 ;
	    RECT 89.4000 101.1000 89.8000 103.1000 ;
	    RECT 90.2000 101.1000 90.6000 103.1000 ;
	    RECT 91.8000 103.1000 92.1000 103.2000 ;
	    RECT 91.8000 101.1000 92.2000 103.1000 ;
	    RECT 93.4000 101.1000 93.8000 105.3000 ;
	    RECT 95.9000 105.1000 98.3000 105.3000 ;
	    RECT 95.0000 104.5000 97.7000 104.8000 ;
	    RECT 95.0000 104.4000 95.4000 104.5000 ;
	    RECT 97.3000 104.4000 97.7000 104.5000 ;
	    RECT 98.0000 104.5000 98.3000 105.1000 ;
	    RECT 99.0000 105.2000 99.3000 105.8000 ;
	    RECT 100.5000 105.7000 100.9000 105.8000 ;
	    RECT 102.2000 105.7000 102.6000 107.4000 ;
	    RECT 100.5000 105.4000 102.6000 105.7000 ;
	    RECT 99.0000 104.9000 100.2000 105.2000 ;
	    RECT 98.7000 104.5000 99.1000 104.6000 ;
	    RECT 98.0000 104.2000 99.1000 104.5000 ;
	    RECT 99.9000 104.4000 100.2000 104.9000 ;
	    RECT 99.9000 104.0000 100.6000 104.4000 ;
	    RECT 96.7000 103.7000 97.1000 103.8000 ;
	    RECT 98.1000 103.7000 98.5000 103.8000 ;
	    RECT 95.0000 103.1000 95.4000 103.5000 ;
	    RECT 96.7000 103.4000 98.5000 103.7000 ;
	    RECT 97.8000 103.1000 98.1000 103.4000 ;
	    RECT 99.8000 103.1000 100.2000 103.5000 ;
	    RECT 95.0000 102.8000 96.0000 103.1000 ;
	    RECT 95.6000 101.1000 96.0000 102.8000 ;
	    RECT 97.8000 101.1000 98.2000 103.1000 ;
	    RECT 99.9000 101.1000 100.5000 103.1000 ;
	    RECT 102.2000 101.1000 102.6000 105.4000 ;
	    RECT 103.0000 107.9000 103.7000 108.4000 ;
	    RECT 105.4000 107.9000 105.8000 109.9000 ;
	    RECT 106.2000 107.9000 106.6000 109.9000 ;
	    RECT 108.3000 108.4000 108.7000 109.9000 ;
	    RECT 108.3000 107.9000 109.0000 108.4000 ;
	    RECT 103.0000 106.2000 103.3000 107.9000 ;
	    RECT 105.4000 107.8000 105.7000 107.9000 ;
	    RECT 104.8000 107.6000 105.7000 107.8000 ;
	    RECT 103.6000 107.5000 105.7000 107.6000 ;
	    RECT 106.3000 107.8000 106.6000 107.9000 ;
	    RECT 106.3000 107.6000 107.2000 107.8000 ;
	    RECT 106.3000 107.5000 108.4000 107.6000 ;
	    RECT 103.6000 107.3000 105.1000 107.5000 ;
	    RECT 106.9000 107.3000 108.4000 107.5000 ;
	    RECT 103.6000 107.2000 104.0000 107.3000 ;
	    RECT 108.0000 107.2000 108.4000 107.3000 ;
	    RECT 103.0000 105.8000 103.4000 106.2000 ;
	    RECT 103.0000 105.1000 103.3000 105.8000 ;
	    RECT 103.7000 105.5000 104.0000 107.2000 ;
	    RECT 105.4000 107.1000 105.8000 107.2000 ;
	    RECT 106.2000 107.1000 106.6000 107.2000 ;
	    RECT 104.4000 106.6000 105.0000 107.0000 ;
	    RECT 105.4000 106.8000 106.6000 107.1000 ;
	    RECT 107.2000 106.9000 107.6000 107.0000 ;
	    RECT 104.6000 106.2000 104.9000 106.6000 ;
	    RECT 105.4000 106.4000 105.8000 106.8000 ;
	    RECT 106.2000 106.4000 106.6000 106.8000 ;
	    RECT 107.1000 106.6000 107.6000 106.9000 ;
	    RECT 107.1000 106.2000 107.4000 106.6000 ;
	    RECT 104.6000 105.8000 105.0000 106.2000 ;
	    RECT 107.0000 105.8000 107.4000 106.2000 ;
	    RECT 108.0000 105.5000 108.3000 107.2000 ;
	    RECT 108.7000 106.2000 109.0000 107.9000 ;
	    RECT 111.0000 107.7000 111.4000 109.9000 ;
	    RECT 113.1000 109.2000 113.7000 109.9000 ;
	    RECT 113.1000 108.9000 113.8000 109.2000 ;
	    RECT 115.4000 108.9000 115.8000 109.9000 ;
	    RECT 117.6000 109.2000 118.0000 109.9000 ;
	    RECT 117.6000 108.9000 118.6000 109.2000 ;
	    RECT 113.4000 108.5000 113.8000 108.9000 ;
	    RECT 115.5000 108.6000 115.8000 108.9000 ;
	    RECT 115.5000 108.3000 116.9000 108.6000 ;
	    RECT 116.5000 108.2000 116.9000 108.3000 ;
	    RECT 117.4000 108.2000 117.8000 108.6000 ;
	    RECT 118.2000 108.5000 118.6000 108.9000 ;
	    RECT 112.5000 107.7000 112.9000 107.8000 ;
	    RECT 111.0000 107.4000 112.9000 107.7000 ;
	    RECT 108.6000 106.1000 109.0000 106.2000 ;
	    RECT 109.4000 106.1000 109.8000 106.2000 ;
	    RECT 108.6000 105.8000 109.8000 106.1000 ;
	    RECT 103.7000 105.2000 104.9000 105.5000 ;
	    RECT 103.0000 101.1000 103.4000 105.1000 ;
	    RECT 104.6000 103.1000 104.9000 105.2000 ;
	    RECT 107.1000 105.2000 108.3000 105.5000 ;
	    RECT 107.1000 103.1000 107.4000 105.2000 ;
	    RECT 108.7000 105.1000 109.0000 105.8000 ;
	    RECT 104.6000 101.1000 105.0000 103.1000 ;
	    RECT 107.0000 101.1000 107.4000 103.1000 ;
	    RECT 108.6000 101.1000 109.0000 105.1000 ;
	    RECT 111.0000 105.7000 111.4000 107.4000 ;
	    RECT 114.2000 107.1000 114.9000 107.2000 ;
	    RECT 117.4000 107.1000 117.7000 108.2000 ;
	    RECT 119.8000 107.5000 120.2000 109.9000 ;
	    RECT 120.9000 109.2000 121.3000 109.9000 ;
	    RECT 120.6000 108.8000 121.3000 109.2000 ;
	    RECT 120.9000 108.4000 121.3000 108.8000 ;
	    RECT 120.6000 107.9000 121.3000 108.4000 ;
	    RECT 123.0000 107.9000 123.4000 109.9000 ;
	    RECT 123.8000 107.9000 124.2000 109.9000 ;
	    RECT 125.9000 108.4000 126.3000 109.9000 ;
	    RECT 127.0000 109.6000 129.0000 109.9000 ;
	    RECT 125.9000 107.9000 126.6000 108.4000 ;
	    RECT 127.0000 107.9000 127.4000 109.6000 ;
	    RECT 127.8000 107.9000 128.2000 109.3000 ;
	    RECT 128.6000 108.0000 129.0000 109.6000 ;
	    RECT 130.2000 108.0000 130.6000 109.9000 ;
	    RECT 128.6000 107.9000 130.6000 108.0000 ;
	    RECT 119.0000 107.1000 119.8000 107.2000 ;
	    RECT 114.2000 106.8000 119.8000 107.1000 ;
	    RECT 113.4000 106.4000 113.8000 106.5000 ;
	    RECT 111.9000 106.1000 113.8000 106.4000 ;
	    RECT 111.9000 106.0000 112.3000 106.1000 ;
	    RECT 112.7000 105.7000 113.1000 105.8000 ;
	    RECT 111.0000 105.4000 113.1000 105.7000 ;
	    RECT 111.0000 101.1000 111.4000 105.4000 ;
	    RECT 114.3000 105.2000 114.6000 106.8000 ;
	    RECT 117.9000 106.7000 118.3000 106.8000 ;
	    RECT 118.7000 106.2000 119.1000 106.3000 ;
	    RECT 116.6000 105.9000 119.1000 106.2000 ;
	    RECT 120.6000 106.2000 120.9000 107.9000 ;
	    RECT 123.0000 107.8000 123.3000 107.9000 ;
	    RECT 122.4000 107.6000 123.3000 107.8000 ;
	    RECT 121.2000 107.5000 123.3000 107.6000 ;
	    RECT 123.9000 107.8000 124.2000 107.9000 ;
	    RECT 123.9000 107.6000 124.8000 107.8000 ;
	    RECT 123.9000 107.5000 126.0000 107.6000 ;
	    RECT 121.2000 107.3000 122.7000 107.5000 ;
	    RECT 124.5000 107.3000 126.0000 107.5000 ;
	    RECT 121.2000 107.2000 121.6000 107.3000 ;
	    RECT 125.6000 107.2000 126.0000 107.3000 ;
	    RECT 116.6000 105.8000 117.0000 105.9000 ;
	    RECT 120.6000 105.8000 121.0000 106.2000 ;
	    RECT 117.4000 105.5000 120.2000 105.6000 ;
	    RECT 117.3000 105.4000 120.2000 105.5000 ;
	    RECT 113.4000 104.9000 114.6000 105.2000 ;
	    RECT 115.3000 105.3000 120.2000 105.4000 ;
	    RECT 115.3000 105.1000 117.7000 105.3000 ;
	    RECT 113.4000 104.4000 113.7000 104.9000 ;
	    RECT 113.0000 104.0000 113.7000 104.4000 ;
	    RECT 114.5000 104.5000 114.9000 104.6000 ;
	    RECT 115.3000 104.5000 115.6000 105.1000 ;
	    RECT 114.5000 104.2000 115.6000 104.5000 ;
	    RECT 115.9000 104.5000 118.6000 104.8000 ;
	    RECT 115.9000 104.4000 116.3000 104.5000 ;
	    RECT 118.2000 104.4000 118.6000 104.5000 ;
	    RECT 115.1000 103.7000 115.5000 103.8000 ;
	    RECT 116.5000 103.7000 116.9000 103.8000 ;
	    RECT 113.4000 103.1000 113.8000 103.5000 ;
	    RECT 115.1000 103.4000 116.9000 103.7000 ;
	    RECT 115.5000 103.1000 115.8000 103.4000 ;
	    RECT 118.2000 103.1000 118.6000 103.5000 ;
	    RECT 113.1000 101.1000 113.7000 103.1000 ;
	    RECT 115.4000 101.1000 115.8000 103.1000 ;
	    RECT 117.6000 102.8000 118.6000 103.1000 ;
	    RECT 117.6000 101.1000 118.0000 102.8000 ;
	    RECT 119.8000 101.1000 120.2000 105.3000 ;
	    RECT 120.6000 105.1000 120.9000 105.8000 ;
	    RECT 121.3000 105.5000 121.6000 107.2000 ;
	    RECT 122.0000 106.9000 122.4000 107.0000 ;
	    RECT 122.0000 106.6000 122.5000 106.9000 ;
	    RECT 122.2000 106.2000 122.5000 106.6000 ;
	    RECT 123.0000 106.4000 123.4000 107.2000 ;
	    RECT 123.8000 106.4000 124.2000 107.2000 ;
	    RECT 124.8000 106.9000 125.2000 107.0000 ;
	    RECT 124.7000 106.6000 125.2000 106.9000 ;
	    RECT 124.7000 106.2000 125.0000 106.6000 ;
	    RECT 122.2000 105.8000 122.6000 106.2000 ;
	    RECT 124.6000 105.8000 125.0000 106.2000 ;
	    RECT 125.6000 105.5000 125.9000 107.2000 ;
	    RECT 126.3000 106.2000 126.6000 107.9000 ;
	    RECT 127.8000 107.2000 128.1000 107.9000 ;
	    RECT 128.7000 107.7000 130.5000 107.9000 ;
	    RECT 131.0000 107.8000 131.4000 108.6000 ;
	    RECT 129.8000 107.2000 130.2000 107.4000 ;
	    RECT 126.2000 106.1000 126.6000 106.2000 ;
	    RECT 127.0000 106.1000 127.4000 107.2000 ;
	    RECT 127.8000 106.9000 129.0000 107.2000 ;
	    RECT 129.8000 106.9000 130.6000 107.2000 ;
	    RECT 128.6000 106.8000 129.0000 106.9000 ;
	    RECT 130.2000 106.8000 130.6000 106.9000 ;
	    RECT 126.2000 105.8000 127.4000 106.1000 ;
	    RECT 127.8000 105.8000 128.2000 106.6000 ;
	    RECT 121.3000 105.2000 122.5000 105.5000 ;
	    RECT 120.6000 101.1000 121.0000 105.1000 ;
	    RECT 122.2000 103.1000 122.5000 105.2000 ;
	    RECT 124.7000 105.2000 125.9000 105.5000 ;
	    RECT 124.7000 103.1000 125.0000 105.2000 ;
	    RECT 126.3000 105.1000 126.6000 105.8000 ;
	    RECT 128.7000 105.1000 129.0000 106.8000 ;
	    RECT 129.4000 105.8000 129.8000 106.6000 ;
	    RECT 131.8000 106.1000 132.2000 109.9000 ;
	    RECT 133.9000 107.9000 134.7000 109.9000 ;
	    RECT 136.9000 108.2000 137.3000 109.9000 ;
	    RECT 140.3000 109.2000 140.7000 109.9000 ;
	    RECT 140.3000 108.8000 141.0000 109.2000 ;
	    RECT 140.3000 108.2000 140.7000 108.8000 ;
	    RECT 136.9000 107.9000 137.8000 108.2000 ;
	    RECT 133.4000 106.8000 133.8000 107.2000 ;
	    RECT 133.5000 106.6000 133.8000 106.8000 ;
	    RECT 133.5000 106.2000 133.9000 106.6000 ;
	    RECT 134.2000 106.2000 134.5000 107.9000 ;
	    RECT 135.0000 107.1000 135.4000 107.2000 ;
	    RECT 135.8000 107.1000 136.2000 107.2000 ;
	    RECT 135.0000 106.8000 136.2000 107.1000 ;
	    RECT 135.0000 106.4000 135.4000 106.8000 ;
	    RECT 132.6000 106.1000 133.0000 106.2000 ;
	    RECT 131.8000 105.8000 133.0000 106.1000 ;
	    RECT 122.2000 101.1000 122.6000 103.1000 ;
	    RECT 124.6000 101.1000 125.0000 103.1000 ;
	    RECT 126.2000 101.1000 126.6000 105.1000 ;
	    RECT 128.3000 101.1000 129.3000 105.1000 ;
	    RECT 131.8000 101.1000 132.2000 105.8000 ;
	    RECT 132.6000 105.4000 133.0000 105.8000 ;
	    RECT 134.2000 105.8000 134.6000 106.2000 ;
	    RECT 135.8000 106.1000 136.2000 106.2000 ;
	    RECT 137.4000 106.1000 137.8000 107.9000 ;
	    RECT 139.8000 107.9000 140.7000 108.2000 ;
	    RECT 138.2000 106.8000 138.6000 107.6000 ;
	    RECT 139.0000 106.8000 139.4000 107.6000 ;
	    RECT 135.4000 105.8000 137.8000 106.1000 ;
	    RECT 134.2000 105.7000 134.5000 105.8000 ;
	    RECT 133.5000 105.4000 134.5000 105.7000 ;
	    RECT 135.4000 105.6000 135.8000 105.8000 ;
	    RECT 133.5000 105.1000 133.8000 105.4000 ;
	    RECT 132.6000 101.4000 133.0000 105.1000 ;
	    RECT 133.4000 101.7000 133.8000 105.1000 ;
	    RECT 134.2000 104.8000 136.2000 105.1000 ;
	    RECT 134.2000 101.4000 134.6000 104.8000 ;
	    RECT 132.6000 101.1000 134.6000 101.4000 ;
	    RECT 135.8000 101.1000 136.2000 104.8000 ;
	    RECT 136.6000 104.4000 137.0000 105.2000 ;
	    RECT 137.4000 101.1000 137.8000 105.8000 ;
	    RECT 139.8000 101.1000 140.2000 107.9000 ;
	    RECT 140.6000 105.1000 141.0000 105.2000 ;
	    RECT 141.4000 105.1000 141.8000 109.9000 ;
	    RECT 142.2000 107.8000 142.6000 108.6000 ;
	    RECT 143.0000 107.5000 143.4000 109.9000 ;
	    RECT 145.2000 109.2000 145.6000 109.9000 ;
	    RECT 144.6000 108.9000 145.6000 109.2000 ;
	    RECT 147.4000 108.9000 147.8000 109.9000 ;
	    RECT 149.5000 109.2000 150.1000 109.9000 ;
	    RECT 149.4000 108.9000 150.1000 109.2000 ;
	    RECT 144.6000 108.5000 145.0000 108.9000 ;
	    RECT 147.4000 108.6000 147.7000 108.9000 ;
	    RECT 145.4000 108.2000 145.8000 108.6000 ;
	    RECT 146.3000 108.3000 147.7000 108.6000 ;
	    RECT 149.4000 108.5000 149.8000 108.9000 ;
	    RECT 146.3000 108.2000 146.7000 108.3000 ;
	    RECT 143.4000 107.1000 144.2000 107.2000 ;
	    RECT 145.5000 107.1000 145.8000 108.2000 ;
	    RECT 150.3000 107.7000 150.7000 107.8000 ;
	    RECT 151.8000 107.7000 152.2000 109.9000 ;
	    RECT 150.3000 107.4000 152.2000 107.7000 ;
	    RECT 146.2000 107.1000 146.6000 107.2000 ;
	    RECT 148.3000 107.1000 148.7000 107.2000 ;
	    RECT 143.4000 106.8000 148.9000 107.1000 ;
	    RECT 144.9000 106.7000 145.3000 106.8000 ;
	    RECT 144.1000 106.2000 144.5000 106.3000 ;
	    RECT 145.4000 106.2000 145.8000 106.3000 ;
	    RECT 144.1000 105.9000 146.6000 106.2000 ;
	    RECT 146.2000 105.8000 146.6000 105.9000 ;
	    RECT 140.6000 104.8000 141.8000 105.1000 ;
	    RECT 140.6000 104.4000 141.0000 104.8000 ;
	    RECT 141.4000 101.1000 141.8000 104.8000 ;
	    RECT 143.0000 105.5000 145.8000 105.6000 ;
	    RECT 143.0000 105.4000 145.9000 105.5000 ;
	    RECT 143.0000 105.3000 147.9000 105.4000 ;
	    RECT 143.0000 101.1000 143.4000 105.3000 ;
	    RECT 145.5000 105.1000 147.9000 105.3000 ;
	    RECT 144.6000 104.5000 147.3000 104.8000 ;
	    RECT 144.6000 104.4000 145.0000 104.5000 ;
	    RECT 146.9000 104.4000 147.3000 104.5000 ;
	    RECT 147.6000 104.5000 147.9000 105.1000 ;
	    RECT 148.6000 105.2000 148.9000 106.8000 ;
	    RECT 149.4000 106.4000 149.8000 106.5000 ;
	    RECT 149.4000 106.1000 151.3000 106.4000 ;
	    RECT 150.9000 106.0000 151.3000 106.1000 ;
	    RECT 150.1000 105.7000 150.5000 105.8000 ;
	    RECT 151.8000 105.7000 152.2000 107.4000 ;
	    RECT 150.1000 105.4000 152.2000 105.7000 ;
	    RECT 148.6000 104.9000 149.8000 105.2000 ;
	    RECT 148.3000 104.5000 148.7000 104.6000 ;
	    RECT 147.6000 104.2000 148.7000 104.5000 ;
	    RECT 149.5000 104.4000 149.8000 104.9000 ;
	    RECT 149.5000 104.0000 150.2000 104.4000 ;
	    RECT 146.3000 103.7000 146.7000 103.8000 ;
	    RECT 147.7000 103.7000 148.1000 103.8000 ;
	    RECT 144.6000 103.1000 145.0000 103.5000 ;
	    RECT 146.3000 103.4000 148.1000 103.7000 ;
	    RECT 147.4000 103.1000 147.7000 103.4000 ;
	    RECT 149.4000 103.1000 149.8000 103.5000 ;
	    RECT 144.6000 102.8000 145.6000 103.1000 ;
	    RECT 145.2000 101.1000 145.6000 102.8000 ;
	    RECT 147.4000 101.1000 147.8000 103.1000 ;
	    RECT 149.5000 101.1000 150.1000 103.1000 ;
	    RECT 151.8000 101.1000 152.2000 105.4000 ;
	    RECT 152.6000 107.7000 153.0000 109.9000 ;
	    RECT 154.7000 109.2000 155.3000 109.9000 ;
	    RECT 154.7000 108.9000 155.4000 109.2000 ;
	    RECT 157.0000 108.9000 157.4000 109.9000 ;
	    RECT 159.2000 109.2000 159.6000 109.9000 ;
	    RECT 159.2000 108.9000 160.2000 109.2000 ;
	    RECT 155.0000 108.5000 155.4000 108.9000 ;
	    RECT 157.1000 108.6000 157.4000 108.9000 ;
	    RECT 157.1000 108.3000 158.5000 108.6000 ;
	    RECT 158.1000 108.2000 158.5000 108.3000 ;
	    RECT 159.0000 108.2000 159.4000 108.6000 ;
	    RECT 159.8000 108.5000 160.2000 108.9000 ;
	    RECT 154.1000 107.7000 154.5000 107.8000 ;
	    RECT 152.6000 107.4000 154.5000 107.7000 ;
	    RECT 152.6000 105.7000 153.0000 107.4000 ;
	    RECT 156.1000 107.1000 156.5000 107.2000 ;
	    RECT 159.0000 107.1000 159.3000 108.2000 ;
	    RECT 161.4000 107.5000 161.8000 109.9000 ;
	    RECT 162.2000 107.5000 162.6000 109.9000 ;
	    RECT 164.4000 109.2000 164.8000 109.9000 ;
	    RECT 163.8000 108.9000 164.8000 109.2000 ;
	    RECT 166.6000 108.9000 167.0000 109.9000 ;
	    RECT 168.7000 109.2000 169.3000 109.9000 ;
	    RECT 168.6000 108.9000 169.3000 109.2000 ;
	    RECT 163.8000 108.5000 164.2000 108.9000 ;
	    RECT 166.6000 108.6000 166.9000 108.9000 ;
	    RECT 164.6000 108.2000 165.0000 108.6000 ;
	    RECT 165.5000 108.3000 166.9000 108.6000 ;
	    RECT 168.6000 108.5000 169.0000 108.9000 ;
	    RECT 165.5000 108.2000 165.9000 108.3000 ;
	    RECT 160.6000 107.1000 161.4000 107.2000 ;
	    RECT 155.9000 106.8000 161.4000 107.1000 ;
	    RECT 162.6000 107.1000 163.4000 107.2000 ;
	    RECT 164.7000 107.1000 165.0000 108.2000 ;
	    RECT 169.5000 107.7000 169.9000 107.8000 ;
	    RECT 171.0000 107.7000 171.4000 109.9000 ;
	    RECT 169.5000 107.4000 171.4000 107.7000 ;
	    RECT 165.4000 107.1000 165.8000 107.2000 ;
	    RECT 167.5000 107.1000 167.9000 107.2000 ;
	    RECT 162.6000 106.8000 168.1000 107.1000 ;
	    RECT 155.0000 106.4000 155.4000 106.5000 ;
	    RECT 153.5000 106.1000 155.4000 106.4000 ;
	    RECT 155.9000 106.2000 156.2000 106.8000 ;
	    RECT 159.5000 106.7000 159.9000 106.8000 ;
	    RECT 164.1000 106.7000 164.5000 106.8000 ;
	    RECT 159.0000 106.2000 159.4000 106.3000 ;
	    RECT 160.3000 106.2000 160.7000 106.3000 ;
	    RECT 153.5000 106.0000 153.9000 106.1000 ;
	    RECT 155.8000 105.8000 156.2000 106.2000 ;
	    RECT 158.2000 105.9000 160.7000 106.2000 ;
	    RECT 163.3000 106.2000 163.7000 106.3000 ;
	    RECT 164.6000 106.2000 165.0000 106.3000 ;
	    RECT 163.3000 105.9000 165.8000 106.2000 ;
	    RECT 158.2000 105.8000 158.6000 105.9000 ;
	    RECT 165.4000 105.8000 165.8000 105.9000 ;
	    RECT 154.3000 105.7000 154.7000 105.8000 ;
	    RECT 152.6000 105.4000 154.7000 105.7000 ;
	    RECT 152.6000 101.1000 153.0000 105.4000 ;
	    RECT 155.9000 105.2000 156.2000 105.8000 ;
	    RECT 159.0000 105.5000 161.8000 105.6000 ;
	    RECT 158.9000 105.4000 161.8000 105.5000 ;
	    RECT 155.0000 104.9000 156.2000 105.2000 ;
	    RECT 156.9000 105.3000 161.8000 105.4000 ;
	    RECT 156.9000 105.1000 159.3000 105.3000 ;
	    RECT 155.0000 104.4000 155.3000 104.9000 ;
	    RECT 154.6000 104.0000 155.3000 104.4000 ;
	    RECT 156.1000 104.5000 156.5000 104.6000 ;
	    RECT 156.9000 104.5000 157.2000 105.1000 ;
	    RECT 156.1000 104.2000 157.2000 104.5000 ;
	    RECT 157.5000 104.5000 160.2000 104.8000 ;
	    RECT 157.5000 104.4000 157.9000 104.5000 ;
	    RECT 159.8000 104.4000 160.2000 104.5000 ;
	    RECT 156.7000 103.7000 157.1000 103.8000 ;
	    RECT 158.1000 103.7000 158.5000 103.8000 ;
	    RECT 155.0000 103.1000 155.4000 103.5000 ;
	    RECT 156.7000 103.4000 158.5000 103.7000 ;
	    RECT 157.1000 103.1000 157.4000 103.4000 ;
	    RECT 159.8000 103.1000 160.2000 103.5000 ;
	    RECT 154.7000 101.1000 155.3000 103.1000 ;
	    RECT 157.0000 101.1000 157.4000 103.1000 ;
	    RECT 159.2000 102.8000 160.2000 103.1000 ;
	    RECT 159.2000 101.1000 159.6000 102.8000 ;
	    RECT 161.4000 101.1000 161.8000 105.3000 ;
	    RECT 162.2000 105.5000 165.0000 105.6000 ;
	    RECT 162.2000 105.4000 165.1000 105.5000 ;
	    RECT 162.2000 105.3000 167.1000 105.4000 ;
	    RECT 162.2000 101.1000 162.6000 105.3000 ;
	    RECT 164.7000 105.1000 167.1000 105.3000 ;
	    RECT 163.8000 104.5000 166.5000 104.8000 ;
	    RECT 163.8000 104.4000 164.2000 104.5000 ;
	    RECT 166.1000 104.4000 166.5000 104.5000 ;
	    RECT 166.8000 104.5000 167.1000 105.1000 ;
	    RECT 167.8000 105.2000 168.1000 106.8000 ;
	    RECT 168.6000 106.4000 169.0000 106.5000 ;
	    RECT 168.6000 106.1000 170.5000 106.4000 ;
	    RECT 170.1000 106.0000 170.5000 106.1000 ;
	    RECT 169.3000 105.7000 169.7000 105.8000 ;
	    RECT 171.0000 105.7000 171.4000 107.4000 ;
	    RECT 169.3000 105.4000 171.4000 105.7000 ;
	    RECT 167.8000 104.9000 169.0000 105.2000 ;
	    RECT 167.5000 104.5000 167.9000 104.6000 ;
	    RECT 166.8000 104.2000 167.9000 104.5000 ;
	    RECT 168.7000 104.4000 169.0000 104.9000 ;
	    RECT 168.7000 104.0000 169.4000 104.4000 ;
	    RECT 165.5000 103.7000 165.9000 103.8000 ;
	    RECT 166.9000 103.7000 167.3000 103.8000 ;
	    RECT 163.8000 103.1000 164.2000 103.5000 ;
	    RECT 165.5000 103.4000 167.3000 103.7000 ;
	    RECT 166.6000 103.1000 166.9000 103.4000 ;
	    RECT 168.6000 103.1000 169.0000 103.5000 ;
	    RECT 163.8000 102.8000 164.8000 103.1000 ;
	    RECT 164.4000 101.1000 164.8000 102.8000 ;
	    RECT 166.6000 101.1000 167.0000 103.1000 ;
	    RECT 168.7000 101.1000 169.3000 103.1000 ;
	    RECT 171.0000 101.1000 171.4000 105.4000 ;
	    RECT 0.6000 96.2000 1.0000 99.9000 ;
	    RECT 0.6000 95.9000 1.7000 96.2000 ;
	    RECT 2.2000 95.9000 2.6000 99.9000 ;
	    RECT 1.4000 95.6000 1.7000 95.9000 ;
	    RECT 1.4000 95.2000 2.0000 95.6000 ;
	    RECT 1.4000 93.7000 1.7000 95.2000 ;
	    RECT 2.3000 94.8000 2.6000 95.9000 ;
	    RECT 0.6000 93.4000 1.7000 93.7000 ;
	    RECT 0.6000 91.1000 1.0000 93.4000 ;
	    RECT 2.2000 91.1000 2.6000 94.8000 ;
	    RECT 3.8000 96.1000 4.2000 99.9000 ;
	    RECT 4.6000 96.1000 5.0000 96.6000 ;
	    RECT 3.8000 95.8000 5.0000 96.1000 ;
	    RECT 3.8000 91.1000 4.2000 95.8000 ;
	    RECT 5.4000 93.1000 5.8000 99.9000 ;
	    RECT 7.0000 95.6000 7.4000 99.9000 ;
	    RECT 9.1000 96.2000 9.5000 99.9000 ;
	    RECT 10.2000 97.9000 10.6000 99.9000 ;
	    RECT 10.3000 97.8000 10.6000 97.9000 ;
	    RECT 11.8000 97.9000 12.2000 99.9000 ;
	    RECT 11.8000 97.8000 12.1000 97.9000 ;
	    RECT 10.3000 97.5000 12.1000 97.8000 ;
	    RECT 10.3000 96.2000 10.6000 97.5000 ;
	    RECT 11.0000 96.4000 11.4000 97.2000 ;
	    RECT 9.1000 95.9000 9.8000 96.2000 ;
	    RECT 7.0000 95.4000 9.0000 95.6000 ;
	    RECT 7.0000 95.3000 9.1000 95.4000 ;
	    RECT 8.7000 95.0000 9.1000 95.3000 ;
	    RECT 9.5000 95.2000 9.8000 95.9000 ;
	    RECT 10.2000 95.8000 10.6000 96.2000 ;
	    RECT 8.0000 94.2000 8.4000 94.6000 ;
	    RECT 6.2000 94.1000 6.6000 94.2000 ;
	    RECT 7.8000 94.1000 8.3000 94.2000 ;
	    RECT 6.2000 93.8000 8.3000 94.1000 ;
	    RECT 6.2000 93.4000 6.6000 93.8000 ;
	    RECT 8.8000 93.5000 9.1000 95.0000 ;
	    RECT 9.4000 94.8000 9.8000 95.2000 ;
	    RECT 9.5000 94.2000 9.8000 94.8000 ;
	    RECT 9.4000 93.8000 9.8000 94.2000 ;
	    RECT 10.3000 94.2000 10.6000 95.8000 ;
	    RECT 12.6000 95.4000 13.0000 96.2000 ;
	    RECT 13.4000 95.6000 13.8000 99.9000 ;
	    RECT 15.5000 96.2000 15.9000 99.9000 ;
	    RECT 16.6000 97.1000 17.0000 97.2000 ;
	    RECT 17.4000 97.1000 17.8000 99.9000 ;
	    RECT 16.6000 96.8000 17.8000 97.1000 ;
	    RECT 15.5000 95.9000 16.2000 96.2000 ;
	    RECT 13.4000 95.4000 15.4000 95.6000 ;
	    RECT 13.4000 95.3000 15.5000 95.4000 ;
	    RECT 11.4000 94.8000 12.2000 95.2000 ;
	    RECT 15.1000 95.0000 15.5000 95.3000 ;
	    RECT 15.9000 95.2000 16.2000 95.9000 ;
	    RECT 10.3000 94.1000 11.1000 94.2000 ;
	    RECT 10.3000 93.9000 11.2000 94.1000 ;
	    RECT 4.9000 92.8000 5.8000 93.1000 ;
	    RECT 7.9000 93.2000 9.1000 93.5000 ;
	    RECT 4.9000 91.1000 5.3000 92.8000 ;
	    RECT 7.9000 92.1000 8.2000 93.2000 ;
	    RECT 9.5000 93.1000 9.8000 93.8000 ;
	    RECT 7.8000 91.1000 8.2000 92.1000 ;
	    RECT 9.4000 91.1000 9.8000 93.1000 ;
	    RECT 10.8000 92.1000 11.2000 93.9000 ;
	    RECT 15.2000 93.5000 15.5000 95.0000 ;
	    RECT 15.8000 94.8000 16.2000 95.2000 ;
	    RECT 15.9000 94.2000 16.2000 94.8000 ;
	    RECT 15.8000 93.8000 16.2000 94.2000 ;
	    RECT 14.3000 93.2000 15.5000 93.5000 ;
	    RECT 13.4000 92.4000 13.8000 93.2000 ;
	    RECT 11.8000 92.1000 12.2000 92.2000 ;
	    RECT 14.3000 92.1000 14.6000 93.2000 ;
	    RECT 15.9000 93.1000 16.2000 93.8000 ;
	    RECT 16.6000 93.4000 17.0000 94.2000 ;
	    RECT 10.8000 91.8000 12.2000 92.1000 ;
	    RECT 10.8000 91.1000 11.2000 91.8000 ;
	    RECT 14.2000 91.1000 14.6000 92.1000 ;
	    RECT 15.8000 91.1000 16.2000 93.1000 ;
	    RECT 17.4000 93.1000 17.8000 96.8000 ;
	    RECT 18.2000 96.1000 18.6000 96.6000 ;
	    RECT 19.8000 96.1000 20.2000 99.9000 ;
	    RECT 20.6000 97.9000 21.0000 99.9000 ;
	    RECT 20.7000 97.8000 21.0000 97.9000 ;
	    RECT 22.2000 97.9000 22.6000 99.9000 ;
	    RECT 22.2000 97.8000 22.5000 97.9000 ;
	    RECT 20.7000 97.5000 22.5000 97.8000 ;
	    RECT 20.7000 96.2000 21.0000 97.5000 ;
	    RECT 21.4000 96.4000 21.8000 97.2000 ;
	    RECT 23.8000 96.2000 24.2000 99.9000 ;
	    RECT 18.2000 95.8000 20.2000 96.1000 ;
	    RECT 20.6000 95.8000 21.0000 96.2000 ;
	    RECT 17.4000 92.8000 18.3000 93.1000 ;
	    RECT 17.9000 91.1000 18.3000 92.8000 ;
	    RECT 19.8000 91.1000 20.2000 95.8000 ;
	    RECT 20.7000 94.2000 21.0000 95.8000 ;
	    RECT 23.0000 95.4000 23.4000 96.2000 ;
	    RECT 23.8000 95.9000 24.9000 96.2000 ;
	    RECT 25.4000 95.9000 25.8000 99.9000 ;
	    RECT 27.0000 97.9000 27.4000 99.9000 ;
	    RECT 27.1000 97.8000 27.4000 97.9000 ;
	    RECT 28.6000 97.9000 29.0000 99.9000 ;
	    RECT 28.6000 97.8000 28.9000 97.9000 ;
	    RECT 30.2000 97.8000 30.6000 99.9000 ;
	    RECT 31.8000 97.9000 32.2000 99.9000 ;
	    RECT 31.8000 97.8000 32.1000 97.9000 ;
	    RECT 27.1000 97.5000 28.9000 97.8000 ;
	    RECT 30.3000 97.5000 32.1000 97.8000 ;
	    RECT 27.8000 96.4000 28.2000 97.2000 ;
	    RECT 28.6000 96.2000 28.9000 97.5000 ;
	    RECT 31.0000 96.4000 31.4000 97.2000 ;
	    RECT 31.8000 96.2000 32.1000 97.5000 ;
	    RECT 32.9000 96.2000 33.3000 99.9000 ;
	    RECT 24.6000 95.6000 24.9000 95.9000 ;
	    RECT 24.6000 95.2000 25.2000 95.6000 ;
	    RECT 21.8000 94.8000 22.6000 95.2000 ;
	    RECT 20.7000 94.1000 21.5000 94.2000 ;
	    RECT 20.7000 93.9000 21.6000 94.1000 ;
	    RECT 21.2000 91.1000 21.6000 93.9000 ;
	    RECT 24.6000 93.7000 24.9000 95.2000 ;
	    RECT 25.5000 94.8000 25.8000 95.9000 ;
	    RECT 26.2000 95.4000 26.6000 96.2000 ;
	    RECT 28.6000 95.8000 29.0000 96.2000 ;
	    RECT 31.8000 95.8000 32.2000 96.2000 ;
	    RECT 32.6000 95.9000 33.3000 96.2000 ;
	    RECT 28.6000 95.2000 28.9000 95.8000 ;
	    RECT 27.0000 94.8000 27.8000 95.2000 ;
	    RECT 28.6000 94.8000 29.0000 95.2000 ;
	    RECT 30.2000 94.8000 31.0000 95.2000 ;
	    RECT 23.8000 93.4000 24.9000 93.7000 ;
	    RECT 23.8000 91.1000 24.2000 93.4000 ;
	    RECT 25.4000 91.1000 25.8000 94.8000 ;
	    RECT 28.6000 94.2000 28.9000 94.8000 ;
	    RECT 31.8000 94.2000 32.1000 95.8000 ;
	    RECT 28.1000 94.1000 28.9000 94.2000 ;
	    RECT 31.3000 94.1000 32.1000 94.2000 ;
	    RECT 28.0000 93.9000 28.9000 94.1000 ;
	    RECT 31.2000 93.9000 32.1000 94.1000 ;
	    RECT 32.6000 95.2000 32.9000 95.9000 ;
	    RECT 35.0000 95.6000 35.4000 99.9000 ;
	    RECT 35.8000 97.9000 36.2000 99.9000 ;
	    RECT 35.9000 97.8000 36.2000 97.9000 ;
	    RECT 37.4000 97.9000 37.8000 99.9000 ;
	    RECT 37.4000 97.8000 37.7000 97.9000 ;
	    RECT 35.9000 97.5000 37.7000 97.8000 ;
	    RECT 35.9000 96.2000 36.2000 97.5000 ;
	    RECT 36.6000 96.4000 37.0000 97.2000 ;
	    RECT 35.8000 95.8000 36.2000 96.2000 ;
	    RECT 33.4000 95.4000 35.4000 95.6000 ;
	    RECT 33.3000 95.3000 35.4000 95.4000 ;
	    RECT 32.6000 94.8000 33.0000 95.2000 ;
	    RECT 33.3000 95.0000 33.7000 95.3000 ;
	    RECT 28.0000 91.1000 28.4000 93.9000 ;
	    RECT 31.2000 91.1000 31.6000 93.9000 ;
	    RECT 32.6000 93.1000 32.9000 94.8000 ;
	    RECT 33.3000 93.5000 33.6000 95.0000 ;
	    RECT 35.9000 94.2000 36.2000 95.8000 ;
	    RECT 38.2000 95.4000 38.6000 96.2000 ;
	    RECT 39.8000 96.1000 40.2000 99.9000 ;
	    RECT 41.4000 97.1000 41.8000 99.9000 ;
	    RECT 41.4000 96.8000 42.5000 97.1000 ;
	    RECT 40.6000 96.1000 41.0000 96.6000 ;
	    RECT 39.8000 95.8000 41.0000 96.1000 ;
	    RECT 37.0000 94.8000 37.8000 95.2000 ;
	    RECT 35.9000 94.1000 36.7000 94.2000 ;
	    RECT 35.9000 93.9000 37.7000 94.1000 ;
	    RECT 36.4000 93.8000 37.7000 93.9000 ;
	    RECT 33.3000 93.2000 34.5000 93.5000 ;
	    RECT 32.6000 91.1000 33.0000 93.1000 ;
	    RECT 34.2000 92.1000 34.5000 93.2000 ;
	    RECT 35.0000 92.4000 35.4000 93.2000 ;
	    RECT 34.2000 91.1000 34.6000 92.1000 ;
	    RECT 36.4000 91.1000 36.8000 93.8000 ;
	    RECT 37.4000 93.2000 37.7000 93.8000 ;
	    RECT 37.4000 92.8000 37.8000 93.2000 ;
	    RECT 39.8000 91.1000 40.2000 95.8000 ;
	    RECT 41.4000 93.1000 41.8000 96.8000 ;
	    RECT 42.2000 96.2000 42.5000 96.8000 ;
	    RECT 42.2000 95.8000 42.6000 96.2000 ;
	    RECT 43.0000 95.6000 43.4000 99.9000 ;
	    RECT 45.1000 96.2000 45.5000 99.9000 ;
	    RECT 46.2000 97.9000 46.6000 99.9000 ;
	    RECT 46.3000 97.8000 46.6000 97.9000 ;
	    RECT 47.8000 97.9000 48.2000 99.9000 ;
	    RECT 47.8000 97.8000 48.1000 97.9000 ;
	    RECT 46.3000 97.5000 48.1000 97.8000 ;
	    RECT 46.3000 96.2000 46.6000 97.5000 ;
	    RECT 47.0000 96.4000 47.4000 97.2000 ;
	    RECT 45.1000 95.9000 45.8000 96.2000 ;
	    RECT 43.0000 95.4000 45.0000 95.6000 ;
	    RECT 43.0000 95.3000 45.1000 95.4000 ;
	    RECT 44.7000 95.0000 45.1000 95.3000 ;
	    RECT 45.5000 95.2000 45.8000 95.9000 ;
	    RECT 46.2000 95.8000 46.6000 96.2000 ;
	    RECT 44.0000 94.2000 44.4000 94.6000 ;
	    RECT 42.2000 94.1000 42.6000 94.2000 ;
	    RECT 43.0000 94.1000 43.4000 94.2000 ;
	    RECT 42.2000 93.8000 43.4000 94.1000 ;
	    RECT 43.8000 93.8000 44.3000 94.2000 ;
	    RECT 42.2000 93.4000 42.6000 93.8000 ;
	    RECT 44.8000 93.5000 45.1000 95.0000 ;
	    RECT 45.4000 94.8000 45.8000 95.2000 ;
	    RECT 40.9000 92.8000 41.8000 93.1000 ;
	    RECT 43.9000 93.2000 45.1000 93.5000 ;
	    RECT 40.9000 91.1000 41.3000 92.8000 ;
	    RECT 43.9000 92.1000 44.2000 93.2000 ;
	    RECT 45.5000 93.1000 45.8000 94.8000 ;
	    RECT 46.3000 94.2000 46.6000 95.8000 ;
	    RECT 48.6000 95.4000 49.0000 96.2000 ;
	    RECT 50.2000 96.1000 50.6000 99.9000 ;
	    RECT 51.8000 97.1000 52.2000 99.9000 ;
	    RECT 51.8000 96.8000 52.9000 97.1000 ;
	    RECT 51.0000 96.1000 51.4000 96.6000 ;
	    RECT 50.2000 95.8000 51.4000 96.1000 ;
	    RECT 47.4000 94.8000 48.2000 95.2000 ;
	    RECT 46.3000 94.1000 47.1000 94.2000 ;
	    RECT 46.3000 93.9000 47.2000 94.1000 ;
	    RECT 43.8000 91.1000 44.2000 92.1000 ;
	    RECT 45.4000 91.1000 45.8000 93.1000 ;
	    RECT 46.8000 91.1000 47.2000 93.9000 ;
	    RECT 50.2000 91.1000 50.6000 95.8000 ;
	    RECT 51.8000 93.1000 52.2000 96.8000 ;
	    RECT 52.6000 96.2000 52.9000 96.8000 ;
	    RECT 52.6000 95.8000 53.0000 96.2000 ;
	    RECT 53.4000 95.6000 53.8000 99.9000 ;
	    RECT 55.5000 96.2000 55.9000 99.9000 ;
	    RECT 57.4000 97.9000 57.8000 99.9000 ;
	    RECT 57.5000 97.8000 57.8000 97.9000 ;
	    RECT 59.0000 97.9000 59.4000 99.9000 ;
	    RECT 59.8000 99.1000 60.2000 99.2000 ;
	    RECT 61.4000 99.1000 61.8000 99.9000 ;
	    RECT 59.8000 98.8000 61.8000 99.1000 ;
	    RECT 59.0000 97.8000 59.3000 97.9000 ;
	    RECT 57.5000 97.5000 59.3000 97.8000 ;
	    RECT 58.2000 96.4000 58.6000 97.2000 ;
	    RECT 59.0000 97.1000 59.3000 97.5000 ;
	    RECT 59.8000 97.1000 60.2000 97.2000 ;
	    RECT 59.0000 96.8000 60.2000 97.1000 ;
	    RECT 59.0000 96.2000 59.3000 96.8000 ;
	    RECT 55.5000 95.9000 56.2000 96.2000 ;
	    RECT 53.4000 95.4000 55.4000 95.6000 ;
	    RECT 53.4000 95.3000 55.5000 95.4000 ;
	    RECT 55.1000 95.0000 55.5000 95.3000 ;
	    RECT 55.9000 95.2000 56.2000 95.9000 ;
	    RECT 56.6000 95.4000 57.0000 96.2000 ;
	    RECT 59.0000 95.8000 59.4000 96.2000 ;
	    RECT 52.6000 94.1000 53.0000 94.2000 ;
	    RECT 52.6000 93.8000 53.7000 94.1000 ;
	    RECT 52.6000 93.4000 53.0000 93.8000 ;
	    RECT 51.3000 92.8000 52.2000 93.1000 ;
	    RECT 53.4000 93.2000 53.7000 93.8000 ;
	    RECT 55.2000 93.5000 55.5000 95.0000 ;
	    RECT 55.8000 94.8000 56.2000 95.2000 ;
	    RECT 57.4000 94.8000 58.2000 95.2000 ;
	    RECT 54.3000 93.2000 55.5000 93.5000 ;
	    RECT 51.3000 91.1000 51.7000 92.8000 ;
	    RECT 53.4000 92.4000 53.8000 93.2000 ;
	    RECT 54.3000 92.1000 54.6000 93.2000 ;
	    RECT 55.9000 93.1000 56.2000 94.8000 ;
	    RECT 59.0000 94.2000 59.3000 95.8000 ;
	    RECT 58.5000 94.1000 59.3000 94.2000 ;
	    RECT 54.2000 91.1000 54.6000 92.1000 ;
	    RECT 55.8000 91.1000 56.2000 93.1000 ;
	    RECT 58.4000 93.9000 59.3000 94.1000 ;
	    RECT 58.4000 91.1000 58.8000 93.9000 ;
	    RECT 61.4000 91.1000 61.8000 98.8000 ;
	    RECT 63.8000 96.1000 64.2000 99.9000 ;
	    RECT 64.6000 96.1000 65.0000 96.6000 ;
	    RECT 63.8000 95.8000 65.0000 96.1000 ;
	    RECT 65.4000 96.1000 65.8000 99.9000 ;
	    RECT 66.2000 96.8000 66.6000 97.2000 ;
	    RECT 66.2000 96.1000 66.5000 96.8000 ;
	    RECT 65.4000 95.8000 66.5000 96.1000 ;
	    RECT 63.8000 91.1000 64.2000 95.8000 ;
	    RECT 65.4000 93.1000 65.8000 95.8000 ;
	    RECT 67.0000 95.6000 67.4000 99.9000 ;
	    RECT 69.1000 96.2000 69.5000 99.9000 ;
	    RECT 70.2000 97.9000 70.6000 99.9000 ;
	    RECT 70.3000 97.8000 70.6000 97.9000 ;
	    RECT 71.8000 97.8000 72.2000 99.9000 ;
	    RECT 73.4000 97.9000 73.8000 99.9000 ;
	    RECT 73.5000 97.8000 73.8000 97.9000 ;
	    RECT 75.0000 97.9000 75.4000 99.9000 ;
	    RECT 75.0000 97.8000 75.3000 97.9000 ;
	    RECT 70.3000 97.5000 72.1000 97.8000 ;
	    RECT 73.5000 97.5000 75.3000 97.8000 ;
	    RECT 70.3000 96.2000 70.6000 97.5000 ;
	    RECT 71.0000 96.4000 71.4000 97.2000 ;
	    RECT 73.5000 96.2000 73.8000 97.5000 ;
	    RECT 74.2000 96.4000 74.6000 97.2000 ;
	    RECT 69.1000 95.9000 69.8000 96.2000 ;
	    RECT 67.0000 95.4000 69.0000 95.6000 ;
	    RECT 67.0000 95.3000 69.1000 95.4000 ;
	    RECT 68.7000 95.0000 69.1000 95.3000 ;
	    RECT 69.5000 95.2000 69.8000 95.9000 ;
	    RECT 70.2000 95.8000 70.6000 96.2000 ;
	    RECT 73.4000 95.8000 73.8000 96.2000 ;
	    RECT 75.0000 96.1000 75.4000 96.2000 ;
	    RECT 75.8000 96.1000 76.2000 96.2000 ;
	    RECT 75.0000 95.8000 76.2000 96.1000 ;
	    RECT 66.2000 94.1000 66.6000 94.2000 ;
	    RECT 66.2000 93.8000 67.3000 94.1000 ;
	    RECT 66.2000 93.4000 66.6000 93.8000 ;
	    RECT 64.9000 92.8000 65.8000 93.1000 ;
	    RECT 67.0000 93.2000 67.3000 93.8000 ;
	    RECT 68.8000 93.5000 69.1000 95.0000 ;
	    RECT 69.4000 94.8000 69.8000 95.2000 ;
	    RECT 69.5000 94.2000 69.8000 94.8000 ;
	    RECT 69.4000 93.8000 69.8000 94.2000 ;
	    RECT 70.3000 94.2000 70.6000 95.8000 ;
	    RECT 71.4000 94.8000 72.2000 95.2000 ;
	    RECT 73.5000 94.2000 73.8000 95.8000 ;
	    RECT 75.8000 95.4000 76.2000 95.8000 ;
	    RECT 76.6000 95.6000 77.0000 99.9000 ;
	    RECT 78.7000 96.2000 79.1000 99.9000 ;
	    RECT 78.7000 95.9000 79.4000 96.2000 ;
	    RECT 76.6000 95.4000 78.6000 95.6000 ;
	    RECT 76.6000 95.3000 78.7000 95.4000 ;
	    RECT 74.6000 94.8000 75.4000 95.2000 ;
	    RECT 78.3000 95.0000 78.7000 95.3000 ;
	    RECT 79.1000 95.2000 79.4000 95.9000 ;
	    RECT 79.8000 96.1000 80.2000 96.2000 ;
	    RECT 80.6000 96.1000 81.0000 99.9000 ;
	    RECT 82.2000 97.9000 82.6000 99.9000 ;
	    RECT 82.3000 97.8000 82.6000 97.9000 ;
	    RECT 83.8000 97.9000 84.2000 99.9000 ;
	    RECT 83.8000 97.8000 84.1000 97.9000 ;
	    RECT 82.3000 97.5000 84.1000 97.8000 ;
	    RECT 83.0000 96.4000 83.4000 97.2000 ;
	    RECT 83.8000 96.2000 84.1000 97.5000 ;
	    RECT 79.8000 95.8000 81.0000 96.1000 ;
	    RECT 70.3000 94.1000 71.1000 94.2000 ;
	    RECT 73.5000 94.1000 74.3000 94.2000 ;
	    RECT 70.3000 93.9000 71.2000 94.1000 ;
	    RECT 73.5000 93.9000 74.4000 94.1000 ;
	    RECT 67.9000 93.2000 69.1000 93.5000 ;
	    RECT 64.9000 91.1000 65.3000 92.8000 ;
	    RECT 67.0000 92.4000 67.4000 93.2000 ;
	    RECT 67.9000 92.1000 68.2000 93.2000 ;
	    RECT 69.5000 93.1000 69.8000 93.8000 ;
	    RECT 67.8000 91.1000 68.2000 92.1000 ;
	    RECT 69.4000 91.1000 69.8000 93.1000 ;
	    RECT 70.8000 91.1000 71.2000 93.9000 ;
	    RECT 74.0000 92.1000 74.4000 93.9000 ;
	    RECT 78.4000 93.5000 78.7000 95.0000 ;
	    RECT 79.0000 95.1000 79.4000 95.2000 ;
	    RECT 79.0000 94.8000 80.1000 95.1000 ;
	    RECT 77.5000 93.2000 78.7000 93.5000 ;
	    RECT 76.6000 92.4000 77.0000 93.2000 ;
	    RECT 75.0000 92.1000 75.4000 92.2000 ;
	    RECT 77.5000 92.1000 77.8000 93.2000 ;
	    RECT 79.1000 93.1000 79.4000 94.8000 ;
	    RECT 79.8000 94.2000 80.1000 94.8000 ;
	    RECT 79.8000 93.8000 80.2000 94.2000 ;
	    RECT 74.0000 91.8000 75.4000 92.1000 ;
	    RECT 74.0000 91.1000 74.4000 91.8000 ;
	    RECT 77.4000 91.1000 77.8000 92.1000 ;
	    RECT 79.0000 91.1000 79.4000 93.1000 ;
	    RECT 80.6000 91.1000 81.0000 95.8000 ;
	    RECT 81.4000 95.4000 81.8000 96.2000 ;
	    RECT 83.8000 95.8000 84.2000 96.2000 ;
	    RECT 84.6000 95.8000 85.0000 96.6000 ;
	    RECT 82.2000 94.8000 83.0000 95.2000 ;
	    RECT 83.8000 94.2000 84.1000 95.8000 ;
	    RECT 83.3000 94.1000 84.1000 94.2000 ;
	    RECT 83.2000 93.9000 84.1000 94.1000 ;
	    RECT 83.2000 91.1000 83.6000 93.9000 ;
	    RECT 85.4000 93.1000 85.8000 99.9000 ;
	    RECT 87.8000 97.9000 88.2000 99.9000 ;
	    RECT 87.9000 97.8000 88.2000 97.9000 ;
	    RECT 89.4000 97.9000 89.8000 99.9000 ;
	    RECT 91.0000 97.9000 91.4000 99.9000 ;
	    RECT 89.4000 97.8000 89.7000 97.9000 ;
	    RECT 87.9000 97.5000 89.7000 97.8000 ;
	    RECT 91.1000 97.8000 91.4000 97.9000 ;
	    RECT 92.6000 97.9000 93.0000 99.9000 ;
	    RECT 92.6000 97.8000 92.9000 97.9000 ;
	    RECT 91.1000 97.5000 92.9000 97.8000 ;
	    RECT 88.6000 96.4000 89.0000 97.2000 ;
	    RECT 89.4000 96.2000 89.7000 97.5000 ;
	    RECT 91.0000 97.1000 91.4000 97.2000 ;
	    RECT 91.8000 97.1000 92.2000 97.2000 ;
	    RECT 91.0000 96.8000 92.2000 97.1000 ;
	    RECT 91.8000 96.4000 92.2000 96.8000 ;
	    RECT 92.6000 96.2000 92.9000 97.5000 ;
	    RECT 89.4000 95.8000 89.8000 96.2000 ;
	    RECT 92.6000 95.8000 93.0000 96.2000 ;
	    RECT 87.8000 94.8000 88.6000 95.2000 ;
	    RECT 89.4000 94.2000 89.7000 95.8000 ;
	    RECT 91.0000 94.8000 92.2000 95.2000 ;
	    RECT 92.6000 94.2000 92.9000 95.8000 ;
	    RECT 93.4000 95.6000 93.8000 99.9000 ;
	    RECT 95.5000 96.2000 95.9000 99.9000 ;
	    RECT 96.6000 97.9000 97.0000 99.9000 ;
	    RECT 96.7000 97.8000 97.0000 97.9000 ;
	    RECT 98.2000 97.9000 98.6000 99.9000 ;
	    RECT 98.2000 97.8000 98.5000 97.9000 ;
	    RECT 96.7000 97.5000 98.5000 97.8000 ;
	    RECT 96.7000 96.2000 97.0000 97.5000 ;
	    RECT 97.4000 96.4000 97.8000 97.2000 ;
	    RECT 99.8000 96.2000 100.2000 99.9000 ;
	    RECT 101.4000 96.2000 101.8000 99.9000 ;
	    RECT 95.5000 95.9000 96.2000 96.2000 ;
	    RECT 93.4000 95.4000 95.4000 95.6000 ;
	    RECT 93.4000 95.3000 95.5000 95.4000 ;
	    RECT 95.1000 95.0000 95.5000 95.3000 ;
	    RECT 95.9000 95.2000 96.2000 95.9000 ;
	    RECT 96.6000 95.8000 97.0000 96.2000 ;
	    RECT 86.2000 93.4000 86.6000 94.2000 ;
	    RECT 88.9000 94.1000 89.7000 94.2000 ;
	    RECT 92.1000 94.1000 92.9000 94.2000 ;
	    RECT 88.8000 93.9000 89.7000 94.1000 ;
	    RECT 92.0000 93.9000 92.9000 94.1000 ;
	    RECT 84.9000 92.8000 85.8000 93.1000 ;
	    RECT 84.9000 91.1000 85.3000 92.8000 ;
	    RECT 88.8000 91.1000 89.2000 93.9000 ;
	    RECT 92.0000 91.1000 92.4000 93.9000 ;
	    RECT 95.2000 93.5000 95.5000 95.0000 ;
	    RECT 95.8000 94.8000 96.2000 95.2000 ;
	    RECT 94.3000 93.2000 95.5000 93.5000 ;
	    RECT 93.4000 92.4000 93.8000 93.2000 ;
	    RECT 94.3000 92.1000 94.6000 93.2000 ;
	    RECT 95.9000 93.1000 96.2000 94.8000 ;
	    RECT 96.7000 94.2000 97.0000 95.8000 ;
	    RECT 99.0000 95.4000 99.4000 96.2000 ;
	    RECT 99.8000 95.9000 101.8000 96.2000 ;
	    RECT 102.2000 95.9000 102.6000 99.9000 ;
	    RECT 103.0000 95.9000 103.4000 99.9000 ;
	    RECT 103.8000 96.2000 104.2000 99.9000 ;
	    RECT 105.4000 96.2000 105.8000 99.9000 ;
	    RECT 103.8000 95.9000 105.8000 96.2000 ;
	    RECT 106.2000 96.2000 106.6000 99.9000 ;
	    RECT 107.8000 96.2000 108.2000 99.9000 ;
	    RECT 106.2000 95.9000 108.2000 96.2000 ;
	    RECT 108.6000 95.9000 109.0000 99.9000 ;
	    RECT 109.4000 96.2000 109.8000 99.9000 ;
	    RECT 111.0000 96.2000 111.4000 99.9000 ;
	    RECT 109.4000 95.9000 111.4000 96.2000 ;
	    RECT 111.8000 95.9000 112.2000 99.9000 ;
	    RECT 114.2000 96.2000 114.6000 99.9000 ;
	    RECT 115.8000 96.2000 116.2000 99.9000 ;
	    RECT 114.2000 95.9000 116.2000 96.2000 ;
	    RECT 116.6000 95.9000 117.0000 99.9000 ;
	    RECT 100.2000 95.2000 100.6000 95.4000 ;
	    RECT 102.2000 95.2000 102.5000 95.9000 ;
	    RECT 103.1000 95.2000 103.4000 95.9000 ;
	    RECT 105.0000 95.2000 105.4000 95.4000 ;
	    RECT 106.6000 95.2000 107.0000 95.4000 ;
	    RECT 108.6000 95.2000 108.9000 95.9000 ;
	    RECT 109.8000 95.2000 110.2000 95.4000 ;
	    RECT 111.8000 95.2000 112.1000 95.9000 ;
	    RECT 114.6000 95.2000 115.0000 95.4000 ;
	    RECT 116.6000 95.2000 116.9000 95.9000 ;
	    RECT 117.4000 95.7000 117.8000 99.9000 ;
	    RECT 119.6000 98.2000 120.0000 99.9000 ;
	    RECT 119.0000 97.9000 120.0000 98.2000 ;
	    RECT 121.8000 97.9000 122.2000 99.9000 ;
	    RECT 123.9000 97.9000 124.5000 99.9000 ;
	    RECT 119.0000 97.5000 119.4000 97.9000 ;
	    RECT 121.8000 97.6000 122.1000 97.9000 ;
	    RECT 120.7000 97.3000 122.5000 97.6000 ;
	    RECT 123.8000 97.5000 124.2000 97.9000 ;
	    RECT 120.7000 97.2000 121.1000 97.3000 ;
	    RECT 122.1000 97.2000 122.5000 97.3000 ;
	    RECT 119.0000 96.5000 119.4000 96.6000 ;
	    RECT 121.3000 96.5000 121.7000 96.6000 ;
	    RECT 119.0000 96.2000 121.7000 96.5000 ;
	    RECT 122.0000 96.5000 123.1000 96.8000 ;
	    RECT 122.0000 95.9000 122.3000 96.5000 ;
	    RECT 122.7000 96.4000 123.1000 96.5000 ;
	    RECT 123.9000 96.6000 124.6000 97.0000 ;
	    RECT 123.9000 96.1000 124.2000 96.6000 ;
	    RECT 119.9000 95.7000 122.3000 95.9000 ;
	    RECT 117.4000 95.6000 122.3000 95.7000 ;
	    RECT 123.0000 95.8000 124.2000 96.1000 ;
	    RECT 117.4000 95.5000 120.3000 95.6000 ;
	    RECT 117.4000 95.4000 120.2000 95.5000 ;
	    RECT 97.8000 94.8000 98.6000 95.2000 ;
	    RECT 99.8000 94.9000 100.6000 95.2000 ;
	    RECT 101.4000 94.9000 102.6000 95.2000 ;
	    RECT 99.8000 94.8000 100.2000 94.9000 ;
	    RECT 96.7000 94.1000 97.5000 94.2000 ;
	    RECT 96.7000 93.9000 97.6000 94.1000 ;
	    RECT 94.2000 91.1000 94.6000 92.1000 ;
	    RECT 95.8000 91.1000 96.2000 93.1000 ;
	    RECT 97.2000 92.1000 97.6000 93.9000 ;
	    RECT 100.6000 93.8000 101.0000 94.6000 ;
	    RECT 101.4000 93.1000 101.7000 94.9000 ;
	    RECT 102.2000 94.8000 102.6000 94.9000 ;
	    RECT 103.0000 94.9000 104.2000 95.2000 ;
	    RECT 105.0000 94.9000 105.8000 95.2000 ;
	    RECT 103.0000 94.8000 103.4000 94.9000 ;
	    RECT 102.2000 94.2000 102.5000 94.8000 ;
	    RECT 102.2000 93.8000 102.6000 94.2000 ;
	    RECT 102.2000 93.1000 102.6000 93.2000 ;
	    RECT 103.0000 93.1000 103.4000 93.2000 ;
	    RECT 103.9000 93.1000 104.2000 94.9000 ;
	    RECT 105.4000 94.8000 105.8000 94.9000 ;
	    RECT 106.2000 94.9000 107.0000 95.2000 ;
	    RECT 107.8000 94.9000 109.0000 95.2000 ;
	    RECT 106.2000 94.8000 106.6000 94.9000 ;
	    RECT 104.6000 93.8000 105.0000 94.6000 ;
	    RECT 107.0000 93.8000 107.4000 94.6000 ;
	    RECT 98.2000 92.1000 98.6000 92.2000 ;
	    RECT 97.2000 91.8000 98.6000 92.1000 ;
	    RECT 97.2000 91.1000 97.6000 91.8000 ;
	    RECT 101.4000 91.1000 101.8000 93.1000 ;
	    RECT 102.2000 92.8000 103.4000 93.1000 ;
	    RECT 102.1000 92.4000 102.5000 92.8000 ;
	    RECT 103.1000 92.4000 103.5000 92.8000 ;
	    RECT 103.8000 91.1000 104.2000 93.1000 ;
	    RECT 107.8000 93.1000 108.1000 94.9000 ;
	    RECT 108.6000 94.8000 109.0000 94.9000 ;
	    RECT 109.4000 94.9000 110.2000 95.2000 ;
	    RECT 111.0000 94.9000 112.2000 95.2000 ;
	    RECT 109.4000 94.8000 109.8000 94.9000 ;
	    RECT 110.2000 93.8000 110.6000 94.6000 ;
	    RECT 107.8000 91.1000 108.2000 93.1000 ;
	    RECT 108.6000 92.8000 109.0000 93.2000 ;
	    RECT 111.0000 93.1000 111.3000 94.9000 ;
	    RECT 111.8000 94.8000 112.2000 94.9000 ;
	    RECT 114.2000 94.9000 115.0000 95.2000 ;
	    RECT 115.8000 94.9000 117.0000 95.2000 ;
	    RECT 120.6000 95.1000 121.0000 95.2000 ;
	    RECT 114.2000 94.8000 114.6000 94.9000 ;
	    RECT 115.0000 93.8000 115.4000 94.6000 ;
	    RECT 115.8000 94.1000 116.1000 94.9000 ;
	    RECT 116.6000 94.8000 117.0000 94.9000 ;
	    RECT 118.5000 94.8000 121.0000 95.1000 ;
	    RECT 118.5000 94.7000 118.9000 94.8000 ;
	    RECT 119.8000 94.7000 120.2000 94.8000 ;
	    RECT 119.3000 94.2000 119.7000 94.3000 ;
	    RECT 123.0000 94.2000 123.3000 95.8000 ;
	    RECT 126.2000 95.6000 126.6000 99.9000 ;
	    RECT 124.5000 95.3000 126.6000 95.6000 ;
	    RECT 124.5000 95.2000 124.9000 95.3000 ;
	    RECT 125.3000 94.9000 125.7000 95.0000 ;
	    RECT 123.8000 94.6000 125.7000 94.9000 ;
	    RECT 123.8000 94.5000 124.2000 94.6000 ;
	    RECT 116.6000 94.1000 117.0000 94.2000 ;
	    RECT 115.8000 93.8000 117.0000 94.1000 ;
	    RECT 117.8000 93.9000 123.3000 94.2000 ;
	    RECT 117.8000 93.8000 118.6000 93.9000 ;
	    RECT 111.8000 93.1000 112.2000 93.2000 ;
	    RECT 113.4000 93.1000 113.8000 93.2000 ;
	    RECT 108.5000 92.4000 108.9000 92.8000 ;
	    RECT 111.0000 91.1000 111.4000 93.1000 ;
	    RECT 111.8000 92.8000 113.8000 93.1000 ;
	    RECT 115.8000 93.1000 116.1000 93.8000 ;
	    RECT 111.7000 92.4000 112.1000 92.8000 ;
	    RECT 115.8000 91.1000 116.2000 93.1000 ;
	    RECT 116.6000 92.8000 117.0000 93.2000 ;
	    RECT 116.5000 92.4000 116.9000 92.8000 ;
	    RECT 117.4000 91.1000 117.8000 93.5000 ;
	    RECT 119.9000 92.8000 120.2000 93.9000 ;
	    RECT 122.7000 93.8000 123.1000 93.9000 ;
	    RECT 126.2000 93.6000 126.6000 95.3000 ;
	    RECT 124.7000 93.3000 126.6000 93.6000 ;
	    RECT 124.7000 93.2000 125.1000 93.3000 ;
	    RECT 119.0000 92.1000 119.4000 92.5000 ;
	    RECT 119.8000 92.4000 120.2000 92.8000 ;
	    RECT 120.7000 92.7000 121.1000 92.8000 ;
	    RECT 120.7000 92.4000 122.1000 92.7000 ;
	    RECT 121.8000 92.1000 122.1000 92.4000 ;
	    RECT 123.8000 92.1000 124.2000 92.5000 ;
	    RECT 119.0000 91.8000 120.0000 92.1000 ;
	    RECT 119.6000 91.1000 120.0000 91.8000 ;
	    RECT 121.8000 91.1000 122.2000 92.1000 ;
	    RECT 123.8000 91.8000 124.5000 92.1000 ;
	    RECT 123.9000 91.1000 124.5000 91.8000 ;
	    RECT 126.2000 91.1000 126.6000 93.3000 ;
	    RECT 127.0000 95.6000 127.4000 99.9000 ;
	    RECT 129.1000 97.9000 129.7000 99.9000 ;
	    RECT 131.4000 97.9000 131.8000 99.9000 ;
	    RECT 133.6000 98.2000 134.0000 99.9000 ;
	    RECT 133.6000 97.9000 134.6000 98.2000 ;
	    RECT 129.4000 97.5000 129.8000 97.9000 ;
	    RECT 131.5000 97.6000 131.8000 97.9000 ;
	    RECT 131.1000 97.3000 132.9000 97.6000 ;
	    RECT 134.2000 97.5000 134.6000 97.9000 ;
	    RECT 131.1000 97.2000 131.5000 97.3000 ;
	    RECT 132.5000 97.2000 132.9000 97.3000 ;
	    RECT 129.0000 96.6000 129.7000 97.0000 ;
	    RECT 129.4000 96.1000 129.7000 96.6000 ;
	    RECT 130.5000 96.5000 131.6000 96.8000 ;
	    RECT 130.5000 96.4000 130.9000 96.5000 ;
	    RECT 129.4000 95.8000 130.6000 96.1000 ;
	    RECT 127.0000 95.3000 129.1000 95.6000 ;
	    RECT 127.0000 93.6000 127.4000 95.3000 ;
	    RECT 128.7000 95.2000 129.1000 95.3000 ;
	    RECT 130.3000 95.2000 130.6000 95.8000 ;
	    RECT 131.3000 95.9000 131.6000 96.5000 ;
	    RECT 131.9000 96.5000 132.3000 96.6000 ;
	    RECT 134.2000 96.5000 134.6000 96.6000 ;
	    RECT 131.9000 96.2000 134.6000 96.5000 ;
	    RECT 131.3000 95.7000 133.7000 95.9000 ;
	    RECT 135.8000 95.7000 136.2000 99.9000 ;
	    RECT 136.6000 95.8000 137.0000 96.6000 ;
	    RECT 131.3000 95.6000 136.2000 95.7000 ;
	    RECT 133.3000 95.5000 136.2000 95.6000 ;
	    RECT 133.4000 95.4000 136.2000 95.5000 ;
	    RECT 127.9000 94.9000 128.3000 95.0000 ;
	    RECT 127.9000 94.6000 129.8000 94.9000 ;
	    RECT 130.2000 94.8000 130.6000 95.2000 ;
	    RECT 132.6000 95.1000 133.0000 95.2000 ;
	    RECT 132.6000 94.8000 135.1000 95.1000 ;
	    RECT 129.4000 94.5000 129.8000 94.6000 ;
	    RECT 130.3000 94.2000 130.6000 94.8000 ;
	    RECT 134.7000 94.7000 135.1000 94.8000 ;
	    RECT 133.9000 94.2000 134.3000 94.3000 ;
	    RECT 130.3000 93.9000 135.8000 94.2000 ;
	    RECT 130.5000 93.8000 130.9000 93.9000 ;
	    RECT 127.0000 93.3000 128.9000 93.6000 ;
	    RECT 127.0000 91.1000 127.4000 93.3000 ;
	    RECT 128.5000 93.2000 128.9000 93.3000 ;
	    RECT 133.4000 92.8000 133.7000 93.9000 ;
	    RECT 135.0000 93.8000 135.8000 93.9000 ;
	    RECT 132.5000 92.7000 132.9000 92.8000 ;
	    RECT 129.4000 92.1000 129.8000 92.5000 ;
	    RECT 131.5000 92.4000 132.9000 92.7000 ;
	    RECT 133.4000 92.4000 133.8000 92.8000 ;
	    RECT 131.5000 92.1000 131.8000 92.4000 ;
	    RECT 134.2000 92.1000 134.6000 92.5000 ;
	    RECT 129.1000 91.8000 129.8000 92.1000 ;
	    RECT 129.1000 91.1000 129.7000 91.8000 ;
	    RECT 131.4000 91.1000 131.8000 92.1000 ;
	    RECT 133.6000 91.8000 134.6000 92.1000 ;
	    RECT 133.6000 91.1000 134.0000 91.8000 ;
	    RECT 135.8000 91.1000 136.2000 93.5000 ;
	    RECT 137.4000 93.1000 137.8000 99.9000 ;
	    RECT 138.2000 93.4000 138.6000 94.2000 ;
	    RECT 136.9000 92.8000 137.8000 93.1000 ;
	    RECT 136.9000 91.1000 137.3000 92.8000 ;
	    RECT 139.0000 91.1000 139.4000 99.9000 ;
	    RECT 140.6000 96.2000 141.0000 99.9000 ;
	    RECT 140.6000 95.9000 141.7000 96.2000 ;
	    RECT 142.2000 95.9000 142.6000 99.9000 ;
	    RECT 141.4000 95.6000 141.7000 95.9000 ;
	    RECT 141.4000 95.2000 142.0000 95.6000 ;
	    RECT 141.4000 93.7000 141.7000 95.2000 ;
	    RECT 142.3000 94.8000 142.6000 95.9000 ;
	    RECT 140.6000 93.4000 141.7000 93.7000 ;
	    RECT 139.8000 92.4000 140.2000 93.2000 ;
	    RECT 140.6000 91.1000 141.0000 93.4000 ;
	    RECT 142.2000 91.1000 142.6000 94.8000 ;
	    RECT 143.0000 95.6000 143.4000 99.9000 ;
	    RECT 145.1000 97.9000 145.7000 99.9000 ;
	    RECT 147.4000 97.9000 147.8000 99.9000 ;
	    RECT 149.6000 98.2000 150.0000 99.9000 ;
	    RECT 149.6000 97.9000 150.6000 98.2000 ;
	    RECT 145.4000 97.5000 145.8000 97.9000 ;
	    RECT 147.5000 97.6000 147.8000 97.9000 ;
	    RECT 147.1000 97.3000 148.9000 97.6000 ;
	    RECT 150.2000 97.5000 150.6000 97.9000 ;
	    RECT 147.1000 97.2000 147.5000 97.3000 ;
	    RECT 148.5000 97.2000 148.9000 97.3000 ;
	    RECT 145.0000 96.6000 145.7000 97.0000 ;
	    RECT 145.4000 96.1000 145.7000 96.6000 ;
	    RECT 146.5000 96.5000 147.6000 96.8000 ;
	    RECT 146.5000 96.4000 146.9000 96.5000 ;
	    RECT 145.4000 95.8000 146.6000 96.1000 ;
	    RECT 143.0000 95.3000 145.1000 95.6000 ;
	    RECT 143.0000 93.6000 143.4000 95.3000 ;
	    RECT 144.7000 95.2000 145.1000 95.3000 ;
	    RECT 146.3000 95.2000 146.6000 95.8000 ;
	    RECT 147.3000 95.9000 147.6000 96.5000 ;
	    RECT 147.9000 96.5000 148.3000 96.6000 ;
	    RECT 150.2000 96.5000 150.6000 96.6000 ;
	    RECT 147.9000 96.2000 150.6000 96.5000 ;
	    RECT 147.3000 95.7000 149.7000 95.9000 ;
	    RECT 151.8000 95.7000 152.2000 99.9000 ;
	    RECT 147.3000 95.6000 152.2000 95.7000 ;
	    RECT 153.4000 95.6000 153.8000 99.9000 ;
	    RECT 155.0000 95.6000 155.4000 99.9000 ;
	    RECT 156.6000 95.6000 157.0000 99.9000 ;
	    RECT 158.2000 95.6000 158.6000 99.9000 ;
	    RECT 149.3000 95.5000 152.2000 95.6000 ;
	    RECT 149.4000 95.4000 152.2000 95.5000 ;
	    RECT 152.6000 95.2000 153.8000 95.6000 ;
	    RECT 154.3000 95.2000 155.4000 95.6000 ;
	    RECT 155.9000 95.2000 157.0000 95.6000 ;
	    RECT 157.7000 95.2000 158.6000 95.6000 ;
	    RECT 159.8000 95.7000 160.2000 99.9000 ;
	    RECT 162.0000 98.2000 162.4000 99.9000 ;
	    RECT 161.4000 97.9000 162.4000 98.2000 ;
	    RECT 164.2000 97.9000 164.6000 99.9000 ;
	    RECT 166.3000 97.9000 166.9000 99.9000 ;
	    RECT 161.4000 97.5000 161.8000 97.9000 ;
	    RECT 164.2000 97.6000 164.5000 97.9000 ;
	    RECT 163.1000 97.3000 164.9000 97.6000 ;
	    RECT 166.2000 97.5000 166.6000 97.9000 ;
	    RECT 163.1000 97.2000 163.5000 97.3000 ;
	    RECT 164.5000 97.2000 164.9000 97.3000 ;
	    RECT 161.4000 96.5000 161.8000 96.6000 ;
	    RECT 163.7000 96.5000 164.1000 96.6000 ;
	    RECT 161.4000 96.2000 164.1000 96.5000 ;
	    RECT 164.4000 96.5000 165.5000 96.8000 ;
	    RECT 164.4000 95.9000 164.7000 96.5000 ;
	    RECT 165.1000 96.4000 165.5000 96.5000 ;
	    RECT 166.3000 96.6000 167.0000 97.0000 ;
	    RECT 166.3000 96.1000 166.6000 96.6000 ;
	    RECT 162.3000 95.7000 164.7000 95.9000 ;
	    RECT 159.8000 95.6000 164.7000 95.7000 ;
	    RECT 165.4000 95.8000 166.6000 96.1000 ;
	    RECT 159.8000 95.5000 162.7000 95.6000 ;
	    RECT 159.8000 95.4000 162.6000 95.5000 ;
	    RECT 143.9000 94.9000 144.3000 95.0000 ;
	    RECT 143.9000 94.6000 145.8000 94.9000 ;
	    RECT 146.2000 94.8000 146.6000 95.2000 ;
	    RECT 148.6000 95.1000 149.0000 95.2000 ;
	    RECT 148.6000 94.8000 151.1000 95.1000 ;
	    RECT 145.4000 94.5000 145.8000 94.6000 ;
	    RECT 146.3000 94.2000 146.6000 94.8000 ;
	    RECT 150.7000 94.7000 151.1000 94.8000 ;
	    RECT 149.9000 94.2000 150.3000 94.3000 ;
	    RECT 146.3000 93.9000 151.8000 94.2000 ;
	    RECT 146.5000 93.8000 146.9000 93.9000 ;
	    RECT 143.0000 93.3000 144.9000 93.6000 ;
	    RECT 143.0000 91.1000 143.4000 93.3000 ;
	    RECT 144.5000 93.2000 144.9000 93.3000 ;
	    RECT 149.4000 92.8000 149.7000 93.9000 ;
	    RECT 151.0000 93.8000 151.8000 93.9000 ;
	    RECT 152.6000 93.8000 153.0000 95.2000 ;
	    RECT 154.3000 94.5000 154.7000 95.2000 ;
	    RECT 155.9000 94.5000 156.3000 95.2000 ;
	    RECT 157.7000 94.5000 158.1000 95.2000 ;
	    RECT 163.0000 95.1000 163.4000 95.2000 ;
	    RECT 164.6000 95.1000 165.0000 95.2000 ;
	    RECT 160.9000 94.8000 165.0000 95.1000 ;
	    RECT 160.9000 94.7000 161.3000 94.8000 ;
	    RECT 153.4000 94.1000 154.7000 94.5000 ;
	    RECT 155.1000 94.1000 156.3000 94.5000 ;
	    RECT 156.8000 94.1000 158.1000 94.5000 ;
	    RECT 161.7000 94.2000 162.1000 94.3000 ;
	    RECT 165.4000 94.2000 165.7000 95.8000 ;
	    RECT 168.6000 95.6000 169.0000 99.9000 ;
	    RECT 166.9000 95.3000 169.0000 95.6000 ;
	    RECT 166.9000 95.2000 167.3000 95.3000 ;
	    RECT 167.7000 94.9000 168.1000 95.0000 ;
	    RECT 166.2000 94.6000 168.1000 94.9000 ;
	    RECT 166.2000 94.5000 166.6000 94.6000 ;
	    RECT 154.3000 93.8000 154.7000 94.1000 ;
	    RECT 155.9000 93.8000 156.3000 94.1000 ;
	    RECT 157.7000 93.8000 158.1000 94.1000 ;
	    RECT 160.2000 93.9000 165.7000 94.2000 ;
	    RECT 160.2000 93.8000 161.0000 93.9000 ;
	    RECT 148.5000 92.7000 148.9000 92.8000 ;
	    RECT 145.4000 92.1000 145.8000 92.5000 ;
	    RECT 147.5000 92.4000 148.9000 92.7000 ;
	    RECT 149.4000 92.4000 149.8000 92.8000 ;
	    RECT 147.5000 92.1000 147.8000 92.4000 ;
	    RECT 150.2000 92.1000 150.6000 92.5000 ;
	    RECT 145.1000 91.8000 145.8000 92.1000 ;
	    RECT 145.1000 91.1000 145.7000 91.8000 ;
	    RECT 147.4000 91.1000 147.8000 92.1000 ;
	    RECT 149.6000 91.8000 150.6000 92.1000 ;
	    RECT 149.6000 91.1000 150.0000 91.8000 ;
	    RECT 151.8000 91.1000 152.2000 93.5000 ;
	    RECT 152.6000 93.4000 153.8000 93.8000 ;
	    RECT 154.3000 93.4000 155.4000 93.8000 ;
	    RECT 155.9000 93.4000 157.0000 93.8000 ;
	    RECT 157.7000 93.4000 158.6000 93.8000 ;
	    RECT 153.4000 91.1000 153.8000 93.4000 ;
	    RECT 155.0000 91.1000 155.4000 93.4000 ;
	    RECT 156.6000 91.1000 157.0000 93.4000 ;
	    RECT 158.2000 91.1000 158.6000 93.4000 ;
	    RECT 159.8000 91.1000 160.2000 93.5000 ;
	    RECT 162.3000 92.8000 162.6000 93.9000 ;
	    RECT 165.1000 93.8000 165.5000 93.9000 ;
	    RECT 168.6000 93.6000 169.0000 95.3000 ;
	    RECT 167.1000 93.3000 169.0000 93.6000 ;
	    RECT 167.1000 93.2000 167.5000 93.3000 ;
	    RECT 161.4000 92.1000 161.8000 92.5000 ;
	    RECT 162.2000 92.4000 162.6000 92.8000 ;
	    RECT 163.1000 92.7000 163.5000 92.8000 ;
	    RECT 163.1000 92.4000 164.5000 92.7000 ;
	    RECT 164.2000 92.1000 164.5000 92.4000 ;
	    RECT 166.2000 92.1000 166.6000 92.5000 ;
	    RECT 161.4000 91.8000 162.4000 92.1000 ;
	    RECT 162.0000 91.1000 162.4000 91.8000 ;
	    RECT 164.2000 91.1000 164.6000 92.1000 ;
	    RECT 166.2000 91.8000 166.9000 92.1000 ;
	    RECT 166.3000 91.1000 166.9000 91.8000 ;
	    RECT 168.6000 91.1000 169.0000 93.3000 ;
	    RECT 169.4000 95.9000 169.8000 99.9000 ;
	    RECT 171.0000 97.9000 171.4000 99.9000 ;
	    RECT 169.4000 95.2000 169.7000 95.9000 ;
	    RECT 171.0000 95.8000 171.3000 97.9000 ;
	    RECT 170.1000 95.5000 171.3000 95.8000 ;
	    RECT 169.4000 94.8000 169.8000 95.2000 ;
	    RECT 169.4000 93.1000 169.7000 94.8000 ;
	    RECT 170.1000 93.8000 170.4000 95.5000 ;
	    RECT 171.0000 94.8000 171.4000 95.2000 ;
	    RECT 171.0000 94.4000 171.3000 94.8000 ;
	    RECT 170.8000 94.1000 171.3000 94.4000 ;
	    RECT 170.8000 94.0000 171.2000 94.1000 ;
	    RECT 171.8000 93.8000 172.2000 94.6000 ;
	    RECT 170.0000 93.7000 170.4000 93.8000 ;
	    RECT 170.0000 93.5000 171.5000 93.7000 ;
	    RECT 170.0000 93.4000 172.1000 93.5000 ;
	    RECT 171.2000 93.2000 172.1000 93.4000 ;
	    RECT 171.8000 93.1000 172.1000 93.2000 ;
	    RECT 169.4000 92.6000 170.1000 93.1000 ;
	    RECT 169.7000 92.2000 170.1000 92.6000 ;
	    RECT 169.4000 91.8000 170.1000 92.2000 ;
	    RECT 169.7000 91.1000 170.1000 91.8000 ;
	    RECT 171.8000 91.1000 172.2000 93.1000 ;
	    RECT 0.6000 84.1000 1.0000 84.2000 ;
	    RECT 1.4000 84.1000 1.8000 89.9000 ;
	    RECT 3.5000 88.2000 3.9000 89.9000 ;
	    RECT 3.0000 87.9000 3.9000 88.2000 ;
	    RECT 2.2000 86.8000 2.6000 87.6000 ;
	    RECT 0.6000 83.8000 1.8000 84.1000 ;
	    RECT 1.4000 81.1000 1.8000 83.8000 ;
	    RECT 3.0000 81.1000 3.4000 87.9000 ;
	    RECT 3.8000 85.1000 4.2000 85.2000 ;
	    RECT 4.6000 85.1000 5.0000 89.9000 ;
	    RECT 7.0000 88.9000 7.4000 89.9000 ;
	    RECT 6.2000 87.8000 6.6000 88.6000 ;
	    RECT 7.1000 87.8000 7.4000 88.9000 ;
	    RECT 8.6000 87.9000 9.0000 89.9000 ;
	    RECT 7.1000 87.5000 8.3000 87.8000 ;
	    RECT 8.0000 86.0000 8.3000 87.5000 ;
	    RECT 8.7000 87.2000 9.0000 87.9000 ;
	    RECT 8.6000 86.8000 9.0000 87.2000 ;
	    RECT 10.0000 87.1000 10.4000 89.9000 ;
	    RECT 13.2000 87.1000 13.6000 89.9000 ;
	    RECT 8.7000 86.2000 9.0000 86.8000 ;
	    RECT 7.9000 85.7000 8.3000 86.0000 ;
	    RECT 8.6000 85.8000 9.0000 86.2000 ;
	    RECT 3.8000 84.8000 5.0000 85.1000 ;
	    RECT 3.8000 84.4000 4.2000 84.8000 ;
	    RECT 4.6000 81.1000 5.0000 84.8000 ;
	    RECT 6.2000 85.6000 8.3000 85.7000 ;
	    RECT 6.2000 85.4000 8.2000 85.6000 ;
	    RECT 6.2000 81.1000 6.6000 85.4000 ;
	    RECT 8.7000 85.1000 9.0000 85.8000 ;
	    RECT 9.5000 86.9000 10.4000 87.1000 ;
	    RECT 12.7000 86.9000 13.6000 87.1000 ;
	    RECT 9.5000 86.8000 10.3000 86.9000 ;
	    RECT 12.7000 86.8000 13.5000 86.9000 ;
	    RECT 9.5000 85.2000 9.8000 86.8000 ;
	    RECT 10.6000 85.8000 11.4000 86.2000 ;
	    RECT 12.7000 85.2000 13.0000 86.8000 ;
	    RECT 13.8000 85.8000 14.6000 86.2000 ;
	    RECT 8.3000 84.8000 9.0000 85.1000 ;
	    RECT 9.4000 84.8000 9.8000 85.2000 ;
	    RECT 12.6000 84.8000 13.0000 85.2000 ;
	    RECT 15.0000 84.8000 15.4000 85.6000 ;
	    RECT 16.6000 85.1000 17.0000 89.9000 ;
	    RECT 18.7000 88.2000 19.1000 89.9000 ;
	    RECT 20.6000 88.9000 21.0000 89.9000 ;
	    RECT 18.2000 87.9000 19.1000 88.2000 ;
	    RECT 17.4000 86.8000 17.8000 87.6000 ;
	    RECT 18.2000 87.1000 18.6000 87.9000 ;
	    RECT 19.8000 87.8000 20.2000 88.6000 ;
	    RECT 20.7000 87.8000 21.0000 88.9000 ;
	    RECT 22.2000 87.9000 22.6000 89.9000 ;
	    RECT 20.7000 87.5000 21.9000 87.8000 ;
	    RECT 19.0000 87.1000 19.4000 87.2000 ;
	    RECT 18.2000 86.8000 19.4000 87.1000 ;
	    RECT 17.4000 85.8000 17.8000 86.2000 ;
	    RECT 17.4000 85.1000 17.7000 85.8000 ;
	    RECT 16.6000 84.8000 17.7000 85.1000 ;
	    RECT 8.3000 81.1000 8.7000 84.8000 ;
	    RECT 9.5000 83.5000 9.8000 84.8000 ;
	    RECT 10.2000 83.8000 10.6000 84.6000 ;
	    RECT 12.7000 83.5000 13.0000 84.8000 ;
	    RECT 13.4000 83.8000 13.8000 84.6000 ;
	    RECT 9.5000 83.2000 11.3000 83.5000 ;
	    RECT 9.5000 83.1000 9.8000 83.2000 ;
	    RECT 9.4000 81.1000 9.8000 83.1000 ;
	    RECT 11.0000 83.1000 11.3000 83.2000 ;
	    RECT 12.7000 83.2000 14.5000 83.5000 ;
	    RECT 12.7000 83.1000 13.0000 83.2000 ;
	    RECT 11.0000 81.1000 11.4000 83.1000 ;
	    RECT 12.6000 81.1000 13.0000 83.1000 ;
	    RECT 14.2000 83.1000 14.5000 83.2000 ;
	    RECT 14.2000 81.1000 14.6000 83.1000 ;
	    RECT 16.6000 81.1000 17.0000 84.8000 ;
	    RECT 18.2000 81.1000 18.6000 86.8000 ;
	    RECT 21.6000 86.0000 21.9000 87.5000 ;
	    RECT 22.3000 86.2000 22.6000 87.9000 ;
	    RECT 24.8000 87.2000 25.2000 89.9000 ;
	    RECT 24.6000 87.1000 25.2000 87.2000 ;
	    RECT 28.0000 87.1000 28.4000 89.9000 ;
	    RECT 30.0000 88.1000 30.4000 89.9000 ;
	    RECT 32.9000 89.2000 33.3000 89.9000 ;
	    RECT 32.6000 88.8000 33.3000 89.2000 ;
	    RECT 32.9000 88.2000 33.3000 88.8000 ;
	    RECT 30.0000 87.8000 31.3000 88.1000 ;
	    RECT 32.9000 87.9000 33.8000 88.2000 ;
	    RECT 30.0000 87.1000 30.4000 87.8000 ;
	    RECT 24.6000 86.8000 25.7000 87.1000 ;
	    RECT 28.0000 86.9000 28.9000 87.1000 ;
	    RECT 28.1000 86.8000 28.9000 86.9000 ;
	    RECT 21.5000 85.7000 21.9000 86.0000 ;
	    RECT 22.2000 85.8000 22.6000 86.2000 ;
	    RECT 23.8000 85.8000 24.6000 86.2000 ;
	    RECT 19.8000 85.6000 21.9000 85.7000 ;
	    RECT 19.8000 85.4000 21.8000 85.6000 ;
	    RECT 19.0000 84.4000 19.4000 85.2000 ;
	    RECT 19.8000 81.1000 20.2000 85.4000 ;
	    RECT 22.3000 85.1000 22.6000 85.8000 ;
	    RECT 21.9000 84.8000 22.6000 85.1000 ;
	    RECT 23.0000 84.8000 23.4000 85.6000 ;
	    RECT 25.4000 85.2000 25.7000 86.8000 ;
	    RECT 27.0000 85.8000 27.8000 86.2000 ;
	    RECT 28.6000 85.2000 28.9000 86.8000 ;
	    RECT 29.5000 86.9000 30.4000 87.1000 ;
	    RECT 31.0000 87.2000 31.3000 87.8000 ;
	    RECT 29.5000 86.8000 30.3000 86.9000 ;
	    RECT 31.0000 86.8000 31.4000 87.2000 ;
	    RECT 29.5000 85.2000 29.8000 86.8000 ;
	    RECT 30.6000 85.8000 31.4000 86.2000 ;
	    RECT 25.4000 84.8000 25.8000 85.2000 ;
	    RECT 28.6000 84.8000 29.0000 85.2000 ;
	    RECT 29.4000 84.8000 29.8000 85.2000 ;
	    RECT 31.8000 84.8000 32.2000 85.6000 ;
	    RECT 21.9000 81.1000 22.3000 84.8000 ;
	    RECT 24.6000 83.8000 25.0000 84.6000 ;
	    RECT 25.4000 83.5000 25.7000 84.8000 ;
	    RECT 27.8000 83.8000 28.2000 84.6000 ;
	    RECT 28.6000 83.5000 28.9000 84.8000 ;
	    RECT 23.9000 83.2000 25.7000 83.5000 ;
	    RECT 27.1000 83.2000 28.9000 83.5000 ;
	    RECT 23.9000 83.1000 24.2000 83.2000 ;
	    RECT 23.8000 81.1000 24.2000 83.1000 ;
	    RECT 25.4000 83.1000 25.7000 83.2000 ;
	    RECT 25.4000 81.1000 25.8000 83.1000 ;
	    RECT 27.0000 81.1000 27.4000 83.2000 ;
	    RECT 28.6000 83.1000 28.9000 83.2000 ;
	    RECT 29.5000 83.5000 29.8000 84.8000 ;
	    RECT 30.2000 83.8000 30.6000 84.6000 ;
	    RECT 32.6000 84.4000 33.0000 85.2000 ;
	    RECT 29.5000 83.2000 31.3000 83.5000 ;
	    RECT 29.5000 83.1000 29.8000 83.2000 ;
	    RECT 28.6000 81.1000 29.0000 83.1000 ;
	    RECT 29.4000 81.1000 29.8000 83.1000 ;
	    RECT 31.0000 83.1000 31.3000 83.2000 ;
	    RECT 31.0000 81.1000 31.4000 83.1000 ;
	    RECT 33.4000 81.1000 33.8000 87.9000 ;
	    RECT 35.0000 87.9000 35.4000 89.9000 ;
	    RECT 36.6000 88.9000 37.0000 89.9000 ;
	    RECT 34.2000 86.8000 34.6000 87.6000 ;
	    RECT 35.0000 86.2000 35.3000 87.9000 ;
	    RECT 36.6000 87.8000 36.9000 88.9000 ;
	    RECT 37.4000 87.8000 37.8000 88.6000 ;
	    RECT 39.5000 88.2000 39.9000 89.9000 ;
	    RECT 39.0000 87.9000 39.9000 88.2000 ;
	    RECT 35.7000 87.5000 36.9000 87.8000 ;
	    RECT 35.0000 86.1000 35.4000 86.2000 ;
	    RECT 34.2000 85.8000 35.4000 86.1000 ;
	    RECT 35.7000 86.0000 36.0000 87.5000 ;
	    RECT 34.2000 85.2000 34.5000 85.8000 ;
	    RECT 34.2000 84.8000 34.6000 85.2000 ;
	    RECT 35.0000 85.1000 35.3000 85.8000 ;
	    RECT 35.7000 85.7000 36.1000 86.0000 ;
	    RECT 35.7000 85.6000 37.8000 85.7000 ;
	    RECT 35.8000 85.4000 37.8000 85.6000 ;
	    RECT 35.0000 84.8000 35.7000 85.1000 ;
	    RECT 35.3000 81.1000 35.7000 84.8000 ;
	    RECT 37.4000 81.1000 37.8000 85.4000 ;
	    RECT 39.0000 81.1000 39.4000 87.9000 ;
	    RECT 42.4000 87.1000 42.8000 89.9000 ;
	    RECT 45.6000 87.1000 46.0000 89.9000 ;
	    RECT 42.4000 86.9000 43.3000 87.1000 ;
	    RECT 45.6000 86.9000 46.5000 87.1000 ;
	    RECT 42.5000 86.8000 43.3000 86.9000 ;
	    RECT 45.7000 86.8000 46.5000 86.9000 ;
	    RECT 41.4000 85.8000 42.2000 86.2000 ;
	    RECT 43.0000 85.2000 43.3000 86.8000 ;
	    RECT 44.6000 85.8000 45.4000 86.2000 ;
	    RECT 39.8000 84.4000 40.2000 85.2000 ;
	    RECT 43.0000 84.8000 43.4000 85.2000 ;
	    RECT 43.8000 84.8000 44.2000 85.6000 ;
	    RECT 46.2000 85.2000 46.5000 86.8000 ;
	    RECT 46.2000 84.8000 46.6000 85.2000 ;
	    RECT 47.8000 85.1000 48.2000 89.9000 ;
	    RECT 49.9000 88.2000 50.3000 89.9000 ;
	    RECT 51.8000 88.9000 52.2000 89.9000 ;
	    RECT 49.4000 87.9000 50.3000 88.2000 ;
	    RECT 48.6000 86.8000 49.0000 87.6000 ;
	    RECT 48.6000 85.8000 49.0000 86.2000 ;
	    RECT 48.6000 85.1000 48.9000 85.8000 ;
	    RECT 47.8000 84.8000 48.9000 85.1000 ;
	    RECT 42.2000 83.8000 42.6000 84.6000 ;
	    RECT 43.0000 84.1000 43.3000 84.8000 ;
	    RECT 45.4000 84.1000 45.8000 84.6000 ;
	    RECT 43.0000 83.8000 45.8000 84.1000 ;
	    RECT 43.0000 83.5000 43.3000 83.8000 ;
	    RECT 46.2000 83.5000 46.5000 84.8000 ;
	    RECT 41.5000 83.2000 43.3000 83.5000 ;
	    RECT 41.5000 83.1000 41.8000 83.2000 ;
	    RECT 41.4000 81.1000 41.8000 83.1000 ;
	    RECT 43.0000 83.1000 43.3000 83.2000 ;
	    RECT 44.7000 83.2000 46.5000 83.5000 ;
	    RECT 44.7000 83.1000 45.0000 83.2000 ;
	    RECT 43.0000 81.1000 43.4000 83.1000 ;
	    RECT 44.6000 81.1000 45.0000 83.1000 ;
	    RECT 46.2000 83.1000 46.5000 83.2000 ;
	    RECT 46.2000 81.1000 46.6000 83.1000 ;
	    RECT 47.8000 81.1000 48.2000 84.8000 ;
	    RECT 48.6000 84.1000 49.0000 84.2000 ;
	    RECT 49.4000 84.1000 49.8000 87.9000 ;
	    RECT 51.0000 87.8000 51.4000 88.6000 ;
	    RECT 51.9000 87.8000 52.2000 88.9000 ;
	    RECT 53.4000 87.9000 53.8000 89.9000 ;
	    RECT 51.9000 87.5000 53.1000 87.8000 ;
	    RECT 52.8000 86.0000 53.1000 87.5000 ;
	    RECT 53.5000 86.2000 53.8000 87.9000 ;
	    RECT 54.8000 87.1000 55.2000 89.9000 ;
	    RECT 58.2000 88.9000 58.6000 89.9000 ;
	    RECT 57.4000 87.8000 57.8000 88.6000 ;
	    RECT 58.3000 87.8000 58.6000 88.9000 ;
	    RECT 59.8000 87.9000 60.2000 89.9000 ;
	    RECT 58.3000 87.5000 59.5000 87.8000 ;
	    RECT 52.7000 85.7000 53.1000 86.0000 ;
	    RECT 53.4000 85.8000 53.8000 86.2000 ;
	    RECT 51.0000 85.6000 53.1000 85.7000 ;
	    RECT 51.0000 85.4000 53.0000 85.6000 ;
	    RECT 50.2000 84.4000 50.6000 85.2000 ;
	    RECT 48.6000 83.8000 49.8000 84.1000 ;
	    RECT 49.4000 81.1000 49.8000 83.8000 ;
	    RECT 51.0000 81.1000 51.4000 85.4000 ;
	    RECT 53.5000 85.1000 53.8000 85.8000 ;
	    RECT 54.3000 86.9000 55.2000 87.1000 ;
	    RECT 54.3000 86.8000 55.1000 86.9000 ;
	    RECT 54.3000 85.2000 54.6000 86.8000 ;
	    RECT 55.4000 85.8000 56.2000 86.2000 ;
	    RECT 59.2000 86.0000 59.5000 87.5000 ;
	    RECT 59.9000 86.2000 60.2000 87.9000 ;
	    RECT 59.1000 85.7000 59.5000 86.0000 ;
	    RECT 59.8000 86.1000 60.2000 86.2000 ;
	    RECT 61.4000 86.1000 61.8000 86.2000 ;
	    RECT 59.8000 85.8000 61.8000 86.1000 ;
	    RECT 57.4000 85.6000 59.5000 85.7000 ;
	    RECT 53.1000 84.8000 53.8000 85.1000 ;
	    RECT 54.2000 84.8000 54.6000 85.2000 ;
	    RECT 56.6000 84.8000 57.0000 85.6000 ;
	    RECT 57.4000 85.4000 59.4000 85.6000 ;
	    RECT 53.1000 81.1000 53.5000 84.8000 ;
	    RECT 54.3000 83.5000 54.6000 84.8000 ;
	    RECT 55.0000 83.8000 55.4000 84.6000 ;
	    RECT 54.3000 83.2000 56.1000 83.5000 ;
	    RECT 54.3000 83.1000 54.6000 83.2000 ;
	    RECT 54.2000 81.1000 54.6000 83.1000 ;
	    RECT 55.8000 83.1000 56.1000 83.2000 ;
	    RECT 55.8000 81.1000 56.2000 83.1000 ;
	    RECT 57.4000 81.1000 57.8000 85.4000 ;
	    RECT 59.9000 85.1000 60.2000 85.8000 ;
	    RECT 59.5000 84.8000 60.2000 85.1000 ;
	    RECT 59.5000 81.1000 59.9000 84.8000 ;
	    RECT 62.2000 84.1000 62.6000 84.2000 ;
	    RECT 63.0000 84.1000 63.4000 89.9000 ;
	    RECT 63.8000 87.6000 64.2000 89.9000 ;
	    RECT 63.8000 87.3000 64.9000 87.6000 ;
	    RECT 64.6000 85.8000 64.9000 87.3000 ;
	    RECT 65.4000 87.1000 65.8000 89.9000 ;
	    RECT 67.5000 88.2000 67.9000 89.9000 ;
	    RECT 68.9000 89.2000 69.3000 89.9000 ;
	    RECT 68.6000 88.8000 69.3000 89.2000 ;
	    RECT 67.0000 87.9000 67.9000 88.2000 ;
	    RECT 68.9000 88.2000 69.3000 88.8000 ;
	    RECT 68.9000 87.9000 69.8000 88.2000 ;
	    RECT 66.2000 87.1000 66.6000 87.6000 ;
	    RECT 65.4000 86.8000 66.6000 87.1000 ;
	    RECT 65.4000 86.2000 65.8000 86.8000 ;
	    RECT 64.6000 85.4000 65.2000 85.8000 ;
	    RECT 64.6000 85.1000 64.9000 85.4000 ;
	    RECT 65.5000 85.1000 65.8000 86.2000 ;
	    RECT 62.2000 83.8000 63.4000 84.1000 ;
	    RECT 63.0000 81.1000 63.4000 83.8000 ;
	    RECT 63.8000 84.8000 64.9000 85.1000 ;
	    RECT 63.8000 81.1000 64.2000 84.8000 ;
	    RECT 65.4000 81.1000 65.8000 85.1000 ;
	    RECT 67.0000 81.1000 67.4000 87.9000 ;
	    RECT 67.8000 84.4000 68.2000 85.2000 ;
	    RECT 68.6000 84.4000 69.0000 85.2000 ;
	    RECT 69.4000 81.1000 69.8000 87.9000 ;
	    RECT 71.6000 87.2000 72.0000 89.9000 ;
	    RECT 72.6000 87.8000 73.0000 88.2000 ;
	    RECT 71.6000 87.1000 72.2000 87.2000 ;
	    RECT 72.6000 87.1000 72.9000 87.8000 ;
	    RECT 74.8000 87.2000 75.2000 89.9000 ;
	    RECT 74.8000 87.1000 75.4000 87.2000 ;
	    RECT 78.0000 87.1000 78.4000 89.9000 ;
	    RECT 71.1000 86.8000 72.9000 87.1000 ;
	    RECT 74.3000 86.8000 75.4000 87.1000 ;
	    RECT 77.5000 86.9000 78.4000 87.1000 ;
	    RECT 82.4000 87.2000 82.8000 89.9000 ;
	    RECT 84.6000 88.9000 85.0000 89.9000 ;
	    RECT 83.8000 87.8000 84.2000 88.6000 ;
	    RECT 84.7000 87.8000 85.0000 88.9000 ;
	    RECT 86.2000 87.9000 86.6000 89.9000 ;
	    RECT 88.3000 89.2000 88.7000 89.9000 ;
	    RECT 89.7000 89.2000 90.1000 89.9000 ;
	    RECT 88.3000 88.8000 89.0000 89.2000 ;
	    RECT 89.7000 88.8000 90.6000 89.2000 ;
	    RECT 88.3000 88.2000 88.7000 88.8000 ;
	    RECT 84.7000 87.5000 85.9000 87.8000 ;
	    RECT 82.4000 86.9000 83.4000 87.2000 ;
	    RECT 77.5000 86.8000 78.3000 86.9000 ;
	    RECT 82.5000 86.8000 83.4000 86.9000 ;
	    RECT 71.1000 85.2000 71.4000 86.8000 ;
	    RECT 72.2000 85.8000 73.0000 86.2000 ;
	    RECT 71.0000 84.8000 71.4000 85.2000 ;
	    RECT 73.4000 84.8000 73.8000 85.6000 ;
	    RECT 74.3000 85.2000 74.6000 86.8000 ;
	    RECT 75.4000 85.8000 76.2000 86.2000 ;
	    RECT 74.2000 84.8000 74.6000 85.2000 ;
	    RECT 76.6000 84.8000 77.0000 85.6000 ;
	    RECT 77.5000 85.2000 77.8000 86.8000 ;
	    RECT 78.6000 85.8000 79.4000 86.2000 ;
	    RECT 81.4000 85.8000 82.2000 86.2000 ;
	    RECT 77.4000 84.8000 77.8000 85.2000 ;
	    RECT 79.8000 85.1000 80.2000 85.6000 ;
	    RECT 80.6000 85.1000 81.0000 85.6000 ;
	    RECT 79.8000 84.8000 81.0000 85.1000 ;
	    RECT 83.0000 85.2000 83.3000 86.8000 ;
	    RECT 85.6000 86.0000 85.9000 87.5000 ;
	    RECT 86.3000 86.2000 86.6000 87.9000 ;
	    RECT 87.8000 87.9000 88.7000 88.2000 ;
	    RECT 89.7000 88.2000 90.1000 88.8000 ;
	    RECT 89.7000 87.9000 90.6000 88.2000 ;
	    RECT 87.0000 86.8000 87.4000 87.6000 ;
	    RECT 85.5000 85.7000 85.9000 86.0000 ;
	    RECT 86.2000 85.8000 86.6000 86.2000 ;
	    RECT 83.8000 85.6000 85.9000 85.7000 ;
	    RECT 83.8000 85.4000 85.8000 85.6000 ;
	    RECT 83.0000 84.8000 83.4000 85.2000 ;
	    RECT 71.1000 83.5000 71.4000 84.8000 ;
	    RECT 71.8000 83.8000 72.2000 84.6000 ;
	    RECT 74.3000 83.5000 74.6000 84.8000 ;
	    RECT 75.0000 83.8000 75.4000 84.6000 ;
	    RECT 77.5000 83.5000 77.8000 84.8000 ;
	    RECT 78.2000 83.8000 78.6000 84.6000 ;
	    RECT 81.4000 84.1000 81.8000 84.2000 ;
	    RECT 82.2000 84.1000 82.6000 84.6000 ;
	    RECT 81.4000 83.8000 82.6000 84.1000 ;
	    RECT 83.0000 83.5000 83.3000 84.8000 ;
	    RECT 71.1000 83.2000 72.9000 83.5000 ;
	    RECT 71.1000 83.1000 71.4000 83.2000 ;
	    RECT 71.0000 81.1000 71.4000 83.1000 ;
	    RECT 72.6000 83.1000 72.9000 83.2000 ;
	    RECT 74.3000 83.2000 76.1000 83.5000 ;
	    RECT 74.3000 83.1000 74.6000 83.2000 ;
	    RECT 72.6000 81.1000 73.0000 83.1000 ;
	    RECT 74.2000 81.1000 74.6000 83.1000 ;
	    RECT 75.8000 83.1000 76.1000 83.2000 ;
	    RECT 77.5000 83.2000 79.3000 83.5000 ;
	    RECT 77.5000 83.1000 77.8000 83.2000 ;
	    RECT 75.8000 81.1000 76.2000 83.1000 ;
	    RECT 77.4000 81.1000 77.8000 83.1000 ;
	    RECT 79.0000 83.1000 79.3000 83.2000 ;
	    RECT 81.5000 83.2000 83.3000 83.5000 ;
	    RECT 81.5000 83.1000 81.8000 83.2000 ;
	    RECT 79.0000 81.1000 79.4000 83.1000 ;
	    RECT 81.4000 81.1000 81.8000 83.1000 ;
	    RECT 83.0000 83.1000 83.3000 83.2000 ;
	    RECT 83.0000 81.1000 83.4000 83.1000 ;
	    RECT 83.8000 81.1000 84.2000 85.4000 ;
	    RECT 86.3000 85.1000 86.6000 85.8000 ;
	    RECT 85.9000 84.8000 86.6000 85.1000 ;
	    RECT 85.9000 81.1000 86.3000 84.8000 ;
	    RECT 87.8000 81.1000 88.2000 87.9000 ;
	    RECT 88.6000 84.4000 89.0000 85.2000 ;
	    RECT 89.4000 84.4000 89.8000 85.2000 ;
	    RECT 90.2000 81.1000 90.6000 87.9000 ;
	    RECT 91.0000 86.8000 91.4000 87.6000 ;
	    RECT 92.4000 87.1000 92.8000 89.9000 ;
	    RECT 95.6000 87.1000 96.0000 89.9000 ;
	    RECT 98.8000 87.1000 99.2000 89.9000 ;
	    RECT 101.4000 87.5000 101.8000 89.9000 ;
	    RECT 103.6000 89.2000 104.0000 89.9000 ;
	    RECT 103.0000 88.9000 104.0000 89.2000 ;
	    RECT 105.8000 88.9000 106.2000 89.9000 ;
	    RECT 107.9000 89.2000 108.5000 89.9000 ;
	    RECT 107.8000 88.9000 108.5000 89.2000 ;
	    RECT 103.0000 88.5000 103.4000 88.9000 ;
	    RECT 105.8000 88.6000 106.1000 88.9000 ;
	    RECT 103.8000 88.2000 104.2000 88.6000 ;
	    RECT 104.7000 88.3000 106.1000 88.6000 ;
	    RECT 107.8000 88.5000 108.2000 88.9000 ;
	    RECT 104.7000 88.2000 105.1000 88.3000 ;
	    RECT 103.9000 87.2000 104.2000 88.2000 ;
	    RECT 108.7000 87.7000 109.1000 87.8000 ;
	    RECT 110.2000 87.7000 110.6000 89.9000 ;
	    RECT 108.7000 87.4000 110.6000 87.7000 ;
	    RECT 91.9000 86.9000 92.8000 87.1000 ;
	    RECT 95.1000 86.9000 96.0000 87.1000 ;
	    RECT 98.3000 86.9000 99.2000 87.1000 ;
	    RECT 101.8000 87.1000 102.6000 87.2000 ;
	    RECT 103.8000 87.1000 104.2000 87.2000 ;
	    RECT 106.7000 87.1000 107.1000 87.2000 ;
	    RECT 91.9000 86.8000 92.7000 86.9000 ;
	    RECT 95.1000 86.8000 95.9000 86.9000 ;
	    RECT 98.3000 86.8000 99.1000 86.9000 ;
	    RECT 101.8000 86.8000 107.3000 87.1000 ;
	    RECT 91.9000 85.2000 92.2000 86.8000 ;
	    RECT 93.0000 85.8000 93.8000 86.2000 ;
	    RECT 91.8000 84.8000 92.2000 85.2000 ;
	    RECT 94.2000 84.8000 94.6000 85.6000 ;
	    RECT 95.1000 85.2000 95.4000 86.8000 ;
	    RECT 96.2000 85.8000 97.0000 86.2000 ;
	    RECT 95.0000 84.8000 95.4000 85.2000 ;
	    RECT 97.4000 84.8000 97.8000 85.6000 ;
	    RECT 98.3000 85.2000 98.6000 86.8000 ;
	    RECT 103.3000 86.7000 103.7000 86.8000 ;
	    RECT 102.5000 86.2000 102.9000 86.3000 ;
	    RECT 99.4000 85.8000 100.2000 86.2000 ;
	    RECT 102.5000 85.9000 105.0000 86.2000 ;
	    RECT 104.6000 85.8000 105.0000 85.9000 ;
	    RECT 98.2000 84.8000 98.6000 85.2000 ;
	    RECT 100.6000 84.8000 101.0000 85.6000 ;
	    RECT 101.4000 85.5000 104.2000 85.6000 ;
	    RECT 101.4000 85.4000 104.3000 85.5000 ;
	    RECT 101.4000 85.3000 106.3000 85.4000 ;
	    RECT 91.9000 83.5000 92.2000 84.8000 ;
	    RECT 92.6000 83.8000 93.0000 84.6000 ;
	    RECT 95.1000 83.5000 95.4000 84.8000 ;
	    RECT 95.8000 83.8000 96.2000 84.6000 ;
	    RECT 98.3000 83.5000 98.6000 84.8000 ;
	    RECT 99.0000 83.8000 99.4000 84.6000 ;
	    RECT 91.9000 83.2000 93.7000 83.5000 ;
	    RECT 91.9000 83.1000 92.2000 83.2000 ;
	    RECT 91.8000 81.1000 92.2000 83.1000 ;
	    RECT 93.4000 83.1000 93.7000 83.2000 ;
	    RECT 95.1000 83.2000 96.9000 83.5000 ;
	    RECT 95.1000 83.1000 95.4000 83.2000 ;
	    RECT 93.4000 81.1000 93.8000 83.1000 ;
	    RECT 95.0000 81.1000 95.4000 83.1000 ;
	    RECT 96.6000 83.1000 96.9000 83.2000 ;
	    RECT 98.3000 83.2000 100.1000 83.5000 ;
	    RECT 98.3000 83.1000 98.6000 83.2000 ;
	    RECT 96.6000 81.1000 97.0000 83.1000 ;
	    RECT 98.2000 81.1000 98.6000 83.1000 ;
	    RECT 99.8000 83.1000 100.1000 83.2000 ;
	    RECT 99.8000 81.1000 100.2000 83.1000 ;
	    RECT 101.4000 81.1000 101.8000 85.3000 ;
	    RECT 103.9000 85.1000 106.3000 85.3000 ;
	    RECT 103.0000 84.5000 105.7000 84.8000 ;
	    RECT 103.0000 84.4000 103.4000 84.5000 ;
	    RECT 105.3000 84.4000 105.7000 84.5000 ;
	    RECT 106.0000 84.5000 106.3000 85.1000 ;
	    RECT 107.0000 85.2000 107.3000 86.8000 ;
	    RECT 107.8000 86.4000 108.2000 86.5000 ;
	    RECT 107.8000 86.1000 109.7000 86.4000 ;
	    RECT 109.3000 86.0000 109.7000 86.1000 ;
	    RECT 110.2000 86.1000 110.6000 87.4000 ;
	    RECT 111.0000 86.1000 111.4000 86.2000 ;
	    RECT 110.2000 85.8000 111.4000 86.1000 ;
	    RECT 108.5000 85.7000 108.9000 85.8000 ;
	    RECT 110.2000 85.7000 110.6000 85.8000 ;
	    RECT 108.5000 85.4000 110.6000 85.7000 ;
	    RECT 107.0000 84.9000 108.2000 85.2000 ;
	    RECT 106.7000 84.5000 107.1000 84.6000 ;
	    RECT 106.0000 84.2000 107.1000 84.5000 ;
	    RECT 107.9000 84.4000 108.2000 84.9000 ;
	    RECT 107.9000 84.0000 108.6000 84.4000 ;
	    RECT 104.7000 83.7000 105.1000 83.8000 ;
	    RECT 106.1000 83.7000 106.5000 83.8000 ;
	    RECT 103.0000 83.1000 103.4000 83.5000 ;
	    RECT 104.7000 83.4000 106.5000 83.7000 ;
	    RECT 105.8000 83.1000 106.1000 83.4000 ;
	    RECT 107.8000 83.1000 108.2000 83.5000 ;
	    RECT 103.0000 82.8000 104.0000 83.1000 ;
	    RECT 103.6000 81.1000 104.0000 82.8000 ;
	    RECT 105.8000 81.1000 106.2000 83.1000 ;
	    RECT 107.9000 81.1000 108.5000 83.1000 ;
	    RECT 110.2000 81.1000 110.6000 85.4000 ;
	    RECT 111.0000 82.1000 111.4000 82.2000 ;
	    RECT 112.6000 82.1000 113.0000 89.9000 ;
	    RECT 113.4000 87.1000 113.8000 87.6000 ;
	    RECT 114.2000 87.1000 114.6000 89.9000 ;
	    RECT 115.8000 87.6000 116.2000 89.9000 ;
	    RECT 116.9000 89.2000 117.3000 89.9000 ;
	    RECT 116.6000 88.8000 117.3000 89.2000 ;
	    RECT 116.9000 88.4000 117.3000 88.8000 ;
	    RECT 113.4000 86.8000 114.6000 87.1000 ;
	    RECT 111.0000 81.8000 113.0000 82.1000 ;
	    RECT 112.6000 81.1000 113.0000 81.8000 ;
	    RECT 114.2000 86.2000 114.6000 86.8000 ;
	    RECT 115.1000 87.3000 116.2000 87.6000 ;
	    RECT 116.6000 87.9000 117.3000 88.4000 ;
	    RECT 119.0000 87.9000 119.4000 89.9000 ;
	    RECT 114.2000 85.1000 114.5000 86.2000 ;
	    RECT 115.1000 85.8000 115.4000 87.3000 ;
	    RECT 114.8000 85.4000 115.4000 85.8000 ;
	    RECT 115.1000 85.1000 115.4000 85.4000 ;
	    RECT 116.6000 86.2000 116.9000 87.9000 ;
	    RECT 119.0000 87.8000 119.3000 87.9000 ;
	    RECT 118.4000 87.6000 119.3000 87.8000 ;
	    RECT 117.2000 87.5000 119.3000 87.6000 ;
	    RECT 119.8000 87.7000 120.2000 89.9000 ;
	    RECT 121.9000 89.2000 122.5000 89.9000 ;
	    RECT 121.9000 88.9000 122.6000 89.2000 ;
	    RECT 124.2000 88.9000 124.6000 89.9000 ;
	    RECT 126.4000 89.2000 126.8000 89.9000 ;
	    RECT 126.4000 88.9000 127.4000 89.2000 ;
	    RECT 122.2000 88.5000 122.6000 88.9000 ;
	    RECT 124.3000 88.6000 124.6000 88.9000 ;
	    RECT 124.3000 88.3000 125.7000 88.6000 ;
	    RECT 125.3000 88.2000 125.7000 88.3000 ;
	    RECT 126.2000 88.2000 126.6000 88.6000 ;
	    RECT 127.0000 88.5000 127.4000 88.9000 ;
	    RECT 121.3000 87.7000 121.7000 87.8000 ;
	    RECT 117.2000 87.3000 118.7000 87.5000 ;
	    RECT 119.8000 87.4000 121.7000 87.7000 ;
	    RECT 117.2000 87.2000 117.6000 87.3000 ;
	    RECT 116.6000 85.8000 117.0000 86.2000 ;
	    RECT 116.6000 85.1000 116.9000 85.8000 ;
	    RECT 117.3000 85.5000 117.6000 87.2000 ;
	    RECT 118.0000 86.6000 118.6000 87.0000 ;
	    RECT 118.2000 86.2000 118.5000 86.6000 ;
	    RECT 119.0000 86.4000 119.4000 87.2000 ;
	    RECT 118.2000 85.8000 118.6000 86.2000 ;
	    RECT 119.8000 85.7000 120.2000 87.4000 ;
	    RECT 123.3000 87.1000 123.7000 87.2000 ;
	    RECT 126.2000 87.1000 126.5000 88.2000 ;
	    RECT 128.6000 87.5000 129.0000 89.9000 ;
	    RECT 129.4000 87.9000 129.8000 89.9000 ;
	    RECT 131.5000 89.2000 131.9000 89.9000 ;
	    RECT 131.5000 88.8000 132.2000 89.2000 ;
	    RECT 131.5000 88.4000 131.9000 88.8000 ;
	    RECT 131.5000 87.9000 132.2000 88.4000 ;
	    RECT 129.5000 87.8000 129.8000 87.9000 ;
	    RECT 129.5000 87.6000 130.4000 87.8000 ;
	    RECT 129.5000 87.5000 131.6000 87.6000 ;
	    RECT 130.1000 87.3000 131.6000 87.5000 ;
	    RECT 131.2000 87.2000 131.6000 87.3000 ;
	    RECT 127.8000 87.1000 128.6000 87.2000 ;
	    RECT 123.1000 86.8000 128.6000 87.1000 ;
	    RECT 122.2000 86.4000 122.6000 86.5000 ;
	    RECT 120.7000 86.1000 122.6000 86.4000 ;
	    RECT 120.7000 86.0000 121.1000 86.1000 ;
	    RECT 121.5000 85.7000 121.9000 85.8000 ;
	    RECT 117.3000 85.2000 118.5000 85.5000 ;
	    RECT 114.2000 81.1000 114.6000 85.1000 ;
	    RECT 115.1000 84.8000 116.2000 85.1000 ;
	    RECT 115.8000 81.1000 116.2000 84.8000 ;
	    RECT 116.6000 81.1000 117.0000 85.1000 ;
	    RECT 118.2000 83.1000 118.5000 85.2000 ;
	    RECT 119.8000 85.4000 121.9000 85.7000 ;
	    RECT 118.2000 81.1000 118.6000 83.1000 ;
	    RECT 119.8000 81.1000 120.2000 85.4000 ;
	    RECT 123.1000 85.2000 123.4000 86.8000 ;
	    RECT 126.7000 86.7000 127.1000 86.8000 ;
	    RECT 129.4000 86.4000 129.8000 87.2000 ;
	    RECT 130.4000 86.9000 130.8000 87.0000 ;
	    RECT 130.3000 86.6000 130.8000 86.9000 ;
	    RECT 127.5000 86.2000 127.9000 86.3000 ;
	    RECT 130.3000 86.2000 130.6000 86.6000 ;
	    RECT 125.4000 85.9000 127.9000 86.2000 ;
	    RECT 125.4000 85.8000 125.8000 85.9000 ;
	    RECT 130.2000 85.8000 130.6000 86.2000 ;
	    RECT 126.2000 85.5000 129.0000 85.6000 ;
	    RECT 131.2000 85.5000 131.5000 87.2000 ;
	    RECT 131.9000 86.2000 132.2000 87.9000 ;
	    RECT 132.6000 87.5000 133.0000 89.9000 ;
	    RECT 134.8000 89.2000 135.2000 89.9000 ;
	    RECT 134.2000 88.9000 135.2000 89.2000 ;
	    RECT 137.0000 88.9000 137.4000 89.9000 ;
	    RECT 139.1000 89.2000 139.7000 89.9000 ;
	    RECT 139.0000 88.9000 139.7000 89.2000 ;
	    RECT 134.2000 88.5000 134.6000 88.9000 ;
	    RECT 137.0000 88.6000 137.3000 88.9000 ;
	    RECT 135.0000 88.2000 135.4000 88.6000 ;
	    RECT 135.9000 88.3000 137.3000 88.6000 ;
	    RECT 139.0000 88.5000 139.4000 88.9000 ;
	    RECT 135.9000 88.2000 136.3000 88.3000 ;
	    RECT 133.0000 87.1000 133.8000 87.2000 ;
	    RECT 135.1000 87.1000 135.4000 88.2000 ;
	    RECT 139.9000 87.7000 140.3000 87.8000 ;
	    RECT 141.4000 87.7000 141.8000 89.9000 ;
	    RECT 142.3000 88.2000 142.7000 88.6000 ;
	    RECT 142.2000 87.8000 142.6000 88.2000 ;
	    RECT 143.0000 87.9000 143.4000 89.9000 ;
	    RECT 139.9000 87.4000 141.8000 87.7000 ;
	    RECT 137.9000 87.1000 138.3000 87.2000 ;
	    RECT 133.0000 86.8000 138.5000 87.1000 ;
	    RECT 134.5000 86.7000 134.9000 86.8000 ;
	    RECT 131.8000 85.8000 132.2000 86.2000 ;
	    RECT 133.7000 86.2000 134.1000 86.3000 ;
	    RECT 135.0000 86.2000 135.4000 86.3000 ;
	    RECT 133.7000 85.9000 136.2000 86.2000 ;
	    RECT 135.8000 85.8000 136.2000 85.9000 ;
	    RECT 126.1000 85.4000 129.0000 85.5000 ;
	    RECT 122.2000 84.9000 123.4000 85.2000 ;
	    RECT 124.1000 85.3000 129.0000 85.4000 ;
	    RECT 124.1000 85.1000 126.5000 85.3000 ;
	    RECT 122.2000 84.4000 122.5000 84.9000 ;
	    RECT 121.8000 84.0000 122.5000 84.4000 ;
	    RECT 123.3000 84.5000 123.7000 84.6000 ;
	    RECT 124.1000 84.5000 124.4000 85.1000 ;
	    RECT 123.3000 84.2000 124.4000 84.5000 ;
	    RECT 124.7000 84.5000 127.4000 84.8000 ;
	    RECT 124.7000 84.4000 125.1000 84.5000 ;
	    RECT 127.0000 84.4000 127.4000 84.5000 ;
	    RECT 123.9000 83.7000 124.3000 83.8000 ;
	    RECT 125.3000 83.7000 125.7000 83.8000 ;
	    RECT 122.2000 83.1000 122.6000 83.5000 ;
	    RECT 123.9000 83.4000 125.7000 83.7000 ;
	    RECT 124.3000 83.1000 124.6000 83.4000 ;
	    RECT 127.0000 83.1000 127.4000 83.5000 ;
	    RECT 121.9000 81.1000 122.5000 83.1000 ;
	    RECT 124.2000 81.1000 124.6000 83.1000 ;
	    RECT 126.4000 82.8000 127.4000 83.1000 ;
	    RECT 126.4000 81.1000 126.8000 82.8000 ;
	    RECT 128.6000 81.1000 129.0000 85.3000 ;
	    RECT 130.3000 85.2000 131.5000 85.5000 ;
	    RECT 130.3000 83.1000 130.6000 85.2000 ;
	    RECT 131.9000 85.1000 132.2000 85.8000 ;
	    RECT 130.2000 81.1000 130.6000 83.1000 ;
	    RECT 131.8000 81.1000 132.2000 85.1000 ;
	    RECT 132.6000 85.5000 135.4000 85.6000 ;
	    RECT 132.6000 85.4000 135.5000 85.5000 ;
	    RECT 132.6000 85.3000 137.5000 85.4000 ;
	    RECT 132.6000 81.1000 133.0000 85.3000 ;
	    RECT 135.1000 85.1000 137.5000 85.3000 ;
	    RECT 134.2000 84.5000 136.9000 84.8000 ;
	    RECT 134.2000 84.4000 134.6000 84.5000 ;
	    RECT 136.5000 84.4000 136.9000 84.5000 ;
	    RECT 137.2000 84.5000 137.5000 85.1000 ;
	    RECT 138.2000 85.2000 138.5000 86.8000 ;
	    RECT 139.0000 86.4000 139.4000 86.5000 ;
	    RECT 139.0000 86.1000 140.9000 86.4000 ;
	    RECT 140.5000 86.0000 140.9000 86.1000 ;
	    RECT 139.7000 85.7000 140.1000 85.8000 ;
	    RECT 141.4000 85.7000 141.8000 87.4000 ;
	    RECT 142.2000 86.1000 142.6000 86.2000 ;
	    RECT 143.1000 86.1000 143.4000 87.9000 ;
	    RECT 146.2000 87.6000 146.6000 89.9000 ;
	    RECT 147.8000 87.6000 148.2000 89.9000 ;
	    RECT 149.4000 87.6000 149.8000 89.9000 ;
	    RECT 151.0000 87.6000 151.4000 89.9000 ;
	    RECT 152.6000 87.7000 153.0000 89.9000 ;
	    RECT 154.7000 89.2000 155.3000 89.9000 ;
	    RECT 154.7000 88.9000 155.4000 89.2000 ;
	    RECT 157.0000 88.9000 157.4000 89.9000 ;
	    RECT 159.2000 89.2000 159.6000 89.9000 ;
	    RECT 159.2000 88.9000 160.2000 89.2000 ;
	    RECT 155.0000 88.5000 155.4000 88.9000 ;
	    RECT 157.1000 88.6000 157.4000 88.9000 ;
	    RECT 157.1000 88.3000 158.5000 88.6000 ;
	    RECT 158.1000 88.2000 158.5000 88.3000 ;
	    RECT 159.0000 88.2000 159.4000 88.6000 ;
	    RECT 159.8000 88.5000 160.2000 88.9000 ;
	    RECT 154.1000 87.7000 154.5000 87.8000 ;
	    RECT 146.2000 87.2000 147.1000 87.6000 ;
	    RECT 147.8000 87.2000 148.9000 87.6000 ;
	    RECT 149.4000 87.2000 150.5000 87.6000 ;
	    RECT 151.0000 87.2000 152.2000 87.6000 ;
	    RECT 143.8000 86.4000 144.2000 87.2000 ;
	    RECT 146.7000 86.9000 147.1000 87.2000 ;
	    RECT 148.5000 86.9000 148.9000 87.2000 ;
	    RECT 150.1000 86.9000 150.5000 87.2000 ;
	    RECT 146.7000 86.5000 148.0000 86.9000 ;
	    RECT 148.5000 86.5000 149.7000 86.9000 ;
	    RECT 150.1000 86.5000 151.4000 86.9000 ;
	    RECT 144.6000 86.1000 145.0000 86.2000 ;
	    RECT 142.2000 85.8000 143.4000 86.1000 ;
	    RECT 144.2000 85.8000 145.0000 86.1000 ;
	    RECT 146.7000 85.8000 147.1000 86.5000 ;
	    RECT 148.5000 85.8000 148.9000 86.5000 ;
	    RECT 150.1000 85.8000 150.5000 86.5000 ;
	    RECT 151.8000 85.8000 152.2000 87.2000 ;
	    RECT 139.7000 85.4000 141.8000 85.7000 ;
	    RECT 138.2000 84.9000 139.4000 85.2000 ;
	    RECT 137.9000 84.5000 138.3000 84.6000 ;
	    RECT 137.2000 84.2000 138.3000 84.5000 ;
	    RECT 139.1000 84.4000 139.4000 84.9000 ;
	    RECT 139.1000 84.0000 139.8000 84.4000 ;
	    RECT 135.9000 83.7000 136.3000 83.8000 ;
	    RECT 137.3000 83.7000 137.7000 83.8000 ;
	    RECT 134.2000 83.1000 134.6000 83.5000 ;
	    RECT 135.9000 83.4000 137.7000 83.7000 ;
	    RECT 137.0000 83.1000 137.3000 83.4000 ;
	    RECT 139.0000 83.1000 139.4000 83.5000 ;
	    RECT 134.2000 82.8000 135.2000 83.1000 ;
	    RECT 134.8000 81.1000 135.2000 82.8000 ;
	    RECT 137.0000 81.1000 137.4000 83.1000 ;
	    RECT 139.1000 81.1000 139.7000 83.1000 ;
	    RECT 141.4000 81.1000 141.8000 85.4000 ;
	    RECT 142.3000 85.1000 142.6000 85.8000 ;
	    RECT 144.2000 85.6000 144.6000 85.8000 ;
	    RECT 146.2000 85.4000 147.1000 85.8000 ;
	    RECT 147.8000 85.4000 148.9000 85.8000 ;
	    RECT 149.4000 85.4000 150.5000 85.8000 ;
	    RECT 151.0000 85.4000 152.2000 85.8000 ;
	    RECT 152.6000 87.4000 154.5000 87.7000 ;
	    RECT 152.6000 85.7000 153.0000 87.4000 ;
	    RECT 159.0000 87.2000 159.3000 88.2000 ;
	    RECT 161.4000 87.5000 161.8000 89.9000 ;
	    RECT 162.2000 87.9000 162.6000 89.9000 ;
	    RECT 164.3000 89.2000 164.7000 89.9000 ;
	    RECT 165.7000 89.2000 166.1000 89.9000 ;
	    RECT 164.3000 88.8000 165.0000 89.2000 ;
	    RECT 165.4000 88.8000 166.1000 89.2000 ;
	    RECT 164.3000 88.4000 164.7000 88.8000 ;
	    RECT 165.7000 88.4000 166.1000 88.8000 ;
	    RECT 164.3000 87.9000 165.0000 88.4000 ;
	    RECT 162.3000 87.8000 162.6000 87.9000 ;
	    RECT 162.3000 87.6000 163.2000 87.8000 ;
	    RECT 162.3000 87.5000 164.4000 87.6000 ;
	    RECT 162.9000 87.3000 164.4000 87.5000 ;
	    RECT 164.0000 87.2000 164.4000 87.3000 ;
	    RECT 156.1000 87.1000 156.5000 87.2000 ;
	    RECT 159.0000 87.1000 159.4000 87.2000 ;
	    RECT 160.6000 87.1000 161.4000 87.2000 ;
	    RECT 155.9000 86.8000 161.4000 87.1000 ;
	    RECT 155.0000 86.4000 155.4000 86.5000 ;
	    RECT 153.5000 86.1000 155.4000 86.4000 ;
	    RECT 153.5000 86.0000 153.9000 86.1000 ;
	    RECT 154.3000 85.7000 154.7000 85.8000 ;
	    RECT 152.6000 85.4000 154.7000 85.7000 ;
	    RECT 142.2000 81.1000 142.6000 85.1000 ;
	    RECT 143.0000 84.8000 145.0000 85.1000 ;
	    RECT 143.0000 81.1000 143.4000 84.8000 ;
	    RECT 144.6000 81.1000 145.0000 84.8000 ;
	    RECT 146.2000 81.1000 146.6000 85.4000 ;
	    RECT 147.8000 81.1000 148.2000 85.4000 ;
	    RECT 149.4000 81.1000 149.8000 85.4000 ;
	    RECT 151.0000 81.1000 151.4000 85.4000 ;
	    RECT 152.6000 81.1000 153.0000 85.4000 ;
	    RECT 155.9000 85.2000 156.2000 86.8000 ;
	    RECT 159.5000 86.7000 159.9000 86.8000 ;
	    RECT 162.2000 86.4000 162.6000 87.2000 ;
	    RECT 163.2000 86.9000 163.6000 87.0000 ;
	    RECT 163.1000 86.6000 163.6000 86.9000 ;
	    RECT 160.3000 86.2000 160.7000 86.3000 ;
	    RECT 163.1000 86.2000 163.4000 86.6000 ;
	    RECT 157.4000 86.1000 157.8000 86.2000 ;
	    RECT 158.2000 86.1000 160.7000 86.2000 ;
	    RECT 157.4000 85.9000 160.7000 86.1000 ;
	    RECT 157.4000 85.8000 158.6000 85.9000 ;
	    RECT 163.0000 85.8000 163.4000 86.2000 ;
	    RECT 159.0000 85.5000 161.8000 85.6000 ;
	    RECT 164.0000 85.5000 164.3000 87.2000 ;
	    RECT 164.7000 86.2000 165.0000 87.9000 ;
	    RECT 164.6000 85.8000 165.0000 86.2000 ;
	    RECT 158.9000 85.4000 161.8000 85.5000 ;
	    RECT 155.0000 84.9000 156.2000 85.2000 ;
	    RECT 156.9000 85.3000 161.8000 85.4000 ;
	    RECT 156.9000 85.1000 159.3000 85.3000 ;
	    RECT 155.0000 84.4000 155.3000 84.9000 ;
	    RECT 154.6000 84.0000 155.3000 84.4000 ;
	    RECT 156.1000 84.5000 156.5000 84.6000 ;
	    RECT 156.9000 84.5000 157.2000 85.1000 ;
	    RECT 156.1000 84.2000 157.2000 84.5000 ;
	    RECT 157.5000 84.5000 160.2000 84.8000 ;
	    RECT 157.5000 84.4000 157.9000 84.5000 ;
	    RECT 159.8000 84.4000 160.2000 84.5000 ;
	    RECT 156.7000 83.7000 157.1000 83.8000 ;
	    RECT 158.1000 83.7000 158.5000 83.8000 ;
	    RECT 155.0000 83.1000 155.4000 83.5000 ;
	    RECT 156.7000 83.4000 158.5000 83.7000 ;
	    RECT 157.1000 83.1000 157.4000 83.4000 ;
	    RECT 159.8000 83.1000 160.2000 83.5000 ;
	    RECT 154.7000 81.1000 155.3000 83.1000 ;
	    RECT 157.0000 81.1000 157.4000 83.1000 ;
	    RECT 159.2000 82.8000 160.2000 83.1000 ;
	    RECT 159.2000 81.1000 159.6000 82.8000 ;
	    RECT 161.4000 81.1000 161.8000 85.3000 ;
	    RECT 163.1000 85.2000 164.3000 85.5000 ;
	    RECT 163.1000 83.1000 163.4000 85.2000 ;
	    RECT 164.7000 85.1000 165.0000 85.8000 ;
	    RECT 163.0000 81.1000 163.4000 83.1000 ;
	    RECT 164.6000 81.1000 165.0000 85.1000 ;
	    RECT 165.4000 87.9000 166.1000 88.4000 ;
	    RECT 167.8000 87.9000 168.2000 89.9000 ;
	    RECT 165.4000 86.2000 165.7000 87.9000 ;
	    RECT 167.8000 87.8000 168.1000 87.9000 ;
	    RECT 167.2000 87.6000 168.1000 87.8000 ;
	    RECT 166.0000 87.5000 168.1000 87.6000 ;
	    RECT 168.6000 87.6000 169.0000 89.9000 ;
	    RECT 171.3000 89.2000 171.7000 89.9000 ;
	    RECT 171.3000 88.8000 172.2000 89.2000 ;
	    RECT 171.3000 88.2000 171.7000 88.8000 ;
	    RECT 171.3000 87.9000 172.2000 88.2000 ;
	    RECT 166.0000 87.3000 167.5000 87.5000 ;
	    RECT 168.6000 87.3000 169.7000 87.6000 ;
	    RECT 166.0000 87.2000 166.4000 87.3000 ;
	    RECT 165.4000 85.8000 165.8000 86.2000 ;
	    RECT 165.4000 85.1000 165.7000 85.8000 ;
	    RECT 166.1000 85.5000 166.4000 87.2000 ;
	    RECT 166.8000 86.9000 167.2000 87.0000 ;
	    RECT 166.8000 86.6000 167.3000 86.9000 ;
	    RECT 167.0000 86.2000 167.3000 86.6000 ;
	    RECT 167.8000 86.4000 168.2000 87.2000 ;
	    RECT 167.0000 85.8000 167.4000 86.2000 ;
	    RECT 168.6000 85.8000 169.0000 86.6000 ;
	    RECT 169.4000 85.8000 169.7000 87.3000 ;
	    RECT 166.1000 85.2000 167.3000 85.5000 ;
	    RECT 165.4000 81.1000 165.8000 85.1000 ;
	    RECT 167.0000 83.1000 167.3000 85.2000 ;
	    RECT 169.4000 85.4000 170.0000 85.8000 ;
	    RECT 169.4000 85.1000 169.7000 85.4000 ;
	    RECT 168.6000 84.8000 169.7000 85.1000 ;
	    RECT 167.0000 81.1000 167.4000 83.1000 ;
	    RECT 168.6000 81.1000 169.0000 84.8000 ;
	    RECT 171.0000 84.4000 171.4000 85.2000 ;
	    RECT 171.8000 81.1000 172.2000 87.9000 ;
	    RECT 172.6000 86.8000 173.0000 87.6000 ;
	    RECT 0.6000 75.8000 1.0000 76.6000 ;
	    RECT 1.4000 73.1000 1.8000 79.9000 ;
	    RECT 3.3000 76.2000 3.7000 79.9000 ;
	    RECT 3.0000 75.9000 3.7000 76.2000 ;
	    RECT 3.0000 75.2000 3.3000 75.9000 ;
	    RECT 5.4000 75.6000 5.8000 79.9000 ;
	    RECT 6.2000 76.2000 6.6000 79.9000 ;
	    RECT 6.2000 75.9000 7.3000 76.2000 ;
	    RECT 7.8000 75.9000 8.2000 79.9000 ;
	    RECT 8.6000 76.2000 9.0000 79.9000 ;
	    RECT 8.6000 75.9000 9.7000 76.2000 ;
	    RECT 10.2000 75.9000 10.6000 79.9000 ;
	    RECT 3.8000 75.4000 5.8000 75.6000 ;
	    RECT 3.7000 75.3000 5.8000 75.4000 ;
	    RECT 7.0000 75.6000 7.3000 75.9000 ;
	    RECT 3.0000 74.8000 3.4000 75.2000 ;
	    RECT 3.7000 75.0000 4.1000 75.3000 ;
	    RECT 7.0000 75.2000 7.6000 75.6000 ;
	    RECT 2.2000 73.4000 2.6000 74.2000 ;
	    RECT 0.9000 72.8000 1.8000 73.1000 ;
	    RECT 3.0000 73.1000 3.3000 74.8000 ;
	    RECT 3.7000 73.5000 4.0000 75.0000 ;
	    RECT 7.0000 73.7000 7.3000 75.2000 ;
	    RECT 7.9000 74.8000 8.2000 75.9000 ;
	    RECT 3.7000 73.2000 4.9000 73.5000 ;
	    RECT 6.2000 73.4000 7.3000 73.7000 ;
	    RECT 0.9000 72.2000 1.3000 72.8000 ;
	    RECT 0.9000 71.8000 1.8000 72.2000 ;
	    RECT 0.9000 71.1000 1.3000 71.8000 ;
	    RECT 3.0000 71.1000 3.4000 73.1000 ;
	    RECT 4.6000 72.1000 4.9000 73.2000 ;
	    RECT 5.4000 72.4000 5.8000 73.2000 ;
	    RECT 4.6000 71.1000 5.0000 72.1000 ;
	    RECT 6.2000 71.1000 6.6000 73.4000 ;
	    RECT 7.8000 71.1000 8.2000 74.8000 ;
	    RECT 9.4000 75.6000 9.7000 75.9000 ;
	    RECT 9.4000 75.2000 10.0000 75.6000 ;
	    RECT 9.4000 73.7000 9.7000 75.2000 ;
	    RECT 10.3000 74.8000 10.6000 75.9000 ;
	    RECT 8.6000 73.4000 9.7000 73.7000 ;
	    RECT 8.6000 71.1000 9.0000 73.4000 ;
	    RECT 10.2000 71.1000 10.6000 74.8000 ;
	    RECT 11.0000 76.1000 11.4000 79.9000 ;
	    RECT 12.6000 76.1000 13.0000 76.6000 ;
	    RECT 11.0000 75.8000 13.0000 76.1000 ;
	    RECT 11.0000 71.1000 11.4000 75.8000 ;
	    RECT 13.4000 73.1000 13.8000 79.9000 ;
	    RECT 15.0000 75.6000 15.4000 79.9000 ;
	    RECT 17.1000 76.2000 17.5000 79.9000 ;
	    RECT 17.1000 75.9000 17.8000 76.2000 ;
	    RECT 15.0000 75.4000 17.0000 75.6000 ;
	    RECT 15.0000 75.3000 17.1000 75.4000 ;
	    RECT 16.7000 75.0000 17.1000 75.3000 ;
	    RECT 17.5000 75.2000 17.8000 75.9000 ;
	    RECT 14.2000 74.1000 14.6000 74.2000 ;
	    RECT 14.2000 73.8000 15.3000 74.1000 ;
	    RECT 14.2000 73.4000 14.6000 73.8000 ;
	    RECT 12.9000 72.8000 13.8000 73.1000 ;
	    RECT 15.0000 73.2000 15.3000 73.8000 ;
	    RECT 16.8000 73.5000 17.1000 75.0000 ;
	    RECT 17.4000 74.8000 17.8000 75.2000 ;
	    RECT 15.9000 73.2000 17.1000 73.5000 ;
	    RECT 12.9000 72.2000 13.3000 72.8000 ;
	    RECT 15.0000 72.4000 15.4000 73.2000 ;
	    RECT 12.6000 71.8000 13.3000 72.2000 ;
	    RECT 15.9000 72.1000 16.2000 73.2000 ;
	    RECT 17.5000 73.1000 17.8000 74.8000 ;
	    RECT 18.2000 73.4000 18.6000 74.2000 ;
	    RECT 12.9000 71.1000 13.3000 71.8000 ;
	    RECT 15.8000 71.1000 16.2000 72.1000 ;
	    RECT 17.4000 71.1000 17.8000 73.1000 ;
	    RECT 19.0000 73.1000 19.4000 79.9000 ;
	    RECT 19.8000 76.1000 20.2000 76.6000 ;
	    RECT 20.6000 76.1000 21.0000 79.9000 ;
	    RECT 19.8000 75.8000 21.0000 76.1000 ;
	    RECT 19.0000 72.8000 19.9000 73.1000 ;
	    RECT 19.5000 72.2000 19.9000 72.8000 ;
	    RECT 19.0000 71.8000 19.9000 72.2000 ;
	    RECT 19.5000 71.1000 19.9000 71.8000 ;
	    RECT 20.6000 71.1000 21.0000 75.8000 ;
	    RECT 22.2000 73.4000 22.6000 74.2000 ;
	    RECT 23.0000 73.1000 23.4000 79.9000 ;
	    RECT 23.8000 76.1000 24.2000 76.6000 ;
	    RECT 24.6000 76.1000 25.0000 79.9000 ;
	    RECT 23.8000 75.8000 25.0000 76.1000 ;
	    RECT 23.0000 72.8000 23.9000 73.1000 ;
	    RECT 23.5000 72.2000 23.9000 72.8000 ;
	    RECT 23.5000 71.8000 24.2000 72.2000 ;
	    RECT 23.5000 71.1000 23.9000 71.8000 ;
	    RECT 24.6000 71.1000 25.0000 75.8000 ;
	    RECT 27.0000 76.1000 27.4000 79.9000 ;
	    RECT 27.8000 76.1000 28.2000 76.6000 ;
	    RECT 27.0000 75.8000 28.2000 76.1000 ;
	    RECT 27.0000 71.1000 27.4000 75.8000 ;
	    RECT 27.8000 75.1000 28.2000 75.2000 ;
	    RECT 28.6000 75.1000 29.0000 79.9000 ;
	    RECT 30.5000 76.2000 30.9000 79.9000 ;
	    RECT 27.8000 74.8000 29.0000 75.1000 ;
	    RECT 28.6000 73.1000 29.0000 74.8000 ;
	    RECT 30.2000 75.9000 30.9000 76.2000 ;
	    RECT 30.2000 75.2000 30.5000 75.9000 ;
	    RECT 32.6000 75.6000 33.0000 79.9000 ;
	    RECT 31.0000 75.4000 33.0000 75.6000 ;
	    RECT 30.9000 75.3000 33.0000 75.4000 ;
	    RECT 30.2000 74.8000 30.6000 75.2000 ;
	    RECT 30.9000 75.0000 31.3000 75.3000 ;
	    RECT 29.4000 73.4000 29.8000 74.2000 ;
	    RECT 28.1000 72.8000 29.0000 73.1000 ;
	    RECT 30.2000 73.1000 30.5000 74.8000 ;
	    RECT 30.9000 73.5000 31.2000 75.0000 ;
	    RECT 31.6000 74.2000 32.0000 74.6000 ;
	    RECT 31.7000 73.8000 32.2000 74.2000 ;
	    RECT 30.9000 73.2000 32.1000 73.5000 ;
	    RECT 28.1000 71.1000 28.5000 72.8000 ;
	    RECT 30.2000 71.1000 30.6000 73.1000 ;
	    RECT 31.8000 72.1000 32.1000 73.2000 ;
	    RECT 31.8000 71.1000 32.2000 72.1000 ;
	    RECT 33.4000 71.1000 33.8000 79.9000 ;
	    RECT 35.0000 74.1000 35.4000 79.9000 ;
	    RECT 37.9000 79.2000 38.3000 79.9000 ;
	    RECT 37.4000 78.8000 38.3000 79.2000 ;
	    RECT 37.9000 76.2000 38.3000 78.8000 ;
	    RECT 38.6000 76.8000 39.0000 77.2000 ;
	    RECT 38.7000 76.2000 39.0000 76.8000 ;
	    RECT 37.9000 75.9000 38.4000 76.2000 ;
	    RECT 38.7000 75.9000 39.4000 76.2000 ;
	    RECT 35.8000 75.1000 36.2000 75.2000 ;
	    RECT 37.4000 75.1000 37.8000 75.2000 ;
	    RECT 35.8000 74.8000 37.8000 75.1000 ;
	    RECT 37.4000 74.4000 37.8000 74.8000 ;
	    RECT 38.1000 74.2000 38.4000 75.9000 ;
	    RECT 39.0000 75.8000 39.4000 75.9000 ;
	    RECT 36.6000 74.1000 37.0000 74.2000 ;
	    RECT 35.0000 73.8000 37.4000 74.1000 ;
	    RECT 38.1000 73.8000 39.4000 74.2000 ;
	    RECT 35.0000 71.1000 35.4000 73.8000 ;
	    RECT 37.0000 73.6000 37.4000 73.8000 ;
	    RECT 36.7000 73.1000 38.5000 73.3000 ;
	    RECT 39.0000 73.1000 39.3000 73.8000 ;
	    RECT 36.6000 73.0000 38.6000 73.1000 ;
	    RECT 36.6000 71.1000 37.0000 73.0000 ;
	    RECT 38.2000 71.1000 38.6000 73.0000 ;
	    RECT 39.0000 71.1000 39.4000 73.1000 ;
	    RECT 39.8000 71.1000 40.2000 79.9000 ;
	    RECT 42.2000 76.1000 42.6000 79.9000 ;
	    RECT 43.8000 77.1000 44.2000 79.9000 ;
	    RECT 43.8000 76.8000 44.9000 77.1000 ;
	    RECT 43.0000 76.1000 43.4000 76.6000 ;
	    RECT 42.2000 75.8000 43.4000 76.1000 ;
	    RECT 42.2000 71.1000 42.6000 75.8000 ;
	    RECT 43.8000 73.1000 44.2000 76.8000 ;
	    RECT 44.6000 76.2000 44.9000 76.8000 ;
	    RECT 44.6000 75.8000 45.0000 76.2000 ;
	    RECT 45.4000 75.6000 45.8000 79.9000 ;
	    RECT 47.5000 76.2000 47.9000 79.9000 ;
	    RECT 48.6000 77.9000 49.0000 79.9000 ;
	    RECT 48.7000 77.8000 49.0000 77.9000 ;
	    RECT 50.2000 77.9000 50.6000 79.9000 ;
	    RECT 50.2000 77.8000 50.5000 77.9000 ;
	    RECT 48.7000 77.5000 50.5000 77.8000 ;
	    RECT 48.7000 76.2000 49.0000 77.5000 ;
	    RECT 49.4000 76.4000 49.8000 77.2000 ;
	    RECT 47.5000 75.9000 48.2000 76.2000 ;
	    RECT 45.4000 75.4000 47.4000 75.6000 ;
	    RECT 45.4000 75.3000 47.5000 75.4000 ;
	    RECT 47.1000 75.0000 47.5000 75.3000 ;
	    RECT 47.9000 75.2000 48.2000 75.9000 ;
	    RECT 48.6000 75.8000 49.0000 76.2000 ;
	    RECT 46.4000 74.2000 46.8000 74.6000 ;
	    RECT 44.6000 74.1000 45.0000 74.2000 ;
	    RECT 46.2000 74.1000 46.7000 74.2000 ;
	    RECT 44.6000 73.8000 46.7000 74.1000 ;
	    RECT 44.6000 73.4000 45.0000 73.8000 ;
	    RECT 47.2000 73.5000 47.5000 75.0000 ;
	    RECT 47.8000 74.8000 48.2000 75.2000 ;
	    RECT 43.3000 72.8000 44.2000 73.1000 ;
	    RECT 46.3000 73.2000 47.5000 73.5000 ;
	    RECT 43.3000 71.1000 43.7000 72.8000 ;
	    RECT 46.3000 72.1000 46.6000 73.2000 ;
	    RECT 47.9000 73.1000 48.2000 74.8000 ;
	    RECT 48.7000 74.2000 49.0000 75.8000 ;
	    RECT 51.0000 75.4000 51.4000 76.2000 ;
	    RECT 51.8000 75.6000 52.2000 79.9000 ;
	    RECT 53.9000 76.2000 54.3000 79.9000 ;
	    RECT 53.9000 75.9000 54.6000 76.2000 ;
	    RECT 54.2000 75.8000 54.6000 75.9000 ;
	    RECT 51.8000 75.4000 53.8000 75.6000 ;
	    RECT 51.8000 75.3000 53.9000 75.4000 ;
	    RECT 49.8000 74.8000 50.6000 75.2000 ;
	    RECT 53.5000 75.0000 53.9000 75.3000 ;
	    RECT 54.3000 75.2000 54.6000 75.8000 ;
	    RECT 48.7000 74.1000 49.5000 74.2000 ;
	    RECT 48.7000 73.9000 49.6000 74.1000 ;
	    RECT 46.2000 71.1000 46.6000 72.1000 ;
	    RECT 47.8000 71.1000 48.2000 73.1000 ;
	    RECT 49.2000 71.1000 49.6000 73.9000 ;
	    RECT 53.6000 73.5000 53.9000 75.0000 ;
	    RECT 54.2000 74.8000 54.6000 75.2000 ;
	    RECT 52.7000 73.2000 53.9000 73.5000 ;
	    RECT 51.8000 72.4000 52.2000 73.2000 ;
	    RECT 52.7000 72.1000 53.0000 73.2000 ;
	    RECT 54.3000 73.1000 54.6000 74.8000 ;
	    RECT 52.6000 71.1000 53.0000 72.1000 ;
	    RECT 54.2000 71.1000 54.6000 73.1000 ;
	    RECT 55.0000 75.9000 55.4000 79.9000 ;
	    RECT 56.6000 76.2000 57.0000 79.9000 ;
	    RECT 57.4000 77.9000 57.8000 79.9000 ;
	    RECT 57.5000 77.8000 57.8000 77.9000 ;
	    RECT 59.0000 77.9000 59.4000 79.9000 ;
	    RECT 62.2000 77.9000 62.6000 79.9000 ;
	    RECT 59.0000 77.8000 59.3000 77.9000 ;
	    RECT 57.5000 77.5000 59.3000 77.8000 ;
	    RECT 62.3000 77.8000 62.6000 77.9000 ;
	    RECT 63.8000 77.9000 64.2000 79.9000 ;
	    RECT 63.8000 77.8000 64.1000 77.9000 ;
	    RECT 62.3000 77.5000 64.1000 77.8000 ;
	    RECT 57.5000 76.2000 57.8000 77.5000 ;
	    RECT 58.2000 76.4000 58.6000 77.2000 ;
	    RECT 62.3000 76.2000 62.6000 77.5000 ;
	    RECT 63.0000 76.4000 63.4000 77.2000 ;
	    RECT 55.9000 75.9000 57.0000 76.2000 ;
	    RECT 55.0000 74.8000 55.3000 75.9000 ;
	    RECT 55.9000 75.6000 56.2000 75.9000 ;
	    RECT 57.4000 75.8000 57.8000 76.2000 ;
	    RECT 62.2000 75.8000 62.6000 76.2000 ;
	    RECT 65.4000 76.2000 65.8000 79.9000 ;
	    RECT 65.4000 75.9000 66.5000 76.2000 ;
	    RECT 67.0000 75.9000 67.4000 79.9000 ;
	    RECT 67.8000 77.9000 68.2000 79.9000 ;
	    RECT 67.9000 77.8000 68.2000 77.9000 ;
	    RECT 69.4000 77.9000 69.8000 79.9000 ;
	    RECT 71.0000 77.9000 71.4000 79.9000 ;
	    RECT 69.4000 77.8000 69.7000 77.9000 ;
	    RECT 67.9000 77.5000 69.7000 77.8000 ;
	    RECT 71.1000 77.8000 71.4000 77.9000 ;
	    RECT 72.6000 77.9000 73.0000 79.9000 ;
	    RECT 72.6000 77.8000 72.9000 77.9000 ;
	    RECT 71.1000 77.5000 72.9000 77.8000 ;
	    RECT 67.9000 76.2000 68.2000 77.5000 ;
	    RECT 68.6000 76.4000 69.0000 77.2000 ;
	    RECT 71.1000 76.2000 71.4000 77.5000 ;
	    RECT 71.8000 76.4000 72.2000 77.2000 ;
	    RECT 74.5000 76.2000 74.9000 79.9000 ;
	    RECT 55.6000 75.2000 56.2000 75.6000 ;
	    RECT 55.0000 71.1000 55.4000 74.8000 ;
	    RECT 55.9000 73.7000 56.2000 75.2000 ;
	    RECT 57.5000 74.2000 57.8000 75.8000 ;
	    RECT 58.6000 74.8000 59.4000 75.2000 ;
	    RECT 62.3000 74.2000 62.6000 75.8000 ;
	    RECT 66.2000 75.6000 66.5000 75.9000 ;
	    RECT 66.2000 75.2000 66.8000 75.6000 ;
	    RECT 63.4000 74.8000 64.2000 75.2000 ;
	    RECT 57.5000 74.1000 58.3000 74.2000 ;
	    RECT 62.3000 74.1000 63.1000 74.2000 ;
	    RECT 57.5000 73.9000 58.4000 74.1000 ;
	    RECT 62.3000 73.9000 63.2000 74.1000 ;
	    RECT 55.9000 73.4000 57.0000 73.7000 ;
	    RECT 56.6000 71.1000 57.0000 73.4000 ;
	    RECT 58.0000 71.1000 58.4000 73.9000 ;
	    RECT 62.8000 71.1000 63.2000 73.9000 ;
	    RECT 66.2000 73.7000 66.5000 75.2000 ;
	    RECT 67.1000 74.8000 67.4000 75.9000 ;
	    RECT 67.8000 75.8000 68.2000 76.2000 ;
	    RECT 65.4000 73.4000 66.5000 73.7000 ;
	    RECT 65.4000 71.1000 65.8000 73.4000 ;
	    RECT 67.0000 71.1000 67.4000 74.8000 ;
	    RECT 67.9000 74.2000 68.2000 75.8000 ;
	    RECT 70.2000 75.4000 70.6000 76.2000 ;
	    RECT 71.0000 75.8000 71.4000 76.2000 ;
	    RECT 69.0000 74.8000 69.8000 75.2000 ;
	    RECT 71.1000 74.2000 71.4000 75.8000 ;
	    RECT 74.2000 75.9000 74.9000 76.2000 ;
	    RECT 74.2000 75.2000 74.5000 75.9000 ;
	    RECT 76.6000 75.6000 77.0000 79.9000 ;
	    RECT 75.0000 75.4000 77.0000 75.6000 ;
	    RECT 74.9000 75.3000 77.0000 75.4000 ;
	    RECT 77.4000 75.6000 77.8000 79.9000 ;
	    RECT 79.5000 76.2000 79.9000 79.9000 ;
	    RECT 81.4000 77.9000 81.8000 79.9000 ;
	    RECT 81.5000 77.8000 81.8000 77.9000 ;
	    RECT 83.0000 77.9000 83.4000 79.9000 ;
	    RECT 83.0000 77.8000 83.3000 77.9000 ;
	    RECT 81.5000 77.5000 83.3000 77.8000 ;
	    RECT 82.2000 76.4000 82.6000 77.2000 ;
	    RECT 83.0000 76.2000 83.3000 77.5000 ;
	    RECT 79.5000 75.9000 80.2000 76.2000 ;
	    RECT 77.4000 75.4000 79.4000 75.6000 ;
	    RECT 77.4000 75.3000 79.5000 75.4000 ;
	    RECT 72.2000 74.8000 73.0000 75.2000 ;
	    RECT 74.2000 74.8000 74.6000 75.2000 ;
	    RECT 74.9000 75.0000 75.3000 75.3000 ;
	    RECT 79.1000 75.0000 79.5000 75.3000 ;
	    RECT 79.9000 75.2000 80.2000 75.9000 ;
	    RECT 83.0000 75.8000 83.4000 76.2000 ;
	    RECT 67.9000 74.1000 68.7000 74.2000 ;
	    RECT 71.1000 74.1000 71.9000 74.2000 ;
	    RECT 67.9000 73.9000 68.8000 74.1000 ;
	    RECT 71.1000 73.9000 72.0000 74.1000 ;
	    RECT 68.4000 71.1000 68.8000 73.9000 ;
	    RECT 71.6000 71.1000 72.0000 73.9000 ;
	    RECT 74.2000 73.1000 74.5000 74.8000 ;
	    RECT 74.9000 73.5000 75.2000 75.0000 ;
	    RECT 79.2000 73.5000 79.5000 75.0000 ;
	    RECT 79.8000 74.8000 80.2000 75.2000 ;
	    RECT 81.4000 74.8000 82.2000 75.2000 ;
	    RECT 74.9000 73.2000 76.1000 73.5000 ;
	    RECT 78.3000 73.2000 79.5000 73.5000 ;
	    RECT 74.2000 71.1000 74.6000 73.1000 ;
	    RECT 75.8000 72.1000 76.1000 73.2000 ;
	    RECT 76.6000 73.1000 77.0000 73.2000 ;
	    RECT 77.4000 73.1000 77.8000 73.2000 ;
	    RECT 76.6000 72.8000 77.8000 73.1000 ;
	    RECT 76.6000 72.4000 77.0000 72.8000 ;
	    RECT 77.4000 72.4000 77.8000 72.8000 ;
	    RECT 78.3000 72.1000 78.6000 73.2000 ;
	    RECT 79.9000 73.1000 80.2000 74.8000 ;
	    RECT 83.0000 74.2000 83.3000 75.8000 ;
	    RECT 82.5000 74.1000 83.3000 74.2000 ;
	    RECT 75.8000 71.1000 76.2000 72.1000 ;
	    RECT 78.2000 71.1000 78.6000 72.1000 ;
	    RECT 79.8000 71.1000 80.2000 73.1000 ;
	    RECT 82.4000 73.9000 83.3000 74.1000 ;
	    RECT 82.4000 71.1000 82.8000 73.9000 ;
	    RECT 84.6000 71.1000 85.0000 79.9000 ;
	    RECT 86.2000 71.1000 86.6000 79.9000 ;
	    RECT 87.0000 75.9000 87.4000 79.9000 ;
	    RECT 88.6000 77.9000 89.0000 79.9000 ;
	    RECT 91.0000 77.9000 91.4000 79.9000 ;
	    RECT 87.0000 75.2000 87.3000 75.9000 ;
	    RECT 88.6000 75.8000 88.9000 77.9000 ;
	    RECT 87.7000 75.5000 88.9000 75.8000 ;
	    RECT 91.1000 75.8000 91.4000 77.9000 ;
	    RECT 92.6000 75.9000 93.0000 79.9000 ;
	    RECT 93.4000 77.9000 93.8000 79.9000 ;
	    RECT 93.5000 77.8000 93.8000 77.9000 ;
	    RECT 95.0000 77.9000 95.4000 79.9000 ;
	    RECT 95.0000 77.8000 95.3000 77.9000 ;
	    RECT 93.5000 77.5000 95.3000 77.8000 ;
	    RECT 93.5000 76.2000 93.8000 77.5000 ;
	    RECT 95.0000 77.2000 95.3000 77.5000 ;
	    RECT 94.2000 76.4000 94.6000 77.2000 ;
	    RECT 95.0000 76.8000 95.4000 77.2000 ;
	    RECT 96.6000 76.2000 97.0000 79.9000 ;
	    RECT 98.2000 76.2000 98.6000 79.9000 ;
	    RECT 91.1000 75.5000 92.3000 75.8000 ;
	    RECT 87.0000 74.8000 87.4000 75.2000 ;
	    RECT 87.0000 73.1000 87.3000 74.8000 ;
	    RECT 87.7000 73.8000 88.0000 75.5000 ;
	    RECT 88.6000 74.8000 89.0000 75.2000 ;
	    RECT 91.0000 74.8000 91.4000 75.2000 ;
	    RECT 88.6000 74.4000 88.9000 74.8000 ;
	    RECT 88.4000 74.0000 89.0000 74.4000 ;
	    RECT 89.4000 74.1000 89.8000 74.6000 ;
	    RECT 90.2000 74.1000 90.6000 74.6000 ;
	    RECT 91.1000 74.4000 91.4000 74.8000 ;
	    RECT 91.1000 74.1000 91.6000 74.4000 ;
	    RECT 89.4000 73.8000 90.6000 74.1000 ;
	    RECT 91.2000 74.0000 91.6000 74.1000 ;
	    RECT 92.0000 73.8000 92.3000 75.5000 ;
	    RECT 92.7000 75.2000 93.0000 75.9000 ;
	    RECT 93.4000 75.8000 93.8000 76.2000 ;
	    RECT 92.6000 74.8000 93.0000 75.2000 ;
	    RECT 87.6000 73.7000 88.0000 73.8000 ;
	    RECT 92.0000 73.7000 92.4000 73.8000 ;
	    RECT 87.6000 73.5000 89.1000 73.7000 ;
	    RECT 90.9000 73.5000 92.4000 73.7000 ;
	    RECT 87.6000 73.4000 89.7000 73.5000 ;
	    RECT 88.8000 73.2000 89.7000 73.4000 ;
	    RECT 89.4000 73.1000 89.7000 73.2000 ;
	    RECT 90.3000 73.4000 92.4000 73.5000 ;
	    RECT 90.3000 73.2000 91.2000 73.4000 ;
	    RECT 90.3000 73.1000 90.6000 73.2000 ;
	    RECT 92.7000 73.1000 93.0000 74.8000 ;
	    RECT 93.5000 74.2000 93.8000 75.8000 ;
	    RECT 95.8000 75.4000 96.2000 76.2000 ;
	    RECT 96.6000 75.9000 98.6000 76.2000 ;
	    RECT 99.0000 75.9000 99.4000 79.9000 ;
	    RECT 99.8000 76.2000 100.2000 79.9000 ;
	    RECT 101.4000 76.2000 101.8000 79.9000 ;
	    RECT 99.8000 75.9000 101.8000 76.2000 ;
	    RECT 102.2000 75.9000 102.6000 79.9000 ;
	    RECT 97.0000 75.2000 97.4000 75.4000 ;
	    RECT 99.0000 75.2000 99.3000 75.9000 ;
	    RECT 100.2000 75.2000 100.6000 75.4000 ;
	    RECT 102.2000 75.2000 102.5000 75.9000 ;
	    RECT 103.8000 75.6000 104.2000 79.9000 ;
	    RECT 105.4000 75.6000 105.8000 79.9000 ;
	    RECT 107.0000 75.6000 107.4000 79.9000 ;
	    RECT 108.6000 75.6000 109.0000 79.9000 ;
	    RECT 103.0000 75.2000 104.2000 75.6000 ;
	    RECT 104.7000 75.2000 105.8000 75.6000 ;
	    RECT 106.3000 75.2000 107.4000 75.6000 ;
	    RECT 108.1000 75.2000 109.0000 75.6000 ;
	    RECT 110.2000 75.9000 110.6000 79.9000 ;
	    RECT 111.8000 76.2000 112.2000 79.9000 ;
	    RECT 111.1000 75.9000 112.2000 76.2000 ;
	    RECT 94.6000 74.8000 95.4000 75.2000 ;
	    RECT 96.6000 74.9000 97.4000 75.2000 ;
	    RECT 98.2000 74.9000 99.4000 75.2000 ;
	    RECT 96.6000 74.8000 97.0000 74.9000 ;
	    RECT 93.5000 74.1000 94.3000 74.2000 ;
	    RECT 93.5000 73.9000 94.4000 74.1000 ;
	    RECT 87.0000 72.6000 87.7000 73.1000 ;
	    RECT 87.3000 71.1000 87.7000 72.6000 ;
	    RECT 89.4000 71.1000 89.8000 73.1000 ;
	    RECT 90.2000 71.1000 90.6000 73.1000 ;
	    RECT 92.3000 72.6000 93.0000 73.1000 ;
	    RECT 92.3000 71.1000 92.7000 72.6000 ;
	    RECT 94.0000 71.1000 94.4000 73.9000 ;
	    RECT 97.4000 73.8000 97.8000 74.6000 ;
	    RECT 98.2000 73.1000 98.5000 74.9000 ;
	    RECT 99.0000 74.8000 99.4000 74.9000 ;
	    RECT 99.8000 74.9000 100.6000 75.2000 ;
	    RECT 101.4000 74.9000 102.6000 75.2000 ;
	    RECT 99.8000 74.8000 100.2000 74.9000 ;
	    RECT 100.6000 73.8000 101.0000 74.6000 ;
	    RECT 98.2000 71.1000 98.6000 73.1000 ;
	    RECT 99.0000 72.8000 99.4000 73.2000 ;
	    RECT 101.4000 73.1000 101.7000 74.9000 ;
	    RECT 102.2000 74.8000 102.6000 74.9000 ;
	    RECT 103.0000 73.8000 103.4000 75.2000 ;
	    RECT 104.7000 74.5000 105.1000 75.2000 ;
	    RECT 106.3000 74.5000 106.7000 75.2000 ;
	    RECT 108.1000 74.5000 108.5000 75.2000 ;
	    RECT 103.8000 74.1000 105.1000 74.5000 ;
	    RECT 105.5000 74.1000 106.7000 74.5000 ;
	    RECT 107.2000 74.1000 108.5000 74.5000 ;
	    RECT 104.7000 73.8000 105.1000 74.1000 ;
	    RECT 106.3000 73.8000 106.7000 74.1000 ;
	    RECT 108.1000 73.8000 108.5000 74.1000 ;
	    RECT 110.2000 74.8000 110.5000 75.9000 ;
	    RECT 111.1000 75.6000 111.4000 75.9000 ;
	    RECT 110.8000 75.2000 111.4000 75.6000 ;
	    RECT 114.2000 75.7000 114.6000 79.9000 ;
	    RECT 116.4000 78.2000 116.8000 79.9000 ;
	    RECT 115.8000 77.9000 116.8000 78.2000 ;
	    RECT 118.6000 77.9000 119.0000 79.9000 ;
	    RECT 120.7000 77.9000 121.3000 79.9000 ;
	    RECT 115.8000 77.5000 116.2000 77.9000 ;
	    RECT 118.6000 77.6000 118.9000 77.9000 ;
	    RECT 117.5000 77.3000 119.3000 77.6000 ;
	    RECT 120.6000 77.5000 121.0000 77.9000 ;
	    RECT 117.5000 77.2000 117.9000 77.3000 ;
	    RECT 118.9000 77.2000 119.3000 77.3000 ;
	    RECT 115.8000 76.5000 116.2000 76.6000 ;
	    RECT 118.1000 76.5000 118.5000 76.6000 ;
	    RECT 115.8000 76.2000 118.5000 76.5000 ;
	    RECT 118.8000 76.5000 119.9000 76.8000 ;
	    RECT 118.8000 75.9000 119.1000 76.5000 ;
	    RECT 119.5000 76.4000 119.9000 76.5000 ;
	    RECT 120.7000 76.6000 121.4000 77.0000 ;
	    RECT 120.7000 76.1000 121.0000 76.6000 ;
	    RECT 116.7000 75.7000 119.1000 75.9000 ;
	    RECT 114.2000 75.6000 119.1000 75.7000 ;
	    RECT 119.8000 75.8000 121.0000 76.1000 ;
	    RECT 123.0000 76.1000 123.4000 79.9000 ;
	    RECT 124.6000 77.9000 125.0000 79.9000 ;
	    RECT 123.8000 76.1000 124.2000 76.2000 ;
	    RECT 123.0000 75.8000 124.2000 76.1000 ;
	    RECT 124.7000 75.8000 125.0000 77.9000 ;
	    RECT 126.2000 75.9000 126.6000 79.9000 ;
	    RECT 114.2000 75.5000 117.1000 75.6000 ;
	    RECT 114.2000 75.4000 117.0000 75.5000 ;
	    RECT 103.0000 73.4000 104.2000 73.8000 ;
	    RECT 104.7000 73.4000 105.8000 73.8000 ;
	    RECT 106.3000 73.4000 107.4000 73.8000 ;
	    RECT 108.1000 73.4000 109.0000 73.8000 ;
	    RECT 98.9000 72.4000 99.3000 72.8000 ;
	    RECT 101.4000 71.1000 101.8000 73.1000 ;
	    RECT 102.2000 72.8000 102.6000 73.2000 ;
	    RECT 102.1000 72.4000 102.5000 72.8000 ;
	    RECT 103.8000 71.1000 104.2000 73.4000 ;
	    RECT 105.4000 71.1000 105.8000 73.4000 ;
	    RECT 107.0000 71.1000 107.4000 73.4000 ;
	    RECT 108.6000 71.1000 109.0000 73.4000 ;
	    RECT 110.2000 71.1000 110.6000 74.8000 ;
	    RECT 111.1000 73.7000 111.4000 75.2000 ;
	    RECT 117.4000 75.1000 117.8000 75.2000 ;
	    RECT 115.3000 74.8000 117.8000 75.1000 ;
	    RECT 115.3000 74.7000 115.7000 74.8000 ;
	    RECT 116.6000 74.7000 117.0000 74.8000 ;
	    RECT 116.1000 74.2000 116.5000 74.3000 ;
	    RECT 119.8000 74.2000 120.1000 75.8000 ;
	    RECT 123.0000 75.6000 123.4000 75.8000 ;
	    RECT 121.3000 75.3000 123.4000 75.6000 ;
	    RECT 124.7000 75.5000 125.9000 75.8000 ;
	    RECT 121.3000 75.2000 121.7000 75.3000 ;
	    RECT 122.1000 74.9000 122.5000 75.0000 ;
	    RECT 120.6000 74.6000 122.5000 74.9000 ;
	    RECT 120.6000 74.5000 121.0000 74.6000 ;
	    RECT 114.6000 73.9000 120.1000 74.2000 ;
	    RECT 114.6000 73.8000 115.4000 73.9000 ;
	    RECT 111.1000 73.4000 112.2000 73.7000 ;
	    RECT 111.8000 71.1000 112.2000 73.4000 ;
	    RECT 114.2000 71.1000 114.6000 73.5000 ;
	    RECT 116.7000 72.8000 117.0000 73.9000 ;
	    RECT 118.2000 73.8000 118.6000 73.9000 ;
	    RECT 119.5000 73.8000 119.9000 73.9000 ;
	    RECT 123.0000 73.6000 123.4000 75.3000 ;
	    RECT 124.6000 74.8000 125.0000 75.2000 ;
	    RECT 123.8000 73.8000 124.2000 74.6000 ;
	    RECT 124.7000 74.4000 125.0000 74.8000 ;
	    RECT 124.7000 74.1000 125.2000 74.4000 ;
	    RECT 124.8000 74.0000 125.2000 74.1000 ;
	    RECT 125.6000 73.8000 125.9000 75.5000 ;
	    RECT 126.3000 75.2000 126.6000 75.9000 ;
	    RECT 127.0000 75.7000 127.4000 79.9000 ;
	    RECT 129.2000 78.2000 129.6000 79.9000 ;
	    RECT 128.6000 77.9000 129.6000 78.2000 ;
	    RECT 131.4000 77.9000 131.8000 79.9000 ;
	    RECT 133.5000 77.9000 134.1000 79.9000 ;
	    RECT 128.6000 77.5000 129.0000 77.9000 ;
	    RECT 131.4000 77.6000 131.7000 77.9000 ;
	    RECT 130.3000 77.3000 132.1000 77.6000 ;
	    RECT 133.4000 77.5000 133.8000 77.9000 ;
	    RECT 130.3000 77.2000 130.7000 77.3000 ;
	    RECT 131.7000 77.2000 132.1000 77.3000 ;
	    RECT 128.6000 76.5000 129.0000 76.6000 ;
	    RECT 130.9000 76.5000 131.3000 76.6000 ;
	    RECT 128.6000 76.2000 131.3000 76.5000 ;
	    RECT 131.6000 76.5000 132.7000 76.8000 ;
	    RECT 131.6000 75.9000 131.9000 76.5000 ;
	    RECT 132.3000 76.4000 132.7000 76.5000 ;
	    RECT 133.5000 76.6000 134.2000 77.0000 ;
	    RECT 133.5000 76.1000 133.8000 76.6000 ;
	    RECT 129.5000 75.7000 131.9000 75.9000 ;
	    RECT 127.0000 75.6000 131.9000 75.7000 ;
	    RECT 132.6000 75.8000 133.8000 76.1000 ;
	    RECT 127.0000 75.5000 129.9000 75.6000 ;
	    RECT 127.0000 75.4000 129.8000 75.5000 ;
	    RECT 126.2000 74.8000 126.6000 75.2000 ;
	    RECT 130.2000 75.1000 130.6000 75.2000 ;
	    RECT 125.6000 73.7000 126.0000 73.8000 ;
	    RECT 121.5000 73.3000 123.4000 73.6000 ;
	    RECT 124.5000 73.5000 126.0000 73.7000 ;
	    RECT 121.5000 73.2000 121.9000 73.3000 ;
	    RECT 115.8000 72.1000 116.2000 72.5000 ;
	    RECT 116.6000 72.4000 117.0000 72.8000 ;
	    RECT 117.5000 72.7000 117.9000 72.8000 ;
	    RECT 117.5000 72.4000 118.9000 72.7000 ;
	    RECT 118.6000 72.1000 118.9000 72.4000 ;
	    RECT 120.6000 72.1000 121.0000 72.5000 ;
	    RECT 115.8000 71.8000 116.8000 72.1000 ;
	    RECT 116.4000 71.1000 116.8000 71.8000 ;
	    RECT 118.6000 71.1000 119.0000 72.1000 ;
	    RECT 120.6000 71.8000 121.3000 72.1000 ;
	    RECT 120.7000 71.1000 121.3000 71.8000 ;
	    RECT 123.0000 71.1000 123.4000 73.3000 ;
	    RECT 123.9000 73.4000 126.0000 73.5000 ;
	    RECT 123.9000 73.2000 124.8000 73.4000 ;
	    RECT 123.9000 73.1000 124.2000 73.2000 ;
	    RECT 126.3000 73.1000 126.6000 74.8000 ;
	    RECT 128.1000 74.8000 130.6000 75.1000 ;
	    RECT 128.1000 74.7000 128.5000 74.8000 ;
	    RECT 129.4000 74.7000 129.8000 74.8000 ;
	    RECT 128.9000 74.2000 129.3000 74.3000 ;
	    RECT 132.6000 74.2000 132.9000 75.8000 ;
	    RECT 135.8000 75.6000 136.2000 79.9000 ;
	    RECT 136.6000 76.2000 137.0000 79.9000 ;
	    RECT 138.2000 76.2000 138.6000 79.9000 ;
	    RECT 136.6000 75.9000 138.6000 76.2000 ;
	    RECT 139.0000 75.9000 139.4000 79.9000 ;
	    RECT 139.8000 76.2000 140.2000 79.9000 ;
	    RECT 139.8000 75.9000 140.9000 76.2000 ;
	    RECT 141.4000 75.9000 141.8000 79.9000 ;
	    RECT 134.1000 75.3000 136.2000 75.6000 ;
	    RECT 134.1000 75.2000 134.5000 75.3000 ;
	    RECT 134.9000 74.9000 135.3000 75.0000 ;
	    RECT 133.4000 74.6000 135.3000 74.9000 ;
	    RECT 133.4000 74.5000 133.8000 74.6000 ;
	    RECT 127.4000 73.9000 132.9000 74.2000 ;
	    RECT 127.4000 73.8000 128.2000 73.9000 ;
	    RECT 123.8000 71.1000 124.2000 73.1000 ;
	    RECT 125.9000 72.6000 126.6000 73.1000 ;
	    RECT 125.9000 71.1000 126.3000 72.6000 ;
	    RECT 127.0000 71.1000 127.4000 73.5000 ;
	    RECT 129.5000 72.8000 129.8000 73.9000 ;
	    RECT 132.3000 73.8000 132.7000 73.9000 ;
	    RECT 135.8000 73.6000 136.2000 75.3000 ;
	    RECT 137.0000 75.2000 137.4000 75.4000 ;
	    RECT 139.0000 75.2000 139.3000 75.9000 ;
	    RECT 140.6000 75.6000 140.9000 75.9000 ;
	    RECT 140.6000 75.2000 141.2000 75.6000 ;
	    RECT 136.6000 74.9000 137.4000 75.2000 ;
	    RECT 138.2000 74.9000 139.4000 75.2000 ;
	    RECT 136.6000 74.8000 137.0000 74.9000 ;
	    RECT 137.4000 73.8000 137.8000 74.6000 ;
	    RECT 134.3000 73.3000 136.2000 73.6000 ;
	    RECT 134.3000 73.2000 134.7000 73.3000 ;
	    RECT 128.6000 72.1000 129.0000 72.5000 ;
	    RECT 129.4000 72.4000 129.8000 72.8000 ;
	    RECT 130.3000 72.7000 130.7000 72.8000 ;
	    RECT 130.3000 72.4000 131.7000 72.7000 ;
	    RECT 131.4000 72.1000 131.7000 72.4000 ;
	    RECT 133.4000 72.1000 133.8000 72.5000 ;
	    RECT 128.6000 71.8000 129.6000 72.1000 ;
	    RECT 129.2000 71.1000 129.6000 71.8000 ;
	    RECT 131.4000 71.1000 131.8000 72.1000 ;
	    RECT 133.4000 71.8000 134.1000 72.1000 ;
	    RECT 133.5000 71.1000 134.1000 71.8000 ;
	    RECT 135.8000 71.1000 136.2000 73.3000 ;
	    RECT 138.2000 73.1000 138.5000 74.9000 ;
	    RECT 139.0000 74.8000 139.4000 74.9000 ;
	    RECT 140.6000 73.7000 140.9000 75.2000 ;
	    RECT 141.5000 74.8000 141.8000 75.9000 ;
	    RECT 139.8000 73.4000 140.9000 73.7000 ;
	    RECT 141.4000 74.1000 141.8000 74.8000 ;
	    RECT 142.2000 74.1000 142.6000 74.2000 ;
	    RECT 141.4000 73.8000 142.6000 74.1000 ;
	    RECT 138.2000 71.1000 138.6000 73.1000 ;
	    RECT 139.0000 72.8000 139.4000 73.2000 ;
	    RECT 138.9000 72.4000 139.3000 72.8000 ;
	    RECT 139.8000 71.1000 140.2000 73.4000 ;
	    RECT 141.4000 71.1000 141.8000 73.8000 ;
	    RECT 142.2000 73.4000 142.6000 73.8000 ;
	    RECT 143.0000 71.1000 143.4000 79.9000 ;
	    RECT 143.8000 76.2000 144.2000 79.9000 ;
	    RECT 145.4000 76.2000 145.8000 79.9000 ;
	    RECT 143.8000 75.9000 145.8000 76.2000 ;
	    RECT 146.2000 75.8000 146.6000 79.9000 ;
	    RECT 147.0000 76.2000 147.4000 79.9000 ;
	    RECT 148.6000 76.2000 149.0000 79.9000 ;
	    RECT 147.0000 75.9000 149.0000 76.2000 ;
	    RECT 149.4000 75.9000 149.8000 79.9000 ;
	    RECT 150.2000 75.9000 150.6000 79.9000 ;
	    RECT 151.0000 76.2000 151.4000 79.9000 ;
	    RECT 152.6000 76.2000 153.0000 79.9000 ;
	    RECT 151.0000 75.9000 153.0000 76.2000 ;
	    RECT 144.2000 75.2000 144.6000 75.4000 ;
	    RECT 146.2000 75.2000 146.5000 75.8000 ;
	    RECT 147.4000 75.2000 147.8000 75.4000 ;
	    RECT 149.4000 75.2000 149.7000 75.9000 ;
	    RECT 150.3000 75.2000 150.6000 75.9000 ;
	    RECT 153.4000 75.7000 153.8000 79.9000 ;
	    RECT 155.6000 78.2000 156.0000 79.9000 ;
	    RECT 155.0000 77.9000 156.0000 78.2000 ;
	    RECT 157.8000 77.9000 158.2000 79.9000 ;
	    RECT 159.9000 77.9000 160.5000 79.9000 ;
	    RECT 155.0000 77.5000 155.4000 77.9000 ;
	    RECT 157.8000 77.6000 158.1000 77.9000 ;
	    RECT 156.7000 77.3000 158.5000 77.6000 ;
	    RECT 159.8000 77.5000 160.2000 77.9000 ;
	    RECT 156.7000 77.2000 157.1000 77.3000 ;
	    RECT 158.1000 77.2000 158.5000 77.3000 ;
	    RECT 155.0000 76.5000 155.4000 76.6000 ;
	    RECT 157.3000 76.5000 157.7000 76.6000 ;
	    RECT 155.0000 76.2000 157.7000 76.5000 ;
	    RECT 158.0000 76.5000 159.1000 76.8000 ;
	    RECT 158.0000 75.9000 158.3000 76.5000 ;
	    RECT 158.7000 76.4000 159.1000 76.5000 ;
	    RECT 159.9000 76.6000 160.6000 77.0000 ;
	    RECT 159.9000 76.1000 160.2000 76.6000 ;
	    RECT 155.9000 75.7000 158.3000 75.9000 ;
	    RECT 153.4000 75.6000 158.3000 75.7000 ;
	    RECT 159.0000 75.8000 160.2000 76.1000 ;
	    RECT 153.4000 75.5000 156.3000 75.6000 ;
	    RECT 153.4000 75.4000 156.2000 75.5000 ;
	    RECT 152.2000 75.2000 152.6000 75.4000 ;
	    RECT 159.0000 75.2000 159.3000 75.8000 ;
	    RECT 162.2000 75.6000 162.6000 79.9000 ;
	    RECT 160.5000 75.3000 162.6000 75.6000 ;
	    RECT 163.0000 75.7000 163.4000 79.9000 ;
	    RECT 165.2000 78.2000 165.6000 79.9000 ;
	    RECT 164.6000 77.9000 165.6000 78.2000 ;
	    RECT 167.4000 77.9000 167.8000 79.9000 ;
	    RECT 169.5000 77.9000 170.1000 79.9000 ;
	    RECT 164.6000 77.5000 165.0000 77.9000 ;
	    RECT 167.4000 77.6000 167.7000 77.9000 ;
	    RECT 166.3000 77.3000 168.1000 77.6000 ;
	    RECT 169.4000 77.5000 169.8000 77.9000 ;
	    RECT 166.3000 77.2000 166.7000 77.3000 ;
	    RECT 167.7000 77.2000 168.1000 77.3000 ;
	    RECT 164.6000 76.5000 165.0000 76.6000 ;
	    RECT 166.9000 76.5000 167.3000 76.6000 ;
	    RECT 164.6000 76.2000 167.3000 76.5000 ;
	    RECT 167.6000 76.5000 168.7000 76.8000 ;
	    RECT 167.6000 75.9000 167.9000 76.5000 ;
	    RECT 168.3000 76.4000 168.7000 76.5000 ;
	    RECT 169.5000 76.6000 170.2000 77.0000 ;
	    RECT 169.5000 76.1000 169.8000 76.6000 ;
	    RECT 165.5000 75.7000 167.9000 75.9000 ;
	    RECT 163.0000 75.6000 167.9000 75.7000 ;
	    RECT 168.6000 75.8000 169.8000 76.1000 ;
	    RECT 163.0000 75.5000 165.9000 75.6000 ;
	    RECT 163.0000 75.4000 165.8000 75.5000 ;
	    RECT 160.5000 75.2000 160.9000 75.3000 ;
	    RECT 143.8000 74.9000 144.6000 75.2000 ;
	    RECT 145.4000 74.9000 146.6000 75.2000 ;
	    RECT 143.8000 74.8000 144.2000 74.9000 ;
	    RECT 143.8000 74.1000 144.2000 74.2000 ;
	    RECT 144.6000 74.1000 145.0000 74.6000 ;
	    RECT 143.8000 73.8000 145.0000 74.1000 ;
	    RECT 145.4000 73.1000 145.7000 74.9000 ;
	    RECT 146.2000 74.8000 146.6000 74.9000 ;
	    RECT 147.0000 74.9000 147.8000 75.2000 ;
	    RECT 148.6000 74.9000 149.8000 75.2000 ;
	    RECT 147.0000 74.8000 147.4000 74.9000 ;
	    RECT 147.8000 73.8000 148.2000 74.6000 ;
	    RECT 145.4000 71.1000 145.8000 73.1000 ;
	    RECT 146.2000 72.8000 146.6000 73.2000 ;
	    RECT 148.6000 73.1000 148.9000 74.9000 ;
	    RECT 149.4000 74.8000 149.8000 74.9000 ;
	    RECT 150.2000 74.9000 151.4000 75.2000 ;
	    RECT 152.2000 74.9000 153.0000 75.2000 ;
	    RECT 156.6000 75.1000 157.0000 75.2000 ;
	    RECT 150.2000 74.8000 150.6000 74.9000 ;
	    RECT 149.4000 73.1000 149.8000 73.2000 ;
	    RECT 150.2000 73.1000 150.6000 73.2000 ;
	    RECT 151.1000 73.1000 151.4000 74.9000 ;
	    RECT 152.6000 74.8000 153.0000 74.9000 ;
	    RECT 154.5000 74.8000 157.0000 75.1000 ;
	    RECT 159.0000 74.8000 159.4000 75.2000 ;
	    RECT 161.3000 74.9000 161.7000 75.0000 ;
	    RECT 154.5000 74.7000 154.9000 74.8000 ;
	    RECT 155.8000 74.7000 156.2000 74.8000 ;
	    RECT 151.8000 73.8000 152.2000 74.6000 ;
	    RECT 155.3000 74.2000 155.7000 74.3000 ;
	    RECT 159.0000 74.2000 159.3000 74.8000 ;
	    RECT 159.8000 74.6000 161.7000 74.9000 ;
	    RECT 159.8000 74.5000 160.2000 74.6000 ;
	    RECT 153.8000 73.9000 159.3000 74.2000 ;
	    RECT 153.8000 73.8000 154.6000 73.9000 ;
	    RECT 146.1000 72.4000 146.5000 72.8000 ;
	    RECT 148.6000 71.1000 149.0000 73.1000 ;
	    RECT 149.4000 72.8000 150.6000 73.1000 ;
	    RECT 149.3000 72.4000 149.7000 72.8000 ;
	    RECT 150.3000 72.4000 150.7000 72.8000 ;
	    RECT 151.0000 71.1000 151.4000 73.1000 ;
	    RECT 153.4000 71.1000 153.8000 73.5000 ;
	    RECT 155.9000 72.8000 156.2000 73.9000 ;
	    RECT 158.7000 73.8000 159.1000 73.9000 ;
	    RECT 162.2000 73.6000 162.6000 75.3000 ;
	    RECT 166.2000 75.1000 166.6000 75.2000 ;
	    RECT 164.1000 74.8000 166.6000 75.1000 ;
	    RECT 164.1000 74.7000 164.5000 74.8000 ;
	    RECT 164.9000 74.2000 165.3000 74.3000 ;
	    RECT 168.6000 74.2000 168.9000 75.8000 ;
	    RECT 171.8000 75.6000 172.2000 79.9000 ;
	    RECT 170.1000 75.3000 172.2000 75.6000 ;
	    RECT 170.1000 75.2000 170.5000 75.3000 ;
	    RECT 170.9000 74.9000 171.3000 75.0000 ;
	    RECT 169.4000 74.6000 171.3000 74.9000 ;
	    RECT 169.4000 74.5000 169.8000 74.6000 ;
	    RECT 163.4000 73.9000 168.9000 74.2000 ;
	    RECT 163.4000 73.8000 164.2000 73.9000 ;
	    RECT 160.7000 73.3000 162.6000 73.6000 ;
	    RECT 160.7000 73.2000 161.1000 73.3000 ;
	    RECT 155.0000 72.1000 155.4000 72.5000 ;
	    RECT 155.8000 72.4000 156.2000 72.8000 ;
	    RECT 156.7000 72.7000 157.1000 72.8000 ;
	    RECT 156.7000 72.4000 158.1000 72.7000 ;
	    RECT 157.8000 72.1000 158.1000 72.4000 ;
	    RECT 159.8000 72.1000 160.2000 72.5000 ;
	    RECT 155.0000 71.8000 156.0000 72.1000 ;
	    RECT 155.6000 71.1000 156.0000 71.8000 ;
	    RECT 157.8000 71.1000 158.2000 72.1000 ;
	    RECT 159.8000 71.8000 160.5000 72.1000 ;
	    RECT 159.9000 71.1000 160.5000 71.8000 ;
	    RECT 162.2000 71.1000 162.6000 73.3000 ;
	    RECT 163.0000 71.1000 163.4000 73.5000 ;
	    RECT 165.5000 72.8000 165.8000 73.9000 ;
	    RECT 168.3000 73.8000 168.7000 73.9000 ;
	    RECT 171.8000 73.6000 172.2000 75.3000 ;
	    RECT 170.3000 73.3000 172.2000 73.6000 ;
	    RECT 170.3000 73.2000 170.7000 73.3000 ;
	    RECT 164.6000 72.1000 165.0000 72.5000 ;
	    RECT 165.4000 72.4000 165.8000 72.8000 ;
	    RECT 166.3000 72.7000 166.7000 72.8000 ;
	    RECT 166.3000 72.4000 167.7000 72.7000 ;
	    RECT 167.4000 72.1000 167.7000 72.4000 ;
	    RECT 169.4000 72.1000 169.8000 72.5000 ;
	    RECT 164.6000 71.8000 165.6000 72.1000 ;
	    RECT 165.2000 71.1000 165.6000 71.8000 ;
	    RECT 167.4000 71.1000 167.8000 72.1000 ;
	    RECT 169.4000 71.8000 170.1000 72.1000 ;
	    RECT 169.5000 71.1000 170.1000 71.8000 ;
	    RECT 171.8000 71.1000 172.2000 73.3000 ;
	    RECT 1.2000 67.1000 1.6000 69.9000 ;
	    RECT 0.7000 66.9000 1.6000 67.1000 ;
	    RECT 0.7000 66.8000 1.5000 66.9000 ;
	    RECT 0.7000 65.2000 1.0000 66.8000 ;
	    RECT 1.8000 65.8000 2.6000 66.2000 ;
	    RECT 0.6000 64.8000 1.0000 65.2000 ;
	    RECT 3.0000 64.8000 3.4000 65.6000 ;
	    RECT 0.7000 63.5000 1.0000 64.8000 ;
	    RECT 1.4000 63.8000 1.8000 64.6000 ;
	    RECT 0.7000 63.2000 2.5000 63.5000 ;
	    RECT 0.7000 63.1000 1.0000 63.2000 ;
	    RECT 0.6000 61.1000 1.0000 63.1000 ;
	    RECT 2.2000 63.1000 2.5000 63.2000 ;
	    RECT 2.2000 61.1000 2.6000 63.1000 ;
	    RECT 4.6000 61.1000 5.0000 69.9000 ;
	    RECT 6.2000 68.9000 6.6000 69.9000 ;
	    RECT 5.4000 67.8000 5.8000 68.6000 ;
	    RECT 6.3000 67.8000 6.6000 68.9000 ;
	    RECT 7.8000 67.9000 8.2000 69.9000 ;
	    RECT 6.3000 67.5000 7.5000 67.8000 ;
	    RECT 7.2000 66.0000 7.5000 67.5000 ;
	    RECT 7.9000 67.2000 8.2000 67.9000 ;
	    RECT 7.8000 66.8000 8.2000 67.2000 ;
	    RECT 10.4000 67.1000 10.8000 69.9000 ;
	    RECT 13.6000 67.1000 14.0000 69.9000 ;
	    RECT 15.6000 67.1000 16.0000 69.9000 ;
	    RECT 10.4000 66.9000 11.3000 67.1000 ;
	    RECT 13.6000 66.9000 14.5000 67.1000 ;
	    RECT 10.5000 66.8000 11.3000 66.9000 ;
	    RECT 13.7000 66.8000 14.5000 66.9000 ;
	    RECT 7.9000 66.2000 8.2000 66.8000 ;
	    RECT 7.1000 65.7000 7.5000 66.0000 ;
	    RECT 7.8000 65.8000 8.2000 66.2000 ;
	    RECT 9.4000 65.8000 10.2000 66.2000 ;
	    RECT 5.4000 65.6000 7.5000 65.7000 ;
	    RECT 5.4000 65.4000 7.4000 65.6000 ;
	    RECT 5.4000 61.1000 5.8000 65.4000 ;
	    RECT 7.9000 65.1000 8.2000 65.8000 ;
	    RECT 7.5000 64.8000 8.2000 65.1000 ;
	    RECT 8.6000 64.8000 9.0000 65.6000 ;
	    RECT 11.0000 65.2000 11.3000 66.8000 ;
	    RECT 12.6000 65.8000 13.4000 66.2000 ;
	    RECT 11.0000 64.8000 11.4000 65.2000 ;
	    RECT 7.5000 61.1000 7.9000 64.8000 ;
	    RECT 10.2000 63.8000 10.6000 64.6000 ;
	    RECT 11.0000 64.1000 11.3000 64.8000 ;
	    RECT 12.6000 64.1000 12.9000 65.8000 ;
	    RECT 14.2000 65.2000 14.5000 66.8000 ;
	    RECT 15.1000 66.9000 16.0000 67.1000 ;
	    RECT 20.0000 67.1000 20.4000 69.9000 ;
	    RECT 21.7000 68.2000 22.1000 69.9000 ;
	    RECT 21.4000 67.8000 22.6000 68.2000 ;
	    RECT 21.4000 67.2000 21.7000 67.8000 ;
	    RECT 20.0000 66.9000 20.9000 67.1000 ;
	    RECT 15.1000 66.8000 15.9000 66.9000 ;
	    RECT 20.1000 66.8000 20.9000 66.9000 ;
	    RECT 21.4000 66.8000 21.8000 67.2000 ;
	    RECT 15.1000 65.2000 15.4000 66.8000 ;
	    RECT 16.2000 65.8000 17.0000 66.2000 ;
	    RECT 19.0000 65.8000 20.2000 66.2000 ;
	    RECT 14.2000 64.8000 14.6000 65.2000 ;
	    RECT 15.0000 64.8000 15.4000 65.2000 ;
	    RECT 17.4000 64.8000 17.8000 65.6000 ;
	    RECT 20.6000 65.2000 20.9000 66.8000 ;
	    RECT 20.6000 64.8000 21.0000 65.2000 ;
	    RECT 11.0000 63.8000 12.9000 64.1000 ;
	    RECT 13.4000 63.8000 13.8000 64.6000 ;
	    RECT 11.0000 63.5000 11.3000 63.8000 ;
	    RECT 14.2000 63.5000 14.5000 64.8000 ;
	    RECT 9.5000 63.2000 11.3000 63.5000 ;
	    RECT 9.5000 63.1000 9.8000 63.2000 ;
	    RECT 9.4000 61.1000 9.8000 63.1000 ;
	    RECT 11.0000 63.1000 11.3000 63.2000 ;
	    RECT 12.7000 63.2000 14.5000 63.5000 ;
	    RECT 12.7000 63.1000 13.0000 63.2000 ;
	    RECT 11.0000 61.1000 11.4000 63.1000 ;
	    RECT 12.6000 61.1000 13.0000 63.1000 ;
	    RECT 14.2000 63.1000 14.5000 63.2000 ;
	    RECT 15.1000 63.5000 15.4000 64.8000 ;
	    RECT 15.8000 63.8000 16.2000 64.6000 ;
	    RECT 19.0000 64.1000 19.4000 64.2000 ;
	    RECT 19.8000 64.1000 20.2000 64.6000 ;
	    RECT 19.0000 63.8000 20.2000 64.1000 ;
	    RECT 20.6000 63.5000 20.9000 64.8000 ;
	    RECT 15.1000 63.2000 16.9000 63.5000 ;
	    RECT 15.1000 63.1000 15.4000 63.2000 ;
	    RECT 14.2000 61.1000 14.6000 63.1000 ;
	    RECT 15.0000 61.1000 15.4000 63.1000 ;
	    RECT 16.6000 63.1000 16.9000 63.2000 ;
	    RECT 19.1000 63.2000 20.9000 63.5000 ;
	    RECT 19.1000 63.1000 19.4000 63.2000 ;
	    RECT 16.6000 61.1000 17.0000 63.1000 ;
	    RECT 19.0000 61.1000 19.4000 63.1000 ;
	    RECT 20.6000 63.1000 20.9000 63.2000 ;
	    RECT 20.6000 61.1000 21.0000 63.1000 ;
	    RECT 22.2000 61.1000 22.6000 67.8000 ;
	    RECT 23.0000 66.8000 23.4000 67.6000 ;
	    RECT 24.4000 67.1000 24.8000 69.9000 ;
	    RECT 27.8000 68.9000 28.2000 69.9000 ;
	    RECT 27.0000 67.8000 27.4000 68.6000 ;
	    RECT 27.9000 67.8000 28.2000 68.9000 ;
	    RECT 29.4000 67.9000 29.8000 69.9000 ;
	    RECT 27.9000 67.5000 29.1000 67.8000 ;
	    RECT 23.9000 66.9000 24.8000 67.1000 ;
	    RECT 23.9000 66.8000 24.7000 66.9000 ;
	    RECT 23.9000 65.2000 24.2000 66.8000 ;
	    RECT 25.0000 65.8000 25.8000 66.2000 ;
	    RECT 28.8000 66.0000 29.1000 67.5000 ;
	    RECT 29.5000 66.2000 29.8000 67.9000 ;
	    RECT 32.0000 67.1000 32.4000 69.9000 ;
	    RECT 34.7000 68.2000 35.1000 69.9000 ;
	    RECT 34.2000 67.9000 35.1000 68.2000 ;
	    RECT 32.0000 66.9000 32.9000 67.1000 ;
	    RECT 32.1000 66.8000 32.9000 66.9000 ;
	    RECT 33.4000 66.8000 33.8000 67.6000 ;
	    RECT 28.7000 65.7000 29.1000 66.0000 ;
	    RECT 29.4000 65.8000 29.8000 66.2000 ;
	    RECT 31.0000 65.8000 31.8000 66.2000 ;
	    RECT 27.0000 65.6000 29.1000 65.7000 ;
	    RECT 23.8000 64.8000 24.2000 65.2000 ;
	    RECT 23.9000 63.5000 24.2000 64.8000 ;
	    RECT 24.6000 63.8000 25.0000 65.2000 ;
	    RECT 25.4000 65.1000 25.8000 65.2000 ;
	    RECT 26.2000 65.1000 26.6000 65.6000 ;
	    RECT 25.4000 64.8000 26.6000 65.1000 ;
	    RECT 27.0000 65.4000 29.0000 65.6000 ;
	    RECT 23.9000 63.2000 25.7000 63.5000 ;
	    RECT 23.9000 63.1000 24.2000 63.2000 ;
	    RECT 23.8000 61.1000 24.2000 63.1000 ;
	    RECT 25.4000 63.1000 25.7000 63.2000 ;
	    RECT 25.4000 61.1000 25.8000 63.1000 ;
	    RECT 27.0000 61.1000 27.4000 65.4000 ;
	    RECT 29.5000 65.1000 29.8000 65.8000 ;
	    RECT 29.1000 64.8000 29.8000 65.1000 ;
	    RECT 30.2000 64.8000 30.6000 65.6000 ;
	    RECT 32.6000 65.2000 32.9000 66.8000 ;
	    RECT 32.6000 64.8000 33.0000 65.2000 ;
	    RECT 29.1000 61.1000 29.5000 64.8000 ;
	    RECT 31.0000 63.8000 31.4000 64.2000 ;
	    RECT 31.8000 63.8000 32.2000 64.6000 ;
	    RECT 31.0000 63.5000 31.3000 63.8000 ;
	    RECT 32.6000 63.5000 32.9000 64.8000 ;
	    RECT 31.0000 63.2000 32.9000 63.5000 ;
	    RECT 31.0000 61.1000 31.4000 63.2000 ;
	    RECT 32.6000 63.1000 32.9000 63.2000 ;
	    RECT 32.6000 61.1000 33.0000 63.1000 ;
	    RECT 34.2000 61.1000 34.6000 67.9000 ;
	    RECT 35.0000 65.1000 35.4000 65.2000 ;
	    RECT 35.8000 65.1000 36.2000 69.9000 ;
	    RECT 38.7000 69.2000 39.1000 69.9000 ;
	    RECT 38.7000 68.8000 39.4000 69.2000 ;
	    RECT 38.7000 68.2000 39.1000 68.8000 ;
	    RECT 38.2000 67.9000 39.1000 68.2000 ;
	    RECT 40.1000 68.2000 40.5000 69.9000 ;
	    RECT 40.1000 67.9000 41.0000 68.2000 ;
	    RECT 37.4000 66.8000 37.8000 67.6000 ;
	    RECT 35.0000 64.8000 36.2000 65.1000 ;
	    RECT 35.0000 64.4000 35.4000 64.8000 ;
	    RECT 35.8000 61.1000 36.2000 64.8000 ;
	    RECT 38.2000 61.1000 38.6000 67.9000 ;
	    RECT 40.6000 64.1000 41.0000 67.9000 ;
	    RECT 41.4000 66.8000 41.8000 67.6000 ;
	    RECT 43.0000 67.1000 43.4000 69.9000 ;
	    RECT 43.8000 68.0000 44.2000 69.9000 ;
	    RECT 45.4000 68.0000 45.8000 69.9000 ;
	    RECT 43.8000 67.9000 45.8000 68.0000 ;
	    RECT 46.2000 67.9000 46.6000 69.9000 ;
	    RECT 47.3000 68.2000 47.7000 69.9000 ;
	    RECT 47.3000 67.9000 48.2000 68.2000 ;
	    RECT 43.9000 67.7000 45.7000 67.9000 ;
	    RECT 44.2000 67.2000 44.6000 67.4000 ;
	    RECT 46.2000 67.2000 46.5000 67.9000 ;
	    RECT 43.8000 67.1000 44.6000 67.2000 ;
	    RECT 43.0000 66.9000 44.6000 67.1000 ;
	    RECT 43.0000 66.8000 44.2000 66.9000 ;
	    RECT 45.3000 66.8000 46.6000 67.2000 ;
	    RECT 41.4000 64.1000 41.8000 64.2000 ;
	    RECT 40.6000 63.8000 41.8000 64.1000 ;
	    RECT 40.6000 61.1000 41.0000 63.8000 ;
	    RECT 43.0000 61.1000 43.4000 66.8000 ;
	    RECT 44.6000 65.8000 45.0000 66.6000 ;
	    RECT 45.3000 65.1000 45.6000 66.8000 ;
	    RECT 46.2000 65.1000 46.6000 65.2000 ;
	    RECT 45.1000 64.8000 45.6000 65.1000 ;
	    RECT 45.9000 64.8000 46.6000 65.1000 ;
	    RECT 47.8000 65.1000 48.2000 67.9000 ;
	    RECT 48.6000 66.8000 49.0000 67.6000 ;
	    RECT 49.4000 67.1000 49.8000 67.2000 ;
	    RECT 50.2000 67.1000 50.6000 69.9000 ;
	    RECT 51.0000 67.9000 51.4000 69.9000 ;
	    RECT 51.8000 68.0000 52.2000 69.9000 ;
	    RECT 53.4000 68.0000 53.8000 69.9000 ;
	    RECT 51.8000 67.9000 53.8000 68.0000 ;
	    RECT 51.1000 67.2000 51.4000 67.9000 ;
	    RECT 51.9000 67.7000 53.7000 67.9000 ;
	    RECT 53.0000 67.2000 53.4000 67.4000 ;
	    RECT 49.4000 66.8000 50.6000 67.1000 ;
	    RECT 51.0000 66.8000 52.3000 67.2000 ;
	    RECT 53.0000 66.9000 53.8000 67.2000 ;
	    RECT 53.4000 66.8000 53.8000 66.9000 ;
	    RECT 48.6000 65.1000 49.0000 65.2000 ;
	    RECT 47.8000 64.8000 49.0000 65.1000 ;
	    RECT 45.1000 61.1000 45.5000 64.8000 ;
	    RECT 45.9000 64.2000 46.2000 64.8000 ;
	    RECT 45.8000 63.8000 46.2000 64.2000 ;
	    RECT 47.8000 61.1000 48.2000 64.8000 ;
	    RECT 50.2000 61.1000 50.6000 66.8000 ;
	    RECT 52.0000 65.2000 52.3000 66.8000 ;
	    RECT 52.6000 65.8000 53.0000 66.6000 ;
	    RECT 51.0000 65.1000 51.4000 65.2000 ;
	    RECT 51.0000 64.8000 51.7000 65.1000 ;
	    RECT 52.0000 64.8000 53.0000 65.2000 ;
	    RECT 51.4000 64.2000 51.7000 64.8000 ;
	    RECT 51.4000 63.8000 51.8000 64.2000 ;
	    RECT 52.1000 61.1000 52.5000 64.8000 ;
	    RECT 54.2000 64.1000 54.6000 64.2000 ;
	    RECT 55.0000 64.1000 55.4000 69.9000 ;
	    RECT 57.1000 69.2000 57.5000 69.9000 ;
	    RECT 58.5000 69.2000 58.9000 69.9000 ;
	    RECT 57.1000 68.8000 57.8000 69.2000 ;
	    RECT 58.5000 68.8000 59.4000 69.2000 ;
	    RECT 57.1000 68.2000 57.5000 68.8000 ;
	    RECT 56.6000 67.9000 57.5000 68.2000 ;
	    RECT 58.5000 68.2000 58.9000 68.8000 ;
	    RECT 58.5000 67.9000 59.4000 68.2000 ;
	    RECT 55.8000 66.8000 56.2000 67.6000 ;
	    RECT 54.2000 63.8000 55.4000 64.1000 ;
	    RECT 55.0000 61.1000 55.4000 63.8000 ;
	    RECT 56.6000 61.1000 57.0000 67.9000 ;
	    RECT 57.4000 64.4000 57.8000 65.2000 ;
	    RECT 58.2000 64.4000 58.6000 65.2000 ;
	    RECT 59.0000 61.1000 59.4000 67.9000 ;
	    RECT 63.0000 65.1000 63.4000 69.9000 ;
	    RECT 64.1000 69.2000 64.5000 69.9000 ;
	    RECT 67.5000 69.2000 67.9000 69.9000 ;
	    RECT 64.1000 68.8000 65.0000 69.2000 ;
	    RECT 67.5000 68.8000 68.2000 69.2000 ;
	    RECT 64.1000 68.2000 64.5000 68.8000 ;
	    RECT 67.5000 68.2000 67.9000 68.8000 ;
	    RECT 64.1000 67.9000 65.0000 68.2000 ;
	    RECT 63.8000 65.1000 64.2000 65.2000 ;
	    RECT 63.0000 64.8000 64.2000 65.1000 ;
	    RECT 63.0000 61.1000 63.4000 64.8000 ;
	    RECT 63.8000 64.4000 64.2000 64.8000 ;
	    RECT 64.6000 61.1000 65.0000 67.9000 ;
	    RECT 67.0000 67.9000 67.9000 68.2000 ;
	    RECT 65.4000 67.1000 65.8000 67.6000 ;
	    RECT 66.2000 67.1000 66.6000 67.6000 ;
	    RECT 65.4000 66.8000 66.6000 67.1000 ;
	    RECT 67.0000 61.1000 67.4000 67.9000 ;
	    RECT 67.8000 65.1000 68.2000 65.2000 ;
	    RECT 68.6000 65.1000 69.0000 69.9000 ;
	    RECT 67.8000 64.8000 69.0000 65.1000 ;
	    RECT 70.2000 67.9000 70.6000 69.9000 ;
	    RECT 71.8000 68.9000 72.2000 69.9000 ;
	    RECT 70.2000 66.2000 70.5000 67.9000 ;
	    RECT 71.8000 67.8000 72.1000 68.9000 ;
	    RECT 72.6000 67.8000 73.0000 68.6000 ;
	    RECT 70.9000 67.5000 72.1000 67.8000 ;
	    RECT 70.2000 65.8000 70.6000 66.2000 ;
	    RECT 70.9000 66.0000 71.2000 67.5000 ;
	    RECT 70.2000 65.1000 70.5000 65.8000 ;
	    RECT 70.9000 65.7000 71.3000 66.0000 ;
	    RECT 70.9000 65.6000 73.0000 65.7000 ;
	    RECT 71.0000 65.4000 73.0000 65.6000 ;
	    RECT 70.2000 64.8000 70.9000 65.1000 ;
	    RECT 67.8000 64.4000 68.2000 64.8000 ;
	    RECT 68.6000 61.1000 69.0000 64.8000 ;
	    RECT 70.5000 61.1000 70.9000 64.8000 ;
	    RECT 72.6000 61.1000 73.0000 65.4000 ;
	    RECT 74.2000 65.1000 74.6000 69.9000 ;
	    RECT 75.3000 69.2000 75.7000 69.9000 ;
	    RECT 75.3000 68.8000 76.2000 69.2000 ;
	    RECT 75.3000 68.2000 75.7000 68.8000 ;
	    RECT 75.3000 67.9000 76.2000 68.2000 ;
	    RECT 77.4000 67.9000 77.8000 69.9000 ;
	    RECT 79.5000 69.2000 79.9000 69.9000 ;
	    RECT 79.5000 68.8000 80.2000 69.2000 ;
	    RECT 79.5000 68.4000 79.9000 68.8000 ;
	    RECT 79.5000 67.9000 80.2000 68.4000 ;
	    RECT 80.6000 67.9000 81.0000 69.9000 ;
	    RECT 82.7000 69.2000 83.1000 69.9000 ;
	    RECT 82.7000 68.8000 83.4000 69.2000 ;
	    RECT 82.7000 68.4000 83.1000 68.8000 ;
	    RECT 82.7000 67.9000 83.4000 68.4000 ;
	    RECT 75.0000 65.1000 75.4000 65.2000 ;
	    RECT 74.2000 64.8000 75.4000 65.1000 ;
	    RECT 74.2000 61.1000 74.6000 64.8000 ;
	    RECT 75.0000 64.4000 75.4000 64.8000 ;
	    RECT 75.8000 61.1000 76.2000 67.9000 ;
	    RECT 77.5000 67.8000 77.8000 67.9000 ;
	    RECT 77.5000 67.6000 78.4000 67.8000 ;
	    RECT 76.6000 66.8000 77.0000 67.6000 ;
	    RECT 77.5000 67.5000 79.6000 67.6000 ;
	    RECT 78.1000 67.3000 79.6000 67.5000 ;
	    RECT 79.2000 67.2000 79.6000 67.3000 ;
	    RECT 77.4000 66.4000 77.8000 67.2000 ;
	    RECT 78.4000 66.9000 78.8000 67.0000 ;
	    RECT 78.3000 66.6000 78.8000 66.9000 ;
	    RECT 78.3000 66.2000 78.6000 66.6000 ;
	    RECT 78.2000 65.8000 78.6000 66.2000 ;
	    RECT 79.2000 65.5000 79.5000 67.2000 ;
	    RECT 79.9000 66.2000 80.2000 67.9000 ;
	    RECT 80.7000 67.8000 81.0000 67.9000 ;
	    RECT 80.7000 67.6000 81.6000 67.8000 ;
	    RECT 80.7000 67.5000 82.8000 67.6000 ;
	    RECT 81.3000 67.3000 82.8000 67.5000 ;
	    RECT 82.4000 67.2000 82.8000 67.3000 ;
	    RECT 80.6000 66.4000 81.0000 67.2000 ;
	    RECT 81.6000 66.9000 82.0000 67.0000 ;
	    RECT 81.5000 66.6000 82.0000 66.9000 ;
	    RECT 81.5000 66.2000 81.8000 66.6000 ;
	    RECT 79.8000 65.8000 80.2000 66.2000 ;
	    RECT 81.4000 65.8000 81.8000 66.2000 ;
	    RECT 78.3000 65.2000 79.5000 65.5000 ;
	    RECT 78.3000 63.1000 78.6000 65.2000 ;
	    RECT 79.9000 65.1000 80.2000 65.8000 ;
	    RECT 82.4000 65.5000 82.7000 67.2000 ;
	    RECT 83.1000 66.2000 83.4000 67.9000 ;
	    RECT 83.8000 67.5000 84.2000 69.9000 ;
	    RECT 86.0000 69.2000 86.4000 69.9000 ;
	    RECT 85.4000 68.9000 86.4000 69.2000 ;
	    RECT 88.2000 68.9000 88.6000 69.9000 ;
	    RECT 90.3000 69.2000 90.9000 69.9000 ;
	    RECT 90.2000 68.9000 90.9000 69.2000 ;
	    RECT 85.4000 68.5000 85.8000 68.9000 ;
	    RECT 88.2000 68.6000 88.5000 68.9000 ;
	    RECT 86.2000 68.2000 86.6000 68.6000 ;
	    RECT 87.1000 68.3000 88.5000 68.6000 ;
	    RECT 90.2000 68.5000 90.6000 68.9000 ;
	    RECT 87.1000 68.2000 87.5000 68.3000 ;
	    RECT 84.2000 67.1000 85.0000 67.2000 ;
	    RECT 86.3000 67.1000 86.6000 68.2000 ;
	    RECT 91.0000 67.8000 91.4000 68.2000 ;
	    RECT 91.0000 67.7000 91.5000 67.8000 ;
	    RECT 92.6000 67.7000 93.0000 69.9000 ;
	    RECT 91.0000 67.4000 93.0000 67.7000 ;
	    RECT 89.1000 67.1000 89.5000 67.2000 ;
	    RECT 84.2000 66.8000 89.7000 67.1000 ;
	    RECT 85.7000 66.7000 86.1000 66.8000 ;
	    RECT 83.0000 65.8000 83.4000 66.2000 ;
	    RECT 84.9000 66.2000 85.3000 66.3000 ;
	    RECT 86.2000 66.2000 86.6000 66.3000 ;
	    RECT 84.9000 65.9000 87.4000 66.2000 ;
	    RECT 87.0000 65.8000 87.4000 65.9000 ;
	    RECT 88.6000 66.1000 89.0000 66.2000 ;
	    RECT 89.4000 66.1000 89.7000 66.8000 ;
	    RECT 90.2000 66.4000 90.6000 66.5000 ;
	    RECT 90.2000 66.1000 92.1000 66.4000 ;
	    RECT 88.6000 65.8000 89.7000 66.1000 ;
	    RECT 91.7000 66.0000 92.1000 66.1000 ;
	    RECT 78.2000 61.1000 78.6000 63.1000 ;
	    RECT 79.8000 61.1000 80.2000 65.1000 ;
	    RECT 81.5000 65.2000 82.7000 65.5000 ;
	    RECT 81.5000 63.1000 81.8000 65.2000 ;
	    RECT 83.1000 65.1000 83.4000 65.8000 ;
	    RECT 81.4000 61.1000 81.8000 63.1000 ;
	    RECT 83.0000 61.1000 83.4000 65.1000 ;
	    RECT 83.8000 65.5000 86.6000 65.6000 ;
	    RECT 83.8000 65.4000 86.7000 65.5000 ;
	    RECT 83.8000 65.3000 88.7000 65.4000 ;
	    RECT 83.8000 61.1000 84.2000 65.3000 ;
	    RECT 86.3000 65.1000 88.7000 65.3000 ;
	    RECT 85.4000 64.5000 88.1000 64.8000 ;
	    RECT 85.4000 64.4000 85.8000 64.5000 ;
	    RECT 87.7000 64.4000 88.1000 64.5000 ;
	    RECT 88.4000 64.5000 88.7000 65.1000 ;
	    RECT 89.4000 65.2000 89.7000 65.8000 ;
	    RECT 90.9000 65.7000 91.3000 65.8000 ;
	    RECT 92.6000 65.7000 93.0000 67.4000 ;
	    RECT 95.0000 67.9000 95.4000 69.9000 ;
	    RECT 95.7000 68.2000 96.1000 68.6000 ;
	    RECT 94.2000 66.4000 94.6000 67.2000 ;
	    RECT 93.4000 66.1000 93.8000 66.2000 ;
	    RECT 95.0000 66.1000 95.3000 67.9000 ;
	    RECT 95.8000 67.8000 96.2000 68.2000 ;
	    RECT 96.6000 66.8000 97.0000 67.6000 ;
	    RECT 95.8000 66.1000 96.2000 66.2000 ;
	    RECT 93.4000 65.8000 94.2000 66.1000 ;
	    RECT 95.0000 65.8000 96.2000 66.1000 ;
	    RECT 90.9000 65.4000 93.0000 65.7000 ;
	    RECT 93.8000 65.6000 94.2000 65.8000 ;
	    RECT 89.4000 64.9000 90.6000 65.2000 ;
	    RECT 89.1000 64.5000 89.5000 64.6000 ;
	    RECT 88.4000 64.2000 89.5000 64.5000 ;
	    RECT 90.3000 64.4000 90.6000 64.9000 ;
	    RECT 90.3000 64.0000 91.0000 64.4000 ;
	    RECT 87.1000 63.7000 87.5000 63.8000 ;
	    RECT 88.5000 63.7000 88.9000 63.8000 ;
	    RECT 85.4000 63.1000 85.8000 63.5000 ;
	    RECT 87.1000 63.4000 88.9000 63.7000 ;
	    RECT 88.2000 63.1000 88.5000 63.4000 ;
	    RECT 90.2000 63.1000 90.6000 63.5000 ;
	    RECT 85.4000 62.8000 86.4000 63.1000 ;
	    RECT 86.0000 61.1000 86.4000 62.8000 ;
	    RECT 88.2000 61.1000 88.6000 63.1000 ;
	    RECT 90.3000 61.1000 90.9000 63.1000 ;
	    RECT 92.6000 61.1000 93.0000 65.4000 ;
	    RECT 95.8000 65.2000 96.1000 65.8000 ;
	    RECT 93.4000 64.8000 95.4000 65.1000 ;
	    RECT 93.4000 61.1000 93.8000 64.8000 ;
	    RECT 95.0000 61.1000 95.4000 64.8000 ;
	    RECT 95.8000 61.1000 96.2000 65.2000 ;
	    RECT 97.4000 61.1000 97.8000 69.9000 ;
	    RECT 98.2000 67.9000 98.6000 69.9000 ;
	    RECT 100.3000 68.4000 100.7000 69.9000 ;
	    RECT 100.3000 67.9000 101.0000 68.4000 ;
	    RECT 98.3000 67.8000 98.6000 67.9000 ;
	    RECT 98.3000 67.6000 99.2000 67.8000 ;
	    RECT 98.3000 67.5000 100.4000 67.6000 ;
	    RECT 98.9000 67.3000 100.4000 67.5000 ;
	    RECT 100.0000 67.2000 100.4000 67.3000 ;
	    RECT 98.2000 66.4000 98.6000 67.2000 ;
	    RECT 99.2000 66.9000 99.6000 67.0000 ;
	    RECT 99.1000 66.6000 99.6000 66.9000 ;
	    RECT 99.1000 66.2000 99.4000 66.6000 ;
	    RECT 99.0000 65.8000 99.4000 66.2000 ;
	    RECT 100.0000 65.5000 100.3000 67.2000 ;
	    RECT 100.7000 66.2000 101.0000 67.9000 ;
	    RECT 101.4000 67.5000 101.8000 69.9000 ;
	    RECT 103.6000 69.2000 104.0000 69.9000 ;
	    RECT 103.0000 68.9000 104.0000 69.2000 ;
	    RECT 105.8000 68.9000 106.2000 69.9000 ;
	    RECT 107.9000 69.2000 108.5000 69.9000 ;
	    RECT 107.8000 68.9000 108.5000 69.2000 ;
	    RECT 110.2000 69.1000 110.6000 69.9000 ;
	    RECT 111.0000 69.1000 111.4000 69.2000 ;
	    RECT 103.0000 68.5000 103.4000 68.9000 ;
	    RECT 105.8000 68.6000 106.1000 68.9000 ;
	    RECT 103.8000 68.2000 104.2000 68.6000 ;
	    RECT 104.7000 68.3000 106.1000 68.6000 ;
	    RECT 107.8000 68.5000 108.2000 68.9000 ;
	    RECT 110.2000 68.8000 111.4000 69.1000 ;
	    RECT 104.7000 68.2000 105.1000 68.3000 ;
	    RECT 101.8000 67.1000 102.6000 67.2000 ;
	    RECT 103.9000 67.1000 104.2000 68.2000 ;
	    RECT 108.7000 67.7000 109.1000 67.8000 ;
	    RECT 110.2000 67.7000 110.6000 68.8000 ;
	    RECT 108.7000 67.4000 110.6000 67.7000 ;
	    RECT 106.7000 67.1000 107.1000 67.2000 ;
	    RECT 101.8000 66.8000 107.3000 67.1000 ;
	    RECT 103.3000 66.7000 103.7000 66.8000 ;
	    RECT 100.6000 65.8000 101.0000 66.2000 ;
	    RECT 102.5000 66.2000 102.9000 66.3000 ;
	    RECT 103.8000 66.2000 104.2000 66.3000 ;
	    RECT 102.5000 65.9000 105.0000 66.2000 ;
	    RECT 104.6000 65.8000 105.0000 65.9000 ;
	    RECT 99.1000 65.2000 100.3000 65.5000 ;
	    RECT 99.1000 63.1000 99.4000 65.2000 ;
	    RECT 100.7000 65.1000 101.0000 65.8000 ;
	    RECT 99.0000 61.1000 99.4000 63.1000 ;
	    RECT 100.6000 61.1000 101.0000 65.1000 ;
	    RECT 101.4000 65.5000 104.2000 65.6000 ;
	    RECT 101.4000 65.4000 104.3000 65.5000 ;
	    RECT 101.4000 65.3000 106.3000 65.4000 ;
	    RECT 101.4000 61.1000 101.8000 65.3000 ;
	    RECT 103.9000 65.1000 106.3000 65.3000 ;
	    RECT 103.0000 64.5000 105.7000 64.8000 ;
	    RECT 103.0000 64.4000 103.4000 64.5000 ;
	    RECT 105.3000 64.4000 105.7000 64.5000 ;
	    RECT 106.0000 64.5000 106.3000 65.1000 ;
	    RECT 107.0000 65.2000 107.3000 66.8000 ;
	    RECT 107.8000 66.4000 108.2000 66.5000 ;
	    RECT 107.8000 66.1000 109.7000 66.4000 ;
	    RECT 109.3000 66.0000 109.7000 66.1000 ;
	    RECT 108.5000 65.7000 108.9000 65.8000 ;
	    RECT 110.2000 65.7000 110.6000 67.4000 ;
	    RECT 113.4000 67.6000 113.8000 69.9000 ;
	    RECT 115.0000 67.6000 115.4000 69.9000 ;
	    RECT 116.6000 67.6000 117.0000 69.9000 ;
	    RECT 118.2000 67.6000 118.6000 69.9000 ;
	    RECT 113.4000 67.2000 114.3000 67.6000 ;
	    RECT 115.0000 67.2000 116.1000 67.6000 ;
	    RECT 116.6000 67.2000 117.7000 67.6000 ;
	    RECT 118.2000 67.2000 119.4000 67.6000 ;
	    RECT 119.8000 67.5000 120.2000 69.9000 ;
	    RECT 122.0000 69.2000 122.4000 69.9000 ;
	    RECT 121.4000 68.9000 122.4000 69.2000 ;
	    RECT 124.2000 68.9000 124.6000 69.9000 ;
	    RECT 126.3000 69.2000 126.9000 69.9000 ;
	    RECT 126.2000 68.9000 126.9000 69.2000 ;
	    RECT 121.4000 68.5000 121.8000 68.9000 ;
	    RECT 124.2000 68.6000 124.5000 68.9000 ;
	    RECT 122.2000 68.2000 122.6000 68.6000 ;
	    RECT 123.1000 68.3000 124.5000 68.6000 ;
	    RECT 126.2000 68.5000 126.6000 68.9000 ;
	    RECT 123.1000 68.2000 123.5000 68.3000 ;
	    RECT 113.9000 66.9000 114.3000 67.2000 ;
	    RECT 115.7000 66.9000 116.1000 67.2000 ;
	    RECT 117.3000 66.9000 117.7000 67.2000 ;
	    RECT 113.9000 66.5000 115.2000 66.9000 ;
	    RECT 115.7000 66.5000 116.9000 66.9000 ;
	    RECT 117.3000 66.5000 118.6000 66.9000 ;
	    RECT 113.9000 65.8000 114.3000 66.5000 ;
	    RECT 115.7000 65.8000 116.1000 66.5000 ;
	    RECT 117.3000 65.8000 117.7000 66.5000 ;
	    RECT 119.0000 65.8000 119.4000 67.2000 ;
	    RECT 120.2000 67.1000 121.0000 67.2000 ;
	    RECT 122.3000 67.1000 122.6000 68.2000 ;
	    RECT 127.1000 67.7000 127.5000 67.8000 ;
	    RECT 128.6000 67.7000 129.0000 69.9000 ;
	    RECT 129.7000 69.2000 130.1000 69.9000 ;
	    RECT 129.4000 68.8000 130.1000 69.2000 ;
	    RECT 129.7000 68.4000 130.1000 68.8000 ;
	    RECT 127.1000 67.4000 129.0000 67.7000 ;
	    RECT 125.1000 67.1000 125.5000 67.2000 ;
	    RECT 120.2000 66.8000 125.7000 67.1000 ;
	    RECT 121.7000 66.7000 122.1000 66.8000 ;
	    RECT 120.9000 66.2000 121.3000 66.3000 ;
	    RECT 122.2000 66.2000 122.6000 66.3000 ;
	    RECT 120.9000 65.9000 123.4000 66.2000 ;
	    RECT 123.0000 65.8000 123.4000 65.9000 ;
	    RECT 108.5000 65.4000 110.6000 65.7000 ;
	    RECT 107.0000 64.9000 108.2000 65.2000 ;
	    RECT 106.7000 64.5000 107.1000 64.6000 ;
	    RECT 106.0000 64.2000 107.1000 64.5000 ;
	    RECT 107.9000 64.4000 108.2000 64.9000 ;
	    RECT 107.9000 64.0000 108.6000 64.4000 ;
	    RECT 104.7000 63.7000 105.1000 63.8000 ;
	    RECT 106.1000 63.7000 106.5000 63.8000 ;
	    RECT 103.0000 63.1000 103.4000 63.5000 ;
	    RECT 104.7000 63.4000 106.5000 63.7000 ;
	    RECT 105.8000 63.1000 106.1000 63.4000 ;
	    RECT 107.8000 63.1000 108.2000 63.5000 ;
	    RECT 103.0000 62.8000 104.0000 63.1000 ;
	    RECT 103.6000 61.1000 104.0000 62.8000 ;
	    RECT 105.8000 61.1000 106.2000 63.1000 ;
	    RECT 107.9000 61.1000 108.5000 63.1000 ;
	    RECT 110.2000 61.1000 110.6000 65.4000 ;
	    RECT 113.4000 65.4000 114.3000 65.8000 ;
	    RECT 115.0000 65.4000 116.1000 65.8000 ;
	    RECT 116.6000 65.4000 117.7000 65.8000 ;
	    RECT 118.2000 65.4000 119.4000 65.8000 ;
	    RECT 119.8000 65.5000 122.6000 65.6000 ;
	    RECT 119.8000 65.4000 122.7000 65.5000 ;
	    RECT 113.4000 61.1000 113.8000 65.4000 ;
	    RECT 115.0000 61.1000 115.4000 65.4000 ;
	    RECT 116.6000 61.1000 117.0000 65.4000 ;
	    RECT 118.2000 61.1000 118.6000 65.4000 ;
	    RECT 119.8000 65.3000 124.7000 65.4000 ;
	    RECT 119.8000 61.1000 120.2000 65.3000 ;
	    RECT 122.3000 65.1000 124.7000 65.3000 ;
	    RECT 121.4000 64.5000 124.1000 64.8000 ;
	    RECT 121.4000 64.4000 121.8000 64.5000 ;
	    RECT 123.7000 64.4000 124.1000 64.5000 ;
	    RECT 124.4000 64.5000 124.7000 65.1000 ;
	    RECT 125.4000 65.2000 125.7000 66.8000 ;
	    RECT 126.2000 66.4000 126.6000 66.5000 ;
	    RECT 126.2000 66.1000 128.1000 66.4000 ;
	    RECT 127.7000 66.0000 128.1000 66.1000 ;
	    RECT 126.9000 65.7000 127.3000 65.8000 ;
	    RECT 128.6000 65.7000 129.0000 67.4000 ;
	    RECT 126.9000 65.4000 129.0000 65.7000 ;
	    RECT 125.4000 64.9000 126.6000 65.2000 ;
	    RECT 125.1000 64.5000 125.5000 64.6000 ;
	    RECT 124.4000 64.2000 125.5000 64.5000 ;
	    RECT 126.3000 64.4000 126.6000 64.9000 ;
	    RECT 126.3000 64.0000 127.0000 64.4000 ;
	    RECT 123.1000 63.7000 123.5000 63.8000 ;
	    RECT 124.5000 63.7000 124.9000 63.8000 ;
	    RECT 121.4000 63.1000 121.8000 63.5000 ;
	    RECT 123.1000 63.4000 124.9000 63.7000 ;
	    RECT 124.2000 63.1000 124.5000 63.4000 ;
	    RECT 126.2000 63.1000 126.6000 63.5000 ;
	    RECT 121.4000 62.8000 122.4000 63.1000 ;
	    RECT 122.0000 61.1000 122.4000 62.8000 ;
	    RECT 124.2000 61.1000 124.6000 63.1000 ;
	    RECT 126.3000 61.1000 126.9000 63.1000 ;
	    RECT 128.6000 61.1000 129.0000 65.4000 ;
	    RECT 129.4000 67.9000 130.1000 68.4000 ;
	    RECT 131.8000 67.9000 132.2000 69.9000 ;
	    RECT 129.4000 66.2000 129.7000 67.9000 ;
	    RECT 131.8000 67.8000 132.1000 67.9000 ;
	    RECT 131.2000 67.6000 132.1000 67.8000 ;
	    RECT 130.0000 67.5000 132.1000 67.6000 ;
	    RECT 132.6000 67.5000 133.0000 69.9000 ;
	    RECT 134.8000 69.2000 135.2000 69.9000 ;
	    RECT 134.2000 68.9000 135.2000 69.2000 ;
	    RECT 137.0000 68.9000 137.4000 69.9000 ;
	    RECT 139.1000 69.2000 139.7000 69.9000 ;
	    RECT 139.0000 68.9000 139.7000 69.2000 ;
	    RECT 134.2000 68.5000 134.6000 68.9000 ;
	    RECT 137.0000 68.6000 137.3000 68.9000 ;
	    RECT 135.0000 68.2000 135.4000 68.6000 ;
	    RECT 135.9000 68.3000 137.3000 68.6000 ;
	    RECT 139.0000 68.5000 139.4000 68.9000 ;
	    RECT 135.9000 68.2000 136.3000 68.3000 ;
	    RECT 130.0000 67.3000 131.5000 67.5000 ;
	    RECT 130.0000 67.2000 130.4000 67.3000 ;
	    RECT 129.4000 65.8000 129.8000 66.2000 ;
	    RECT 129.4000 65.1000 129.7000 65.8000 ;
	    RECT 130.1000 65.5000 130.4000 67.2000 ;
	    RECT 130.8000 66.9000 131.2000 67.0000 ;
	    RECT 130.8000 66.6000 131.3000 66.9000 ;
	    RECT 131.0000 66.2000 131.3000 66.6000 ;
	    RECT 131.8000 66.4000 132.2000 67.2000 ;
	    RECT 133.0000 67.1000 133.8000 67.2000 ;
	    RECT 135.1000 67.1000 135.4000 68.2000 ;
	    RECT 139.9000 67.7000 140.3000 67.8000 ;
	    RECT 141.4000 67.7000 141.8000 69.9000 ;
	    RECT 142.2000 67.9000 142.6000 69.9000 ;
	    RECT 144.3000 69.2000 144.7000 69.9000 ;
	    RECT 144.3000 68.8000 145.0000 69.2000 ;
	    RECT 144.3000 68.4000 144.7000 68.8000 ;
	    RECT 144.3000 67.9000 145.0000 68.4000 ;
	    RECT 139.9000 67.4000 141.8000 67.7000 ;
	    RECT 142.3000 67.8000 142.6000 67.9000 ;
	    RECT 142.3000 67.6000 143.2000 67.8000 ;
	    RECT 142.3000 67.5000 144.4000 67.6000 ;
	    RECT 137.9000 67.1000 138.3000 67.2000 ;
	    RECT 133.0000 66.8000 138.5000 67.1000 ;
	    RECT 134.5000 66.7000 134.9000 66.8000 ;
	    RECT 133.7000 66.2000 134.1000 66.3000 ;
	    RECT 131.0000 65.8000 131.4000 66.2000 ;
	    RECT 133.7000 65.9000 136.2000 66.2000 ;
	    RECT 135.8000 65.8000 136.2000 65.9000 ;
	    RECT 132.6000 65.5000 135.4000 65.6000 ;
	    RECT 130.1000 65.2000 131.3000 65.5000 ;
	    RECT 129.4000 61.1000 129.8000 65.1000 ;
	    RECT 131.0000 63.1000 131.3000 65.2000 ;
	    RECT 132.6000 65.4000 135.5000 65.5000 ;
	    RECT 132.6000 65.3000 137.5000 65.4000 ;
	    RECT 131.0000 61.1000 131.4000 63.1000 ;
	    RECT 132.6000 61.1000 133.0000 65.3000 ;
	    RECT 135.1000 65.1000 137.5000 65.3000 ;
	    RECT 134.2000 64.5000 136.9000 64.8000 ;
	    RECT 134.2000 64.4000 134.6000 64.5000 ;
	    RECT 136.5000 64.4000 136.9000 64.5000 ;
	    RECT 137.2000 64.5000 137.5000 65.1000 ;
	    RECT 138.2000 65.2000 138.5000 66.8000 ;
	    RECT 139.0000 66.4000 139.4000 66.5000 ;
	    RECT 139.0000 66.1000 140.9000 66.4000 ;
	    RECT 140.5000 66.0000 140.9000 66.1000 ;
	    RECT 139.7000 65.7000 140.1000 65.8000 ;
	    RECT 141.4000 65.7000 141.8000 67.4000 ;
	    RECT 142.9000 67.3000 144.4000 67.5000 ;
	    RECT 144.0000 67.2000 144.4000 67.3000 ;
	    RECT 142.2000 66.4000 142.6000 67.2000 ;
	    RECT 143.2000 66.9000 143.6000 67.0000 ;
	    RECT 143.1000 66.6000 143.6000 66.9000 ;
	    RECT 143.1000 66.2000 143.4000 66.6000 ;
	    RECT 143.0000 65.8000 143.4000 66.2000 ;
	    RECT 139.7000 65.4000 141.8000 65.7000 ;
	    RECT 144.0000 65.5000 144.3000 67.2000 ;
	    RECT 144.7000 66.2000 145.0000 67.9000 ;
	    RECT 144.6000 65.8000 145.0000 66.2000 ;
	    RECT 138.2000 64.9000 139.4000 65.2000 ;
	    RECT 137.9000 64.5000 138.3000 64.6000 ;
	    RECT 137.2000 64.2000 138.3000 64.5000 ;
	    RECT 139.1000 64.4000 139.4000 64.9000 ;
	    RECT 141.4000 65.1000 141.8000 65.4000 ;
	    RECT 143.1000 65.2000 144.3000 65.5000 ;
	    RECT 142.2000 65.1000 142.6000 65.2000 ;
	    RECT 141.4000 64.8000 142.6000 65.1000 ;
	    RECT 139.1000 64.0000 139.8000 64.4000 ;
	    RECT 135.9000 63.7000 136.3000 63.8000 ;
	    RECT 137.3000 63.7000 137.7000 63.8000 ;
	    RECT 134.2000 63.1000 134.6000 63.5000 ;
	    RECT 135.9000 63.4000 137.7000 63.7000 ;
	    RECT 137.0000 63.1000 137.3000 63.4000 ;
	    RECT 139.0000 63.1000 139.4000 63.5000 ;
	    RECT 134.2000 62.8000 135.2000 63.1000 ;
	    RECT 134.8000 61.1000 135.2000 62.8000 ;
	    RECT 137.0000 61.1000 137.4000 63.1000 ;
	    RECT 139.1000 61.1000 139.7000 63.1000 ;
	    RECT 141.4000 61.1000 141.8000 64.8000 ;
	    RECT 143.1000 63.1000 143.4000 65.2000 ;
	    RECT 144.7000 65.1000 145.0000 65.8000 ;
	    RECT 143.0000 61.1000 143.4000 63.1000 ;
	    RECT 144.6000 61.1000 145.0000 65.1000 ;
	    RECT 145.4000 67.7000 145.8000 69.9000 ;
	    RECT 147.5000 69.2000 148.1000 69.9000 ;
	    RECT 147.5000 68.9000 148.2000 69.2000 ;
	    RECT 149.8000 68.9000 150.2000 69.9000 ;
	    RECT 152.0000 69.2000 152.4000 69.9000 ;
	    RECT 152.0000 68.9000 153.0000 69.2000 ;
	    RECT 147.8000 68.5000 148.2000 68.9000 ;
	    RECT 149.9000 68.6000 150.2000 68.9000 ;
	    RECT 149.9000 68.3000 151.3000 68.6000 ;
	    RECT 150.9000 68.2000 151.3000 68.3000 ;
	    RECT 151.8000 68.2000 152.2000 68.6000 ;
	    RECT 152.6000 68.5000 153.0000 68.9000 ;
	    RECT 146.9000 67.7000 147.3000 67.8000 ;
	    RECT 145.4000 67.4000 147.4000 67.7000 ;
	    RECT 145.4000 65.7000 145.8000 67.4000 ;
	    RECT 147.0000 66.8000 147.4000 67.4000 ;
	    RECT 148.9000 67.1000 149.3000 67.2000 ;
	    RECT 151.8000 67.1000 152.1000 68.2000 ;
	    RECT 154.2000 67.5000 154.6000 69.9000 ;
	    RECT 155.0000 67.9000 155.4000 69.9000 ;
	    RECT 157.1000 69.2000 157.5000 69.9000 ;
	    RECT 157.1000 68.8000 157.8000 69.2000 ;
	    RECT 157.1000 68.4000 157.5000 68.8000 ;
	    RECT 157.1000 67.9000 157.8000 68.4000 ;
	    RECT 155.1000 67.8000 155.4000 67.9000 ;
	    RECT 155.1000 67.6000 156.0000 67.8000 ;
	    RECT 155.1000 67.5000 157.2000 67.6000 ;
	    RECT 155.7000 67.3000 157.2000 67.5000 ;
	    RECT 156.8000 67.2000 157.2000 67.3000 ;
	    RECT 153.4000 67.1000 154.2000 67.2000 ;
	    RECT 148.7000 66.8000 154.2000 67.1000 ;
	    RECT 147.8000 66.4000 148.2000 66.5000 ;
	    RECT 146.3000 66.1000 148.2000 66.4000 ;
	    RECT 146.3000 66.0000 146.7000 66.1000 ;
	    RECT 147.1000 65.7000 147.5000 65.8000 ;
	    RECT 145.4000 65.4000 147.5000 65.7000 ;
	    RECT 145.4000 61.1000 145.8000 65.4000 ;
	    RECT 148.7000 65.2000 149.0000 66.8000 ;
	    RECT 152.3000 66.7000 152.7000 66.8000 ;
	    RECT 155.0000 66.4000 155.4000 67.2000 ;
	    RECT 156.0000 66.9000 156.4000 67.0000 ;
	    RECT 155.9000 66.6000 156.4000 66.9000 ;
	    RECT 153.1000 66.2000 153.5000 66.3000 ;
	    RECT 155.9000 66.2000 156.2000 66.6000 ;
	    RECT 151.0000 65.9000 153.5000 66.2000 ;
	    RECT 151.0000 65.8000 151.4000 65.9000 ;
	    RECT 155.8000 65.8000 156.2000 66.2000 ;
	    RECT 151.8000 65.5000 154.6000 65.6000 ;
	    RECT 156.8000 65.5000 157.1000 67.2000 ;
	    RECT 157.5000 66.2000 157.8000 67.9000 ;
	    RECT 158.2000 67.5000 158.6000 69.9000 ;
	    RECT 160.4000 69.2000 160.8000 69.9000 ;
	    RECT 159.8000 68.9000 160.8000 69.2000 ;
	    RECT 162.6000 68.9000 163.0000 69.9000 ;
	    RECT 164.7000 69.2000 165.3000 69.9000 ;
	    RECT 164.6000 68.9000 165.3000 69.2000 ;
	    RECT 159.8000 68.5000 160.2000 68.9000 ;
	    RECT 162.6000 68.6000 162.9000 68.9000 ;
	    RECT 160.6000 68.2000 161.0000 68.6000 ;
	    RECT 161.5000 68.3000 162.9000 68.6000 ;
	    RECT 164.6000 68.5000 165.0000 68.9000 ;
	    RECT 161.5000 68.2000 161.9000 68.3000 ;
	    RECT 158.6000 67.1000 159.4000 67.2000 ;
	    RECT 160.7000 67.1000 161.0000 68.2000 ;
	    RECT 165.5000 67.7000 165.9000 67.8000 ;
	    RECT 167.0000 67.7000 167.4000 69.9000 ;
	    RECT 165.5000 67.4000 167.4000 67.7000 ;
	    RECT 163.5000 67.1000 164.2000 67.2000 ;
	    RECT 158.6000 66.8000 164.2000 67.1000 ;
	    RECT 160.1000 66.7000 160.5000 66.8000 ;
	    RECT 157.4000 65.8000 157.8000 66.2000 ;
	    RECT 159.3000 66.2000 159.7000 66.3000 ;
	    RECT 160.6000 66.2000 161.0000 66.3000 ;
	    RECT 159.3000 65.9000 161.8000 66.2000 ;
	    RECT 161.4000 65.8000 161.8000 65.9000 ;
	    RECT 151.7000 65.4000 154.6000 65.5000 ;
	    RECT 147.8000 64.9000 149.0000 65.2000 ;
	    RECT 149.7000 65.3000 154.6000 65.4000 ;
	    RECT 149.7000 65.1000 152.1000 65.3000 ;
	    RECT 147.8000 64.4000 148.1000 64.9000 ;
	    RECT 147.4000 64.0000 148.1000 64.4000 ;
	    RECT 148.9000 64.5000 149.3000 64.6000 ;
	    RECT 149.7000 64.5000 150.0000 65.1000 ;
	    RECT 148.9000 64.2000 150.0000 64.5000 ;
	    RECT 150.3000 64.5000 153.0000 64.8000 ;
	    RECT 150.3000 64.4000 150.7000 64.5000 ;
	    RECT 152.6000 64.4000 153.0000 64.5000 ;
	    RECT 149.5000 63.7000 149.9000 63.8000 ;
	    RECT 150.9000 63.7000 151.3000 63.8000 ;
	    RECT 147.8000 63.1000 148.2000 63.5000 ;
	    RECT 149.5000 63.4000 151.3000 63.7000 ;
	    RECT 149.9000 63.1000 150.2000 63.4000 ;
	    RECT 152.6000 63.1000 153.0000 63.5000 ;
	    RECT 147.5000 61.1000 148.1000 63.1000 ;
	    RECT 149.8000 61.1000 150.2000 63.1000 ;
	    RECT 152.0000 62.8000 153.0000 63.1000 ;
	    RECT 152.0000 61.1000 152.4000 62.8000 ;
	    RECT 154.2000 61.1000 154.6000 65.3000 ;
	    RECT 155.9000 65.2000 157.1000 65.5000 ;
	    RECT 155.9000 63.1000 156.2000 65.2000 ;
	    RECT 157.5000 65.1000 157.8000 65.8000 ;
	    RECT 155.8000 61.1000 156.2000 63.1000 ;
	    RECT 157.4000 61.1000 157.8000 65.1000 ;
	    RECT 158.2000 65.5000 161.0000 65.6000 ;
	    RECT 158.2000 65.4000 161.1000 65.5000 ;
	    RECT 158.2000 65.3000 163.1000 65.4000 ;
	    RECT 158.2000 61.1000 158.6000 65.3000 ;
	    RECT 160.7000 65.1000 163.1000 65.3000 ;
	    RECT 159.8000 64.5000 162.5000 64.8000 ;
	    RECT 159.8000 64.4000 160.2000 64.5000 ;
	    RECT 162.1000 64.4000 162.5000 64.5000 ;
	    RECT 162.8000 64.5000 163.1000 65.1000 ;
	    RECT 163.8000 65.2000 164.1000 66.8000 ;
	    RECT 164.6000 66.4000 165.0000 66.5000 ;
	    RECT 164.6000 66.1000 166.5000 66.4000 ;
	    RECT 166.1000 66.0000 166.5000 66.1000 ;
	    RECT 165.3000 65.7000 165.7000 65.8000 ;
	    RECT 167.0000 65.7000 167.4000 67.4000 ;
	    RECT 167.8000 67.6000 168.2000 69.9000 ;
	    RECT 170.2000 67.6000 170.6000 69.9000 ;
	    RECT 167.8000 67.3000 168.9000 67.6000 ;
	    RECT 170.2000 67.3000 171.3000 67.6000 ;
	    RECT 167.8000 65.8000 168.2000 66.6000 ;
	    RECT 168.6000 65.8000 168.9000 67.3000 ;
	    RECT 170.2000 65.8000 170.6000 66.6000 ;
	    RECT 171.0000 65.8000 171.3000 67.3000 ;
	    RECT 165.3000 65.4000 167.4000 65.7000 ;
	    RECT 163.8000 64.9000 165.0000 65.2000 ;
	    RECT 163.5000 64.5000 163.9000 64.6000 ;
	    RECT 162.8000 64.2000 163.9000 64.5000 ;
	    RECT 164.7000 64.4000 165.0000 64.9000 ;
	    RECT 164.7000 64.0000 165.4000 64.4000 ;
	    RECT 161.5000 63.7000 161.9000 63.8000 ;
	    RECT 162.9000 63.7000 163.3000 63.8000 ;
	    RECT 159.8000 63.1000 160.2000 63.5000 ;
	    RECT 161.5000 63.4000 163.3000 63.7000 ;
	    RECT 162.6000 63.1000 162.9000 63.4000 ;
	    RECT 164.6000 63.1000 165.0000 63.5000 ;
	    RECT 159.8000 62.8000 160.8000 63.1000 ;
	    RECT 160.4000 61.1000 160.8000 62.8000 ;
	    RECT 162.6000 61.1000 163.0000 63.1000 ;
	    RECT 164.7000 61.1000 165.3000 63.1000 ;
	    RECT 167.0000 61.1000 167.4000 65.4000 ;
	    RECT 168.6000 65.4000 169.2000 65.8000 ;
	    RECT 171.0000 65.4000 171.6000 65.8000 ;
	    RECT 168.6000 65.1000 168.9000 65.4000 ;
	    RECT 171.0000 65.1000 171.3000 65.4000 ;
	    RECT 167.8000 64.8000 168.9000 65.1000 ;
	    RECT 170.2000 64.8000 171.3000 65.1000 ;
	    RECT 167.8000 61.1000 168.2000 64.8000 ;
	    RECT 170.2000 61.1000 170.6000 64.8000 ;
	    RECT 0.6000 57.9000 1.0000 59.9000 ;
	    RECT 0.7000 57.8000 1.0000 57.9000 ;
	    RECT 2.2000 57.9000 2.6000 59.9000 ;
	    RECT 3.8000 57.9000 4.2000 59.9000 ;
	    RECT 2.2000 57.8000 2.5000 57.9000 ;
	    RECT 0.7000 57.5000 2.5000 57.8000 ;
	    RECT 3.9000 57.8000 4.2000 57.9000 ;
	    RECT 5.4000 57.8000 5.8000 59.9000 ;
	    RECT 3.9000 57.5000 5.7000 57.8000 ;
	    RECT 0.7000 56.2000 1.0000 57.5000 ;
	    RECT 1.4000 56.4000 1.8000 57.2000 ;
	    RECT 3.9000 56.2000 4.2000 57.5000 ;
	    RECT 4.6000 56.4000 5.0000 57.2000 ;
	    RECT 0.6000 55.8000 1.0000 56.2000 ;
	    RECT 0.7000 54.2000 1.0000 55.8000 ;
	    RECT 3.0000 55.4000 3.4000 56.2000 ;
	    RECT 3.8000 55.8000 4.2000 56.2000 ;
	    RECT 1.8000 54.8000 2.6000 55.2000 ;
	    RECT 3.9000 54.2000 4.2000 55.8000 ;
	    RECT 6.2000 55.4000 6.6000 56.2000 ;
	    RECT 5.0000 54.8000 5.8000 55.2000 ;
	    RECT 0.7000 54.1000 1.5000 54.2000 ;
	    RECT 3.9000 54.1000 4.7000 54.2000 ;
	    RECT 0.7000 53.9000 2.5000 54.1000 ;
	    RECT 3.9000 53.9000 4.8000 54.1000 ;
	    RECT 1.2000 53.8000 2.5000 53.9000 ;
	    RECT 1.2000 51.1000 1.6000 53.8000 ;
	    RECT 2.2000 53.2000 2.5000 53.8000 ;
	    RECT 2.2000 52.8000 2.6000 53.2000 ;
	    RECT 4.4000 51.1000 4.8000 53.9000 ;
	    RECT 7.8000 51.1000 8.2000 59.9000 ;
	    RECT 8.6000 54.1000 9.0000 59.9000 ;
	    RECT 11.5000 56.2000 11.9000 59.9000 ;
	    RECT 13.4000 57.9000 13.8000 59.9000 ;
	    RECT 13.5000 57.8000 13.8000 57.9000 ;
	    RECT 15.0000 57.8000 15.4000 59.9000 ;
	    RECT 16.6000 57.9000 17.0000 59.9000 ;
	    RECT 16.7000 57.8000 17.0000 57.9000 ;
	    RECT 18.2000 57.9000 18.6000 59.9000 ;
	    RECT 20.6000 57.9000 21.0000 59.9000 ;
	    RECT 18.2000 57.8000 18.5000 57.9000 ;
	    RECT 13.5000 57.5000 15.3000 57.8000 ;
	    RECT 16.7000 57.5000 18.5000 57.8000 ;
	    RECT 20.7000 57.8000 21.0000 57.9000 ;
	    RECT 22.2000 57.9000 22.6000 59.9000 ;
	    RECT 23.8000 57.9000 24.2000 59.9000 ;
	    RECT 22.2000 57.8000 22.5000 57.9000 ;
	    RECT 20.7000 57.5000 22.5000 57.8000 ;
	    RECT 23.9000 57.8000 24.2000 57.9000 ;
	    RECT 25.4000 57.9000 25.8000 59.9000 ;
	    RECT 27.0000 57.9000 27.4000 59.9000 ;
	    RECT 25.4000 57.8000 25.7000 57.9000 ;
	    RECT 23.9000 57.5000 25.7000 57.8000 ;
	    RECT 27.1000 57.8000 27.4000 57.9000 ;
	    RECT 28.6000 57.9000 29.0000 59.9000 ;
	    RECT 28.6000 57.8000 28.9000 57.9000 ;
	    RECT 27.1000 57.5000 28.9000 57.8000 ;
	    RECT 12.2000 56.8000 12.6000 57.2000 ;
	    RECT 12.3000 56.2000 12.6000 56.8000 ;
	    RECT 13.5000 56.2000 13.8000 57.5000 ;
	    RECT 14.2000 56.4000 14.6000 57.2000 ;
	    RECT 16.7000 56.2000 17.0000 57.5000 ;
	    RECT 17.4000 57.1000 17.8000 57.2000 ;
	    RECT 19.0000 57.1000 19.4000 57.2000 ;
	    RECT 17.4000 56.8000 19.4000 57.1000 ;
	    RECT 17.4000 56.4000 17.8000 56.8000 ;
	    RECT 21.4000 56.4000 21.8000 57.2000 ;
	    RECT 22.2000 56.2000 22.5000 57.5000 ;
	    RECT 24.6000 56.4000 25.0000 57.2000 ;
	    RECT 25.4000 56.2000 25.7000 57.5000 ;
	    RECT 27.8000 56.4000 28.2000 57.2000 ;
	    RECT 28.6000 56.2000 28.9000 57.5000 ;
	    RECT 29.7000 56.2000 30.1000 59.9000 ;
	    RECT 11.5000 55.9000 12.0000 56.2000 ;
	    RECT 12.3000 55.9000 13.0000 56.2000 ;
	    RECT 11.0000 54.4000 11.4000 55.2000 ;
	    RECT 11.7000 54.2000 12.0000 55.9000 ;
	    RECT 12.6000 55.8000 13.0000 55.9000 ;
	    RECT 13.4000 55.8000 13.8000 56.2000 ;
	    RECT 13.5000 54.2000 13.8000 55.8000 ;
	    RECT 15.8000 55.4000 16.2000 56.2000 ;
	    RECT 16.6000 55.8000 17.0000 56.2000 ;
	    RECT 14.6000 54.8000 15.4000 55.2000 ;
	    RECT 16.7000 54.2000 17.0000 55.8000 ;
	    RECT 17.8000 54.8000 18.6000 55.2000 ;
	    RECT 19.0000 54.8000 19.4000 56.2000 ;
	    RECT 19.8000 55.4000 20.2000 56.2000 ;
	    RECT 22.2000 55.8000 22.6000 56.2000 ;
	    RECT 20.6000 54.8000 21.4000 55.2000 ;
	    RECT 22.2000 54.2000 22.5000 55.8000 ;
	    RECT 23.0000 55.4000 23.4000 56.2000 ;
	    RECT 25.4000 55.8000 25.8000 56.2000 ;
	    RECT 28.6000 55.8000 29.0000 56.2000 ;
	    RECT 29.4000 55.9000 30.1000 56.2000 ;
	    RECT 23.8000 54.8000 24.6000 55.2000 ;
	    RECT 25.4000 54.2000 25.7000 55.8000 ;
	    RECT 27.0000 54.8000 27.8000 55.2000 ;
	    RECT 28.6000 54.2000 28.9000 55.8000 ;
	    RECT 10.2000 54.1000 10.6000 54.2000 ;
	    RECT 8.6000 53.8000 11.0000 54.1000 ;
	    RECT 11.7000 53.8000 13.0000 54.2000 ;
	    RECT 13.5000 54.1000 14.3000 54.2000 ;
	    RECT 16.6000 54.1000 17.5000 54.2000 ;
	    RECT 21.7000 54.1000 22.5000 54.2000 ;
	    RECT 24.9000 54.1000 25.7000 54.2000 ;
	    RECT 28.1000 54.1000 28.9000 54.2000 ;
	    RECT 13.5000 53.9000 14.4000 54.1000 ;
	    RECT 8.6000 51.1000 9.0000 53.8000 ;
	    RECT 10.6000 53.6000 11.0000 53.8000 ;
	    RECT 10.3000 53.1000 12.1000 53.3000 ;
	    RECT 12.6000 53.1000 12.9000 53.8000 ;
	    RECT 10.2000 53.0000 12.2000 53.1000 ;
	    RECT 10.2000 51.1000 10.6000 53.0000 ;
	    RECT 11.8000 51.1000 12.2000 53.0000 ;
	    RECT 12.6000 51.1000 13.0000 53.1000 ;
	    RECT 14.0000 51.1000 14.4000 53.9000 ;
	    RECT 16.6000 53.8000 17.6000 54.1000 ;
	    RECT 17.2000 51.1000 17.6000 53.8000 ;
	    RECT 21.6000 53.9000 22.5000 54.1000 ;
	    RECT 24.8000 53.9000 25.7000 54.1000 ;
	    RECT 28.0000 53.9000 28.9000 54.1000 ;
	    RECT 29.4000 55.2000 29.7000 55.9000 ;
	    RECT 31.8000 55.6000 32.2000 59.9000 ;
	    RECT 32.6000 56.2000 33.0000 59.9000 ;
	    RECT 34.2000 56.2000 34.6000 59.9000 ;
	    RECT 32.6000 55.9000 34.6000 56.2000 ;
	    RECT 30.2000 55.4000 32.2000 55.6000 ;
	    RECT 35.0000 55.8000 35.4000 59.9000 ;
	    RECT 35.8000 56.2000 36.2000 59.9000 ;
	    RECT 37.4000 56.2000 37.8000 59.9000 ;
	    RECT 35.8000 55.9000 37.8000 56.2000 ;
	    RECT 38.2000 55.8000 38.6000 59.9000 ;
	    RECT 39.0000 56.2000 39.4000 59.9000 ;
	    RECT 40.6000 56.2000 41.0000 59.9000 ;
	    RECT 39.0000 55.9000 41.0000 56.2000 ;
	    RECT 41.4000 55.8000 41.8000 59.9000 ;
	    RECT 42.2000 56.2000 42.6000 59.9000 ;
	    RECT 43.8000 56.2000 44.2000 59.9000 ;
	    RECT 42.2000 55.9000 44.2000 56.2000 ;
	    RECT 44.6000 55.9000 45.0000 59.9000 ;
	    RECT 30.1000 55.3000 32.2000 55.4000 ;
	    RECT 29.4000 54.8000 29.8000 55.2000 ;
	    RECT 30.1000 55.0000 30.5000 55.3000 ;
	    RECT 33.0000 55.2000 33.4000 55.4000 ;
	    RECT 35.0000 55.2000 35.3000 55.8000 ;
	    RECT 36.2000 55.2000 36.6000 55.4000 ;
	    RECT 38.2000 55.2000 38.5000 55.8000 ;
	    RECT 39.4000 55.2000 39.8000 55.4000 ;
	    RECT 41.4000 55.2000 41.7000 55.8000 ;
	    RECT 42.6000 55.2000 43.0000 55.4000 ;
	    RECT 44.6000 55.2000 44.9000 55.9000 ;
	    RECT 21.6000 53.2000 22.0000 53.9000 ;
	    RECT 21.6000 52.8000 22.6000 53.2000 ;
	    RECT 21.6000 51.1000 22.0000 52.8000 ;
	    RECT 24.8000 51.1000 25.2000 53.9000 ;
	    RECT 28.0000 51.1000 28.4000 53.9000 ;
	    RECT 29.4000 53.1000 29.7000 54.8000 ;
	    RECT 30.1000 53.5000 30.4000 55.0000 ;
	    RECT 32.6000 54.9000 33.4000 55.2000 ;
	    RECT 34.2000 54.9000 35.4000 55.2000 ;
	    RECT 32.6000 54.8000 33.0000 54.9000 ;
	    RECT 33.4000 53.8000 33.8000 54.6000 ;
	    RECT 30.1000 53.2000 31.3000 53.5000 ;
	    RECT 29.4000 51.1000 29.8000 53.1000 ;
	    RECT 31.0000 52.1000 31.3000 53.2000 ;
	    RECT 31.8000 52.4000 32.2000 53.2000 ;
	    RECT 34.2000 53.1000 34.5000 54.9000 ;
	    RECT 35.0000 54.8000 35.4000 54.9000 ;
	    RECT 35.8000 54.9000 36.6000 55.2000 ;
	    RECT 37.4000 54.9000 38.6000 55.2000 ;
	    RECT 35.8000 54.8000 36.2000 54.9000 ;
	    RECT 36.6000 53.8000 37.0000 54.6000 ;
	    RECT 31.0000 51.1000 31.4000 52.1000 ;
	    RECT 34.2000 51.1000 34.6000 53.1000 ;
	    RECT 35.0000 52.8000 35.4000 53.2000 ;
	    RECT 37.4000 53.1000 37.7000 54.9000 ;
	    RECT 38.2000 54.8000 38.6000 54.9000 ;
	    RECT 39.0000 54.9000 39.8000 55.2000 ;
	    RECT 40.6000 54.9000 41.8000 55.2000 ;
	    RECT 39.0000 54.8000 39.4000 54.9000 ;
	    RECT 39.8000 53.8000 40.2000 54.6000 ;
	    RECT 34.9000 52.4000 35.3000 52.8000 ;
	    RECT 37.4000 51.1000 37.8000 53.1000 ;
	    RECT 38.2000 52.8000 38.6000 53.2000 ;
	    RECT 40.6000 53.1000 40.9000 54.9000 ;
	    RECT 41.4000 54.8000 41.8000 54.9000 ;
	    RECT 42.2000 54.9000 43.0000 55.2000 ;
	    RECT 43.8000 54.9000 45.0000 55.2000 ;
	    RECT 42.2000 54.8000 42.6000 54.9000 ;
	    RECT 41.4000 53.8000 41.8000 54.2000 ;
	    RECT 43.0000 53.8000 43.4000 54.6000 ;
	    RECT 41.4000 53.2000 41.7000 53.8000 ;
	    RECT 38.1000 52.4000 38.5000 52.8000 ;
	    RECT 40.6000 51.1000 41.0000 53.1000 ;
	    RECT 41.4000 52.8000 41.8000 53.2000 ;
	    RECT 43.8000 53.1000 44.1000 54.9000 ;
	    RECT 44.6000 54.8000 45.0000 54.9000 ;
	    RECT 44.6000 53.1000 45.0000 53.2000 ;
	    RECT 45.4000 53.1000 45.8000 59.9000 ;
	    RECT 47.0000 55.7000 47.4000 59.9000 ;
	    RECT 49.2000 58.2000 49.6000 59.9000 ;
	    RECT 48.6000 57.9000 49.6000 58.2000 ;
	    RECT 51.4000 57.9000 51.8000 59.9000 ;
	    RECT 53.5000 57.9000 54.1000 59.9000 ;
	    RECT 48.6000 57.5000 49.0000 57.9000 ;
	    RECT 51.4000 57.6000 51.7000 57.9000 ;
	    RECT 50.3000 57.3000 52.1000 57.6000 ;
	    RECT 53.4000 57.5000 53.8000 57.9000 ;
	    RECT 50.3000 57.2000 50.7000 57.3000 ;
	    RECT 51.7000 57.2000 52.1000 57.3000 ;
	    RECT 48.6000 56.5000 49.0000 56.6000 ;
	    RECT 50.9000 56.5000 51.3000 56.6000 ;
	    RECT 48.6000 56.2000 51.3000 56.5000 ;
	    RECT 51.6000 56.5000 52.7000 56.8000 ;
	    RECT 51.6000 55.9000 51.9000 56.5000 ;
	    RECT 52.3000 56.4000 52.7000 56.5000 ;
	    RECT 53.5000 56.6000 54.2000 57.0000 ;
	    RECT 53.5000 56.1000 53.8000 56.6000 ;
	    RECT 49.5000 55.7000 51.9000 55.9000 ;
	    RECT 47.0000 55.6000 51.9000 55.7000 ;
	    RECT 52.6000 55.8000 53.8000 56.1000 ;
	    RECT 47.0000 55.5000 49.9000 55.6000 ;
	    RECT 47.0000 55.4000 49.8000 55.5000 ;
	    RECT 52.6000 55.2000 52.9000 55.8000 ;
	    RECT 55.8000 55.6000 56.2000 59.9000 ;
	    RECT 56.6000 57.9000 57.0000 59.9000 ;
	    RECT 56.7000 57.8000 57.0000 57.9000 ;
	    RECT 58.2000 57.9000 58.6000 59.9000 ;
	    RECT 58.2000 57.8000 58.5000 57.9000 ;
	    RECT 56.7000 57.5000 58.5000 57.8000 ;
	    RECT 56.7000 56.2000 57.0000 57.5000 ;
	    RECT 57.4000 56.4000 57.8000 57.2000 ;
	    RECT 56.6000 55.8000 57.0000 56.2000 ;
	    RECT 54.1000 55.3000 56.2000 55.6000 ;
	    RECT 54.1000 55.2000 54.5000 55.3000 ;
	    RECT 50.2000 55.1000 50.6000 55.2000 ;
	    RECT 48.1000 54.8000 50.6000 55.1000 ;
	    RECT 52.6000 54.8000 53.0000 55.2000 ;
	    RECT 54.9000 54.9000 55.3000 55.0000 ;
	    RECT 48.1000 54.7000 48.5000 54.8000 ;
	    RECT 49.4000 54.7000 49.8000 54.8000 ;
	    RECT 48.9000 54.2000 49.3000 54.3000 ;
	    RECT 52.6000 54.2000 52.9000 54.8000 ;
	    RECT 53.4000 54.6000 55.3000 54.9000 ;
	    RECT 53.4000 54.5000 53.8000 54.6000 ;
	    RECT 46.2000 53.4000 46.6000 54.2000 ;
	    RECT 47.4000 53.9000 52.9000 54.2000 ;
	    RECT 47.4000 53.8000 48.2000 53.9000 ;
	    RECT 41.3000 52.4000 41.7000 52.8000 ;
	    RECT 43.8000 51.1000 44.2000 53.1000 ;
	    RECT 44.6000 52.8000 45.8000 53.1000 ;
	    RECT 44.5000 52.4000 44.9000 52.8000 ;
	    RECT 45.4000 51.1000 45.8000 52.8000 ;
	    RECT 47.0000 51.1000 47.4000 53.5000 ;
	    RECT 49.5000 52.8000 49.8000 53.9000 ;
	    RECT 52.3000 53.8000 52.7000 53.9000 ;
	    RECT 55.8000 53.6000 56.2000 55.3000 ;
	    RECT 56.7000 54.2000 57.0000 55.8000 ;
	    RECT 61.4000 55.7000 61.8000 59.9000 ;
	    RECT 63.6000 58.2000 64.0000 59.9000 ;
	    RECT 63.0000 57.9000 64.0000 58.2000 ;
	    RECT 65.8000 57.9000 66.2000 59.9000 ;
	    RECT 67.9000 57.9000 68.5000 59.9000 ;
	    RECT 63.0000 57.5000 63.4000 57.9000 ;
	    RECT 65.8000 57.6000 66.1000 57.9000 ;
	    RECT 64.7000 57.3000 66.5000 57.6000 ;
	    RECT 67.8000 57.5000 68.2000 57.9000 ;
	    RECT 64.7000 57.2000 65.1000 57.3000 ;
	    RECT 66.1000 57.2000 66.5000 57.3000 ;
	    RECT 63.0000 56.5000 63.4000 56.6000 ;
	    RECT 65.3000 56.5000 65.7000 56.6000 ;
	    RECT 63.0000 56.2000 65.7000 56.5000 ;
	    RECT 66.0000 56.5000 67.1000 56.8000 ;
	    RECT 66.0000 55.9000 66.3000 56.5000 ;
	    RECT 66.7000 56.4000 67.1000 56.5000 ;
	    RECT 67.9000 56.6000 68.6000 57.0000 ;
	    RECT 67.9000 56.1000 68.2000 56.6000 ;
	    RECT 63.9000 55.7000 66.3000 55.9000 ;
	    RECT 61.4000 55.6000 66.3000 55.7000 ;
	    RECT 67.0000 55.8000 68.2000 56.1000 ;
	    RECT 61.4000 55.5000 64.3000 55.6000 ;
	    RECT 61.4000 55.4000 64.2000 55.5000 ;
	    RECT 67.0000 55.2000 67.3000 55.8000 ;
	    RECT 70.2000 55.6000 70.6000 59.9000 ;
	    RECT 71.0000 57.9000 71.4000 59.9000 ;
	    RECT 71.1000 57.8000 71.4000 57.9000 ;
	    RECT 72.6000 57.9000 73.0000 59.9000 ;
	    RECT 74.2000 57.9000 74.6000 59.9000 ;
	    RECT 72.6000 57.8000 72.9000 57.9000 ;
	    RECT 71.1000 57.5000 72.9000 57.8000 ;
	    RECT 74.3000 57.8000 74.6000 57.9000 ;
	    RECT 75.8000 57.9000 76.2000 59.9000 ;
	    RECT 78.2000 57.9000 78.6000 59.9000 ;
	    RECT 75.8000 57.8000 76.1000 57.9000 ;
	    RECT 74.3000 57.5000 76.1000 57.8000 ;
	    RECT 78.3000 57.8000 78.6000 57.9000 ;
	    RECT 79.8000 57.9000 80.2000 59.9000 ;
	    RECT 79.8000 57.8000 80.1000 57.9000 ;
	    RECT 78.3000 57.5000 80.1000 57.8000 ;
	    RECT 71.1000 56.2000 71.4000 57.5000 ;
	    RECT 71.8000 56.4000 72.2000 57.2000 ;
	    RECT 74.3000 56.2000 74.6000 57.5000 ;
	    RECT 75.0000 56.4000 75.4000 57.2000 ;
	    RECT 79.0000 56.4000 79.4000 57.2000 ;
	    RECT 71.0000 55.8000 71.4000 56.2000 ;
	    RECT 74.2000 55.8000 74.6000 56.2000 ;
	    RECT 68.5000 55.3000 70.6000 55.6000 ;
	    RECT 68.5000 55.2000 68.9000 55.3000 ;
	    RECT 57.8000 54.8000 58.6000 55.2000 ;
	    RECT 64.6000 55.1000 65.0000 55.2000 ;
	    RECT 62.5000 54.8000 65.0000 55.1000 ;
	    RECT 67.0000 54.8000 67.4000 55.2000 ;
	    RECT 69.3000 54.9000 69.7000 55.0000 ;
	    RECT 62.5000 54.7000 62.9000 54.8000 ;
	    RECT 63.8000 54.7000 64.2000 54.8000 ;
	    RECT 63.3000 54.2000 63.7000 54.3000 ;
	    RECT 67.0000 54.2000 67.3000 54.8000 ;
	    RECT 67.8000 54.6000 69.7000 54.9000 ;
	    RECT 67.8000 54.5000 68.2000 54.6000 ;
	    RECT 56.7000 54.1000 57.5000 54.2000 ;
	    RECT 56.7000 53.9000 57.6000 54.1000 ;
	    RECT 54.3000 53.3000 56.2000 53.6000 ;
	    RECT 54.3000 53.2000 54.7000 53.3000 ;
	    RECT 48.6000 52.1000 49.0000 52.5000 ;
	    RECT 49.4000 52.4000 49.8000 52.8000 ;
	    RECT 50.3000 52.7000 50.7000 52.8000 ;
	    RECT 50.3000 52.4000 51.7000 52.7000 ;
	    RECT 51.4000 52.1000 51.7000 52.4000 ;
	    RECT 53.4000 52.1000 53.8000 52.5000 ;
	    RECT 48.6000 51.8000 49.6000 52.1000 ;
	    RECT 49.2000 51.1000 49.6000 51.8000 ;
	    RECT 51.4000 51.1000 51.8000 52.1000 ;
	    RECT 53.4000 51.8000 54.1000 52.1000 ;
	    RECT 53.5000 51.1000 54.1000 51.8000 ;
	    RECT 55.8000 51.1000 56.2000 53.3000 ;
	    RECT 57.2000 51.1000 57.6000 53.9000 ;
	    RECT 61.8000 53.9000 67.3000 54.2000 ;
	    RECT 61.8000 53.8000 62.6000 53.9000 ;
	    RECT 61.4000 51.1000 61.8000 53.5000 ;
	    RECT 63.9000 52.8000 64.2000 53.9000 ;
	    RECT 66.7000 53.8000 67.1000 53.9000 ;
	    RECT 70.2000 53.6000 70.6000 55.3000 ;
	    RECT 71.1000 54.2000 71.4000 55.8000 ;
	    RECT 72.2000 54.8000 73.0000 55.2000 ;
	    RECT 74.3000 54.2000 74.6000 55.8000 ;
	    RECT 79.8000 56.2000 80.1000 57.5000 ;
	    RECT 79.8000 55.8000 80.2000 56.2000 ;
	    RECT 75.4000 54.8000 76.2000 55.2000 ;
	    RECT 78.2000 54.8000 79.0000 55.2000 ;
	    RECT 79.8000 54.2000 80.1000 55.8000 ;
	    RECT 80.6000 55.7000 81.0000 59.9000 ;
	    RECT 82.8000 58.2000 83.2000 59.9000 ;
	    RECT 82.2000 57.9000 83.2000 58.2000 ;
	    RECT 85.0000 57.9000 85.4000 59.9000 ;
	    RECT 87.1000 57.9000 87.7000 59.9000 ;
	    RECT 82.2000 57.5000 82.6000 57.9000 ;
	    RECT 85.0000 57.6000 85.3000 57.9000 ;
	    RECT 83.9000 57.3000 85.7000 57.6000 ;
	    RECT 87.0000 57.5000 87.4000 57.9000 ;
	    RECT 83.9000 57.2000 84.3000 57.3000 ;
	    RECT 85.3000 57.2000 85.7000 57.3000 ;
	    RECT 82.2000 56.5000 82.6000 56.6000 ;
	    RECT 84.5000 56.5000 84.9000 56.6000 ;
	    RECT 82.2000 56.2000 84.9000 56.5000 ;
	    RECT 85.2000 56.5000 86.3000 56.8000 ;
	    RECT 85.2000 55.9000 85.5000 56.5000 ;
	    RECT 85.9000 56.4000 86.3000 56.5000 ;
	    RECT 87.1000 56.6000 87.8000 57.0000 ;
	    RECT 87.1000 56.1000 87.4000 56.6000 ;
	    RECT 83.1000 55.7000 85.5000 55.9000 ;
	    RECT 80.6000 55.6000 85.5000 55.7000 ;
	    RECT 86.2000 55.8000 87.4000 56.1000 ;
	    RECT 80.6000 55.5000 83.5000 55.6000 ;
	    RECT 80.6000 55.4000 83.4000 55.5000 ;
	    RECT 86.2000 55.2000 86.5000 55.8000 ;
	    RECT 89.4000 55.6000 89.8000 59.9000 ;
	    RECT 87.7000 55.3000 89.8000 55.6000 ;
	    RECT 90.2000 55.7000 90.6000 59.9000 ;
	    RECT 92.4000 58.2000 92.8000 59.9000 ;
	    RECT 91.8000 57.9000 92.8000 58.2000 ;
	    RECT 94.6000 57.9000 95.0000 59.9000 ;
	    RECT 96.7000 57.9000 97.3000 59.9000 ;
	    RECT 91.8000 57.5000 92.2000 57.9000 ;
	    RECT 94.6000 57.6000 94.9000 57.9000 ;
	    RECT 93.5000 57.3000 95.3000 57.6000 ;
	    RECT 96.6000 57.5000 97.0000 57.9000 ;
	    RECT 93.5000 57.2000 93.9000 57.3000 ;
	    RECT 94.9000 57.2000 95.3000 57.3000 ;
	    RECT 91.8000 56.5000 92.2000 56.6000 ;
	    RECT 94.1000 56.5000 94.5000 56.6000 ;
	    RECT 91.8000 56.2000 94.5000 56.5000 ;
	    RECT 94.8000 56.5000 95.9000 56.8000 ;
	    RECT 94.8000 55.9000 95.1000 56.5000 ;
	    RECT 95.5000 56.4000 95.9000 56.5000 ;
	    RECT 96.7000 56.6000 97.4000 57.0000 ;
	    RECT 96.7000 56.1000 97.0000 56.6000 ;
	    RECT 92.7000 55.7000 95.1000 55.9000 ;
	    RECT 90.2000 55.6000 95.1000 55.7000 ;
	    RECT 95.8000 55.8000 97.0000 56.1000 ;
	    RECT 90.2000 55.5000 93.1000 55.6000 ;
	    RECT 90.2000 55.4000 93.0000 55.5000 ;
	    RECT 87.7000 55.2000 88.1000 55.3000 ;
	    RECT 83.8000 55.1000 84.2000 55.2000 ;
	    RECT 81.7000 54.8000 84.2000 55.1000 ;
	    RECT 86.2000 54.8000 86.6000 55.2000 ;
	    RECT 88.5000 54.9000 88.9000 55.0000 ;
	    RECT 81.7000 54.7000 82.1000 54.8000 ;
	    RECT 83.0000 54.7000 83.4000 54.8000 ;
	    RECT 82.5000 54.2000 82.9000 54.3000 ;
	    RECT 86.2000 54.2000 86.5000 54.8000 ;
	    RECT 87.0000 54.6000 88.9000 54.9000 ;
	    RECT 87.0000 54.5000 87.4000 54.6000 ;
	    RECT 71.1000 54.1000 71.9000 54.2000 ;
	    RECT 74.3000 54.1000 75.1000 54.2000 ;
	    RECT 79.3000 54.1000 80.1000 54.2000 ;
	    RECT 71.1000 53.9000 72.0000 54.1000 ;
	    RECT 74.3000 53.9000 75.2000 54.1000 ;
	    RECT 68.7000 53.3000 70.6000 53.6000 ;
	    RECT 68.7000 53.2000 69.1000 53.3000 ;
	    RECT 63.0000 52.1000 63.4000 52.5000 ;
	    RECT 63.8000 52.4000 64.2000 52.8000 ;
	    RECT 64.7000 52.7000 65.1000 52.8000 ;
	    RECT 64.7000 52.4000 66.1000 52.7000 ;
	    RECT 65.8000 52.1000 66.1000 52.4000 ;
	    RECT 67.8000 52.1000 68.2000 52.5000 ;
	    RECT 63.0000 51.8000 64.0000 52.1000 ;
	    RECT 63.6000 51.1000 64.0000 51.8000 ;
	    RECT 65.8000 51.1000 66.2000 52.1000 ;
	    RECT 67.8000 51.8000 68.5000 52.1000 ;
	    RECT 67.9000 51.1000 68.5000 51.8000 ;
	    RECT 70.2000 51.1000 70.6000 53.3000 ;
	    RECT 71.6000 51.1000 72.0000 53.9000 ;
	    RECT 74.8000 51.1000 75.2000 53.9000 ;
	    RECT 79.2000 53.9000 80.1000 54.1000 ;
	    RECT 81.0000 53.9000 86.5000 54.2000 ;
	    RECT 79.2000 51.1000 79.6000 53.9000 ;
	    RECT 81.0000 53.8000 81.8000 53.9000 ;
	    RECT 80.6000 51.1000 81.0000 53.5000 ;
	    RECT 83.1000 52.8000 83.4000 53.9000 ;
	    RECT 85.9000 53.8000 86.3000 53.9000 ;
	    RECT 89.4000 53.6000 89.8000 55.3000 ;
	    RECT 95.8000 55.2000 96.1000 55.8000 ;
	    RECT 99.0000 55.6000 99.4000 59.9000 ;
	    RECT 97.3000 55.3000 99.4000 55.6000 ;
	    RECT 97.3000 55.2000 97.7000 55.3000 ;
	    RECT 93.4000 55.1000 93.8000 55.2000 ;
	    RECT 95.0000 55.1000 95.4000 55.2000 ;
	    RECT 91.3000 54.8000 95.4000 55.1000 ;
	    RECT 95.8000 54.8000 96.2000 55.2000 ;
	    RECT 98.1000 54.9000 98.5000 55.0000 ;
	    RECT 91.3000 54.7000 91.7000 54.8000 ;
	    RECT 92.1000 54.2000 92.5000 54.3000 ;
	    RECT 95.8000 54.2000 96.1000 54.8000 ;
	    RECT 96.6000 54.6000 98.5000 54.9000 ;
	    RECT 96.6000 54.5000 97.0000 54.6000 ;
	    RECT 90.6000 53.9000 96.1000 54.2000 ;
	    RECT 90.6000 53.8000 91.4000 53.9000 ;
	    RECT 87.9000 53.3000 89.8000 53.6000 ;
	    RECT 87.9000 53.2000 88.3000 53.3000 ;
	    RECT 82.2000 52.1000 82.6000 52.5000 ;
	    RECT 83.0000 52.4000 83.4000 52.8000 ;
	    RECT 83.9000 52.7000 84.3000 52.8000 ;
	    RECT 83.9000 52.4000 85.3000 52.7000 ;
	    RECT 85.0000 52.1000 85.3000 52.4000 ;
	    RECT 87.0000 52.1000 87.4000 52.5000 ;
	    RECT 82.2000 51.8000 83.2000 52.1000 ;
	    RECT 82.8000 51.1000 83.2000 51.8000 ;
	    RECT 85.0000 51.1000 85.4000 52.1000 ;
	    RECT 87.0000 51.8000 87.7000 52.1000 ;
	    RECT 87.1000 51.1000 87.7000 51.8000 ;
	    RECT 89.4000 51.1000 89.8000 53.3000 ;
	    RECT 90.2000 51.1000 90.6000 53.5000 ;
	    RECT 92.7000 52.8000 93.0000 53.9000 ;
	    RECT 95.5000 53.8000 95.9000 53.9000 ;
	    RECT 99.0000 53.6000 99.4000 55.3000 ;
	    RECT 97.5000 53.3000 99.4000 53.6000 ;
	    RECT 97.5000 53.2000 97.9000 53.3000 ;
	    RECT 91.8000 52.1000 92.2000 52.5000 ;
	    RECT 92.6000 52.4000 93.0000 52.8000 ;
	    RECT 93.5000 52.7000 93.9000 52.8000 ;
	    RECT 93.5000 52.4000 94.9000 52.7000 ;
	    RECT 94.6000 52.1000 94.9000 52.4000 ;
	    RECT 96.6000 52.1000 97.0000 52.5000 ;
	    RECT 91.8000 51.8000 92.8000 52.1000 ;
	    RECT 92.4000 51.1000 92.8000 51.8000 ;
	    RECT 94.6000 51.1000 95.0000 52.1000 ;
	    RECT 96.6000 51.8000 97.3000 52.1000 ;
	    RECT 96.7000 51.1000 97.3000 51.8000 ;
	    RECT 99.0000 51.1000 99.4000 53.3000 ;
	    RECT 99.8000 51.1000 100.2000 59.9000 ;
	    RECT 102.2000 55.6000 102.6000 59.9000 ;
	    RECT 103.8000 55.6000 104.2000 59.9000 ;
	    RECT 105.4000 55.6000 105.8000 59.9000 ;
	    RECT 107.0000 55.6000 107.4000 59.9000 ;
	    RECT 108.6000 57.9000 109.0000 59.9000 ;
	    RECT 108.7000 57.8000 109.0000 57.9000 ;
	    RECT 110.2000 57.9000 110.6000 59.9000 ;
	    RECT 110.2000 57.8000 110.5000 57.9000 ;
	    RECT 108.7000 57.5000 110.5000 57.8000 ;
	    RECT 108.7000 56.2000 109.0000 57.5000 ;
	    RECT 109.4000 56.4000 109.8000 57.2000 ;
	    RECT 108.6000 55.8000 109.0000 56.2000 ;
	    RECT 101.4000 55.2000 102.6000 55.6000 ;
	    RECT 103.1000 55.2000 104.2000 55.6000 ;
	    RECT 104.7000 55.2000 105.8000 55.6000 ;
	    RECT 106.5000 55.2000 107.4000 55.6000 ;
	    RECT 101.4000 53.8000 101.8000 55.2000 ;
	    RECT 103.1000 54.5000 103.5000 55.2000 ;
	    RECT 104.7000 54.5000 105.1000 55.2000 ;
	    RECT 106.5000 54.5000 106.9000 55.2000 ;
	    RECT 102.2000 54.1000 103.5000 54.5000 ;
	    RECT 103.9000 54.1000 105.1000 54.5000 ;
	    RECT 105.6000 54.1000 106.9000 54.5000 ;
	    RECT 103.1000 53.8000 103.5000 54.1000 ;
	    RECT 104.7000 53.8000 105.1000 54.1000 ;
	    RECT 106.5000 53.8000 106.9000 54.1000 ;
	    RECT 108.7000 54.2000 109.0000 55.8000 ;
	    RECT 113.4000 55.9000 113.8000 59.9000 ;
	    RECT 115.0000 56.2000 115.4000 59.9000 ;
	    RECT 116.6000 57.9000 117.0000 59.9000 ;
	    RECT 116.7000 57.8000 117.0000 57.9000 ;
	    RECT 118.2000 57.9000 118.6000 59.9000 ;
	    RECT 118.2000 57.8000 118.5000 57.9000 ;
	    RECT 116.7000 57.5000 118.5000 57.8000 ;
	    RECT 117.4000 56.4000 117.8000 57.2000 ;
	    RECT 114.3000 55.9000 115.4000 56.2000 ;
	    RECT 118.2000 56.2000 118.5000 57.5000 ;
	    RECT 109.4000 54.8000 110.6000 55.2000 ;
	    RECT 113.4000 54.8000 113.7000 55.9000 ;
	    RECT 114.3000 55.6000 114.6000 55.9000 ;
	    RECT 114.0000 55.2000 114.6000 55.6000 ;
	    RECT 118.2000 55.8000 118.6000 56.2000 ;
	    RECT 119.8000 56.1000 120.2000 59.9000 ;
	    RECT 120.6000 56.1000 121.0000 56.6000 ;
	    RECT 119.8000 55.8000 121.0000 56.1000 ;
	    RECT 108.7000 54.1000 109.5000 54.2000 ;
	    RECT 112.6000 54.1000 113.0000 54.2000 ;
	    RECT 113.4000 54.1000 113.8000 54.8000 ;
	    RECT 108.7000 53.9000 109.6000 54.1000 ;
	    RECT 101.4000 53.4000 102.6000 53.8000 ;
	    RECT 103.1000 53.4000 104.2000 53.8000 ;
	    RECT 104.7000 53.4000 105.8000 53.8000 ;
	    RECT 106.5000 53.4000 107.4000 53.8000 ;
	    RECT 102.2000 51.1000 102.6000 53.4000 ;
	    RECT 103.8000 51.1000 104.2000 53.4000 ;
	    RECT 105.4000 51.1000 105.8000 53.4000 ;
	    RECT 107.0000 51.1000 107.4000 53.4000 ;
	    RECT 109.2000 51.1000 109.6000 53.9000 ;
	    RECT 112.6000 53.8000 113.8000 54.1000 ;
	    RECT 113.4000 51.1000 113.8000 53.8000 ;
	    RECT 114.3000 53.7000 114.6000 55.2000 ;
	    RECT 116.6000 54.8000 117.4000 55.2000 ;
	    RECT 118.2000 54.2000 118.5000 55.8000 ;
	    RECT 117.7000 54.1000 118.5000 54.2000 ;
	    RECT 117.6000 53.9000 118.5000 54.1000 ;
	    RECT 114.3000 53.4000 115.4000 53.7000 ;
	    RECT 115.0000 51.1000 115.4000 53.4000 ;
	    RECT 117.6000 51.1000 118.0000 53.9000 ;
	    RECT 119.8000 51.1000 120.2000 55.8000 ;
	    RECT 121.4000 53.1000 121.8000 59.9000 ;
	    RECT 123.0000 56.2000 123.4000 59.9000 ;
	    RECT 123.0000 55.9000 124.1000 56.2000 ;
	    RECT 124.6000 55.9000 125.0000 59.9000 ;
	    RECT 123.8000 55.6000 124.1000 55.9000 ;
	    RECT 123.8000 55.2000 124.4000 55.6000 ;
	    RECT 122.2000 53.4000 122.6000 54.2000 ;
	    RECT 123.8000 53.7000 124.1000 55.2000 ;
	    RECT 124.7000 54.8000 125.0000 55.9000 ;
	    RECT 123.0000 53.4000 124.1000 53.7000 ;
	    RECT 124.6000 54.1000 125.0000 54.8000 ;
	    RECT 125.4000 54.1000 125.8000 54.2000 ;
	    RECT 124.6000 53.8000 125.8000 54.1000 ;
	    RECT 120.9000 52.8000 121.8000 53.1000 ;
	    RECT 120.9000 52.2000 121.3000 52.8000 ;
	    RECT 120.6000 51.8000 121.3000 52.2000 ;
	    RECT 120.9000 51.1000 121.3000 51.8000 ;
	    RECT 123.0000 51.1000 123.4000 53.4000 ;
	    RECT 124.6000 51.1000 125.0000 53.8000 ;
	    RECT 125.4000 53.4000 125.8000 53.8000 ;
	    RECT 126.2000 53.1000 126.6000 59.9000 ;
	    RECT 127.0000 56.1000 127.4000 56.6000 ;
	    RECT 127.8000 56.1000 128.2000 59.9000 ;
	    RECT 127.0000 55.8000 128.2000 56.1000 ;
	    RECT 126.2000 52.8000 127.1000 53.1000 ;
	    RECT 126.7000 52.2000 127.1000 52.8000 ;
	    RECT 126.7000 51.8000 127.4000 52.2000 ;
	    RECT 126.7000 51.1000 127.1000 51.8000 ;
	    RECT 127.8000 51.1000 128.2000 55.8000 ;
	    RECT 129.4000 53.4000 129.8000 54.2000 ;
	    RECT 130.2000 53.1000 130.6000 59.9000 ;
	    RECT 131.0000 56.1000 131.4000 56.6000 ;
	    RECT 131.8000 56.1000 132.2000 59.9000 ;
	    RECT 131.0000 55.8000 132.2000 56.1000 ;
	    RECT 130.2000 52.8000 131.1000 53.1000 ;
	    RECT 130.7000 52.2000 131.1000 52.8000 ;
	    RECT 130.7000 51.8000 131.4000 52.2000 ;
	    RECT 130.7000 51.1000 131.1000 51.8000 ;
	    RECT 131.8000 51.1000 132.2000 55.8000 ;
	    RECT 133.4000 51.1000 133.8000 59.9000 ;
	    RECT 135.8000 57.9000 136.2000 59.9000 ;
	    RECT 135.9000 57.8000 136.2000 57.9000 ;
	    RECT 137.4000 57.9000 137.8000 59.9000 ;
	    RECT 137.4000 57.8000 137.7000 57.9000 ;
	    RECT 135.9000 57.5000 137.7000 57.8000 ;
	    RECT 136.6000 56.4000 137.0000 57.2000 ;
	    RECT 137.4000 56.2000 137.7000 57.5000 ;
	    RECT 137.4000 55.8000 137.8000 56.2000 ;
	    RECT 135.8000 54.8000 136.6000 55.2000 ;
	    RECT 137.4000 54.2000 137.7000 55.8000 ;
	    RECT 138.2000 55.6000 138.6000 59.9000 ;
	    RECT 140.3000 56.2000 140.7000 59.9000 ;
	    RECT 142.2000 57.8000 142.6000 59.9000 ;
	    RECT 143.8000 57.9000 144.2000 59.9000 ;
	    RECT 143.8000 57.8000 144.1000 57.9000 ;
	    RECT 142.2000 57.5000 144.1000 57.8000 ;
	    RECT 142.2000 57.2000 142.5000 57.5000 ;
	    RECT 142.2000 56.8000 142.6000 57.2000 ;
	    RECT 143.0000 56.4000 143.4000 57.2000 ;
	    RECT 143.8000 56.2000 144.1000 57.5000 ;
	    RECT 145.4000 57.8000 145.8000 59.9000 ;
	    RECT 147.0000 57.9000 147.4000 59.9000 ;
	    RECT 147.0000 57.8000 147.3000 57.9000 ;
	    RECT 145.4000 57.5000 147.3000 57.8000 ;
	    RECT 145.4000 57.2000 145.7000 57.5000 ;
	    RECT 145.4000 56.8000 145.8000 57.2000 ;
	    RECT 146.2000 56.4000 146.6000 57.2000 ;
	    RECT 147.0000 56.2000 147.3000 57.5000 ;
	    RECT 140.3000 55.9000 141.0000 56.2000 ;
	    RECT 138.2000 55.4000 140.2000 55.6000 ;
	    RECT 138.2000 55.3000 140.3000 55.4000 ;
	    RECT 139.9000 55.0000 140.3000 55.3000 ;
	    RECT 140.7000 55.2000 141.0000 55.9000 ;
	    RECT 141.4000 56.1000 141.8000 56.2000 ;
	    RECT 142.2000 56.1000 142.6000 56.2000 ;
	    RECT 141.4000 55.8000 142.6000 56.1000 ;
	    RECT 143.8000 55.8000 144.2000 56.2000 ;
	    RECT 147.0000 55.8000 147.4000 56.2000 ;
	    RECT 141.4000 55.4000 141.8000 55.8000 ;
	    RECT 136.9000 54.1000 137.7000 54.2000 ;
	    RECT 136.8000 53.9000 137.7000 54.1000 ;
	    RECT 136.8000 51.1000 137.2000 53.9000 ;
	    RECT 140.0000 53.5000 140.3000 55.0000 ;
	    RECT 140.6000 54.8000 141.0000 55.2000 ;
	    RECT 142.2000 54.8000 143.0000 55.2000 ;
	    RECT 139.1000 53.2000 140.3000 53.5000 ;
	    RECT 138.2000 52.4000 138.6000 53.2000 ;
	    RECT 139.1000 52.1000 139.4000 53.2000 ;
	    RECT 140.7000 53.1000 141.0000 54.8000 ;
	    RECT 143.8000 54.2000 144.1000 55.8000 ;
	    RECT 145.4000 54.8000 146.2000 55.2000 ;
	    RECT 147.0000 54.2000 147.3000 55.8000 ;
	    RECT 143.3000 54.1000 144.1000 54.2000 ;
	    RECT 146.5000 54.1000 147.3000 54.2000 ;
	    RECT 139.0000 51.1000 139.4000 52.1000 ;
	    RECT 140.6000 51.1000 141.0000 53.1000 ;
	    RECT 143.2000 53.9000 144.1000 54.1000 ;
	    RECT 146.4000 53.9000 147.3000 54.1000 ;
	    RECT 143.2000 51.1000 143.6000 53.9000 ;
	    RECT 146.4000 51.1000 146.8000 53.9000 ;
	    RECT 147.8000 53.4000 148.2000 54.2000 ;
	    RECT 148.6000 53.1000 149.0000 59.9000 ;
	    RECT 149.4000 56.1000 149.8000 56.6000 ;
	    RECT 150.2000 56.1000 150.6000 59.9000 ;
	    RECT 149.4000 55.8000 150.6000 56.1000 ;
	    RECT 148.6000 52.8000 149.5000 53.1000 ;
	    RECT 149.1000 51.1000 149.5000 52.8000 ;
	    RECT 150.2000 51.1000 150.6000 55.8000 ;
	    RECT 152.6000 53.1000 153.0000 59.9000 ;
	    RECT 153.4000 56.1000 153.8000 56.6000 ;
	    RECT 154.2000 56.1000 154.6000 56.2000 ;
	    RECT 153.4000 55.8000 154.6000 56.1000 ;
	    RECT 154.2000 53.4000 154.6000 54.2000 ;
	    RECT 155.0000 53.1000 155.4000 59.9000 ;
	    RECT 155.8000 56.1000 156.2000 56.6000 ;
	    RECT 157.4000 56.1000 157.8000 59.9000 ;
	    RECT 155.8000 55.8000 157.8000 56.1000 ;
	    RECT 152.6000 52.8000 153.5000 53.1000 ;
	    RECT 155.0000 52.8000 155.9000 53.1000 ;
	    RECT 153.1000 52.2000 153.5000 52.8000 ;
	    RECT 152.6000 51.8000 153.5000 52.2000 ;
	    RECT 153.1000 51.1000 153.5000 51.8000 ;
	    RECT 155.5000 52.2000 155.9000 52.8000 ;
	    RECT 155.5000 51.8000 156.2000 52.2000 ;
	    RECT 155.5000 51.1000 155.9000 51.8000 ;
	    RECT 157.4000 51.1000 157.8000 55.8000 ;
	    RECT 159.0000 54.1000 159.4000 59.9000 ;
	    RECT 161.1000 56.2000 161.5000 59.9000 ;
	    RECT 163.8000 57.9000 164.2000 59.9000 ;
	    RECT 161.8000 56.8000 162.2000 57.2000 ;
	    RECT 161.9000 56.2000 162.2000 56.8000 ;
	    RECT 160.6000 55.8000 161.6000 56.2000 ;
	    RECT 161.9000 55.9000 162.6000 56.2000 ;
	    RECT 162.2000 55.8000 162.6000 55.9000 ;
	    RECT 163.9000 55.8000 164.2000 57.9000 ;
	    RECT 165.4000 55.9000 165.8000 59.9000 ;
	    RECT 159.8000 55.1000 160.2000 55.2000 ;
	    RECT 160.6000 55.1000 161.0000 55.2000 ;
	    RECT 159.8000 54.8000 161.0000 55.1000 ;
	    RECT 160.6000 54.4000 161.0000 54.8000 ;
	    RECT 161.3000 54.2000 161.6000 55.8000 ;
	    RECT 163.9000 55.5000 165.1000 55.8000 ;
	    RECT 163.8000 54.8000 164.2000 55.2000 ;
	    RECT 159.8000 54.1000 160.2000 54.2000 ;
	    RECT 159.0000 53.8000 160.6000 54.1000 ;
	    RECT 161.3000 53.8000 162.6000 54.2000 ;
	    RECT 163.0000 53.8000 163.4000 54.6000 ;
	    RECT 163.9000 54.4000 164.2000 54.8000 ;
	    RECT 163.9000 54.1000 164.4000 54.4000 ;
	    RECT 164.0000 54.0000 164.4000 54.1000 ;
	    RECT 164.8000 53.8000 165.1000 55.5000 ;
	    RECT 165.5000 55.2000 165.8000 55.9000 ;
	    RECT 165.4000 54.8000 165.8000 55.2000 ;
	    RECT 159.0000 51.1000 159.4000 53.8000 ;
	    RECT 160.2000 53.6000 160.6000 53.8000 ;
	    RECT 159.9000 53.1000 161.7000 53.3000 ;
	    RECT 162.2000 53.1000 162.5000 53.8000 ;
	    RECT 164.8000 53.7000 165.2000 53.8000 ;
	    RECT 163.7000 53.5000 165.2000 53.7000 ;
	    RECT 163.1000 53.4000 165.2000 53.5000 ;
	    RECT 163.1000 53.2000 164.0000 53.4000 ;
	    RECT 163.1000 53.1000 163.4000 53.2000 ;
	    RECT 165.5000 53.1000 165.8000 54.8000 ;
	    RECT 159.8000 53.0000 161.8000 53.1000 ;
	    RECT 159.8000 51.1000 160.2000 53.0000 ;
	    RECT 161.4000 51.1000 161.8000 53.0000 ;
	    RECT 162.2000 51.1000 162.6000 53.1000 ;
	    RECT 163.0000 51.1000 163.4000 53.1000 ;
	    RECT 165.1000 52.6000 165.8000 53.1000 ;
	    RECT 167.0000 56.1000 167.4000 59.9000 ;
	    RECT 167.8000 56.1000 168.2000 56.6000 ;
	    RECT 167.0000 55.8000 168.2000 56.1000 ;
	    RECT 165.1000 51.1000 165.5000 52.6000 ;
	    RECT 167.0000 51.1000 167.4000 55.8000 ;
	    RECT 168.6000 53.1000 169.0000 59.9000 ;
	    RECT 170.2000 56.2000 170.6000 59.9000 ;
	    RECT 170.2000 55.9000 171.3000 56.2000 ;
	    RECT 171.0000 55.6000 171.3000 55.9000 ;
	    RECT 171.0000 55.2000 171.6000 55.6000 ;
	    RECT 170.2000 54.4000 170.6000 55.2000 ;
	    RECT 169.4000 53.4000 169.8000 54.2000 ;
	    RECT 171.0000 53.7000 171.3000 55.2000 ;
	    RECT 170.2000 53.4000 171.3000 53.7000 ;
	    RECT 168.1000 52.8000 169.0000 53.1000 ;
	    RECT 168.1000 52.2000 168.5000 52.8000 ;
	    RECT 167.8000 51.8000 168.5000 52.2000 ;
	    RECT 168.1000 51.1000 168.5000 51.8000 ;
	    RECT 170.2000 51.1000 170.6000 53.4000 ;
	    RECT 1.4000 49.1000 1.8000 49.2000 ;
	    RECT 2.4000 49.1000 2.8000 49.9000 ;
	    RECT 1.4000 48.8000 2.8000 49.1000 ;
	    RECT 2.4000 47.1000 2.8000 48.8000 ;
	    RECT 3.8000 47.9000 4.2000 49.9000 ;
	    RECT 5.4000 48.9000 5.8000 49.9000 ;
	    RECT 2.4000 46.9000 3.3000 47.1000 ;
	    RECT 2.5000 46.8000 3.3000 46.9000 ;
	    RECT 1.4000 45.8000 2.2000 46.2000 ;
	    RECT 3.0000 45.2000 3.3000 46.8000 ;
	    RECT 3.8000 46.2000 4.1000 47.9000 ;
	    RECT 5.4000 47.8000 5.7000 48.9000 ;
	    RECT 6.2000 47.8000 6.6000 48.6000 ;
	    RECT 4.5000 47.5000 5.7000 47.8000 ;
	    RECT 3.8000 45.8000 4.2000 46.2000 ;
	    RECT 4.5000 46.0000 4.8000 47.5000 ;
	    RECT 3.0000 44.8000 3.4000 45.2000 ;
	    RECT 3.8000 45.1000 4.1000 45.8000 ;
	    RECT 4.5000 45.7000 4.9000 46.0000 ;
	    RECT 4.5000 45.6000 6.6000 45.7000 ;
	    RECT 4.6000 45.4000 6.6000 45.6000 ;
	    RECT 3.8000 44.8000 4.5000 45.1000 ;
	    RECT 2.2000 43.8000 2.6000 44.6000 ;
	    RECT 3.0000 43.5000 3.3000 44.8000 ;
	    RECT 1.5000 43.2000 3.3000 43.5000 ;
	    RECT 1.5000 43.1000 1.8000 43.2000 ;
	    RECT 1.4000 41.1000 1.8000 43.1000 ;
	    RECT 3.0000 43.1000 3.3000 43.2000 ;
	    RECT 3.0000 41.1000 3.4000 43.1000 ;
	    RECT 4.1000 41.1000 4.5000 44.8000 ;
	    RECT 6.2000 41.1000 6.6000 45.4000 ;
	    RECT 7.0000 45.1000 7.4000 49.9000 ;
	    RECT 8.9000 48.2000 9.3000 49.9000 ;
	    RECT 12.3000 49.2000 12.7000 49.9000 ;
	    RECT 11.8000 48.8000 12.7000 49.2000 ;
	    RECT 12.3000 48.2000 12.7000 48.8000 ;
	    RECT 8.9000 47.9000 9.8000 48.2000 ;
	    RECT 7.8000 46.1000 8.2000 46.2000 ;
	    RECT 9.4000 46.1000 9.8000 47.9000 ;
	    RECT 11.8000 47.9000 12.7000 48.2000 ;
	    RECT 10.2000 46.8000 10.6000 47.6000 ;
	    RECT 7.8000 45.8000 9.8000 46.1000 ;
	    RECT 8.6000 45.1000 9.0000 45.2000 ;
	    RECT 7.0000 44.8000 9.0000 45.1000 ;
	    RECT 7.0000 41.1000 7.4000 44.8000 ;
	    RECT 8.6000 44.4000 9.0000 44.8000 ;
	    RECT 9.4000 41.1000 9.8000 45.8000 ;
	    RECT 11.8000 41.1000 12.2000 47.9000 ;
	    RECT 12.6000 44.4000 13.0000 45.2000 ;
	    RECT 14.2000 45.1000 14.6000 49.9000 ;
	    RECT 16.3000 49.2000 16.7000 49.9000 ;
	    RECT 16.3000 48.8000 17.0000 49.2000 ;
	    RECT 16.3000 48.2000 16.7000 48.8000 ;
	    RECT 15.8000 47.9000 16.7000 48.2000 ;
	    RECT 15.0000 46.8000 15.4000 47.6000 ;
	    RECT 14.2000 44.8000 15.3000 45.1000 ;
	    RECT 14.2000 41.1000 14.6000 44.8000 ;
	    RECT 15.0000 44.2000 15.3000 44.8000 ;
	    RECT 15.0000 43.8000 15.4000 44.2000 ;
	    RECT 15.8000 41.1000 16.2000 47.9000 ;
	    RECT 19.2000 47.1000 19.6000 49.9000 ;
	    RECT 20.6000 47.9000 21.0000 49.9000 ;
	    RECT 22.2000 48.9000 22.6000 49.9000 ;
	    RECT 25.6000 49.2000 26.0000 49.9000 ;
	    RECT 19.2000 46.9000 20.1000 47.1000 ;
	    RECT 19.3000 46.8000 20.1000 46.9000 ;
	    RECT 18.2000 45.8000 19.0000 46.2000 ;
	    RECT 19.8000 45.2000 20.1000 46.8000 ;
	    RECT 20.6000 46.2000 20.9000 47.9000 ;
	    RECT 22.2000 47.8000 22.5000 48.9000 ;
	    RECT 25.6000 48.8000 26.6000 49.2000 ;
	    RECT 23.0000 47.8000 23.4000 48.6000 ;
	    RECT 21.3000 47.5000 22.5000 47.8000 ;
	    RECT 20.6000 45.8000 21.0000 46.2000 ;
	    RECT 21.3000 46.0000 21.6000 47.5000 ;
	    RECT 25.6000 47.1000 26.0000 48.8000 ;
	    RECT 28.3000 48.2000 28.7000 49.9000 ;
	    RECT 27.8000 47.9000 28.7000 48.2000 ;
	    RECT 25.6000 46.9000 26.5000 47.1000 ;
	    RECT 25.7000 46.8000 26.5000 46.9000 ;
	    RECT 27.0000 46.8000 27.4000 47.6000 ;
	    RECT 16.6000 44.4000 17.0000 45.2000 ;
	    RECT 19.8000 44.8000 20.2000 45.2000 ;
	    RECT 20.6000 45.1000 20.9000 45.8000 ;
	    RECT 21.3000 45.7000 21.7000 46.0000 ;
	    RECT 24.6000 45.8000 25.4000 46.2000 ;
	    RECT 21.3000 45.6000 23.4000 45.7000 ;
	    RECT 21.4000 45.4000 23.4000 45.6000 ;
	    RECT 20.6000 44.8000 21.3000 45.1000 ;
	    RECT 19.0000 43.8000 19.4000 44.6000 ;
	    RECT 19.8000 43.5000 20.1000 44.8000 ;
	    RECT 18.3000 43.2000 20.1000 43.5000 ;
	    RECT 18.3000 43.1000 18.6000 43.2000 ;
	    RECT 18.2000 41.1000 18.6000 43.1000 ;
	    RECT 19.8000 43.1000 20.1000 43.2000 ;
	    RECT 19.8000 41.1000 20.2000 43.1000 ;
	    RECT 20.9000 41.1000 21.3000 44.8000 ;
	    RECT 23.0000 41.1000 23.4000 45.4000 ;
	    RECT 26.2000 45.2000 26.5000 46.8000 ;
	    RECT 26.2000 44.8000 26.6000 45.2000 ;
	    RECT 25.4000 43.8000 25.8000 44.6000 ;
	    RECT 26.2000 43.5000 26.5000 44.8000 ;
	    RECT 24.7000 43.2000 26.5000 43.5000 ;
	    RECT 24.7000 43.1000 25.0000 43.2000 ;
	    RECT 24.6000 41.1000 25.0000 43.1000 ;
	    RECT 26.2000 43.1000 26.5000 43.2000 ;
	    RECT 26.2000 41.1000 26.6000 43.1000 ;
	    RECT 27.8000 41.1000 28.2000 47.9000 ;
	    RECT 31.2000 47.1000 31.6000 49.9000 ;
	    RECT 34.4000 47.1000 34.8000 49.9000 ;
	    RECT 35.8000 47.9000 36.2000 49.9000 ;
	    RECT 37.4000 48.9000 37.8000 49.9000 ;
	    RECT 31.2000 46.9000 32.1000 47.1000 ;
	    RECT 34.4000 46.9000 35.3000 47.1000 ;
	    RECT 31.3000 46.8000 32.1000 46.9000 ;
	    RECT 34.5000 46.8000 35.3000 46.9000 ;
	    RECT 30.2000 45.8000 31.0000 46.2000 ;
	    RECT 31.8000 45.2000 32.1000 46.8000 ;
	    RECT 33.4000 45.8000 34.6000 46.2000 ;
	    RECT 35.0000 45.2000 35.3000 46.8000 ;
	    RECT 35.8000 46.2000 36.1000 47.9000 ;
	    RECT 37.4000 47.8000 37.7000 48.9000 ;
	    RECT 38.2000 47.8000 38.6000 48.6000 ;
	    RECT 40.3000 48.2000 40.7000 49.9000 ;
	    RECT 42.7000 48.2000 43.1000 49.9000 ;
	    RECT 45.1000 48.2000 45.5000 49.9000 ;
	    RECT 39.8000 47.9000 40.7000 48.2000 ;
	    RECT 42.2000 47.9000 43.1000 48.2000 ;
	    RECT 44.6000 47.9000 45.5000 48.2000 ;
	    RECT 36.5000 47.5000 37.7000 47.8000 ;
	    RECT 35.8000 45.8000 36.2000 46.2000 ;
	    RECT 36.5000 46.0000 36.8000 47.5000 ;
	    RECT 38.2000 47.1000 38.6000 47.2000 ;
	    RECT 39.0000 47.1000 39.4000 47.6000 ;
	    RECT 38.2000 46.8000 39.4000 47.1000 ;
	    RECT 28.6000 44.4000 29.0000 45.2000 ;
	    RECT 31.8000 44.8000 32.2000 45.2000 ;
	    RECT 35.0000 44.8000 35.4000 45.2000 ;
	    RECT 35.8000 45.1000 36.1000 45.8000 ;
	    RECT 36.5000 45.7000 36.9000 46.0000 ;
	    RECT 36.5000 45.6000 38.6000 45.7000 ;
	    RECT 36.6000 45.4000 38.6000 45.6000 ;
	    RECT 35.8000 44.8000 36.5000 45.1000 ;
	    RECT 31.0000 43.8000 31.4000 44.6000 ;
	    RECT 31.8000 43.5000 32.1000 44.8000 ;
	    RECT 34.2000 43.8000 34.6000 44.6000 ;
	    RECT 35.0000 43.5000 35.3000 44.8000 ;
	    RECT 30.3000 43.2000 32.1000 43.5000 ;
	    RECT 33.5000 43.2000 35.3000 43.5000 ;
	    RECT 30.3000 43.1000 30.6000 43.2000 ;
	    RECT 30.2000 41.1000 30.6000 43.1000 ;
	    RECT 31.8000 43.1000 32.1000 43.2000 ;
	    RECT 31.8000 41.1000 32.2000 43.1000 ;
	    RECT 33.4000 41.1000 33.8000 43.2000 ;
	    RECT 35.0000 43.1000 35.3000 43.2000 ;
	    RECT 35.0000 41.1000 35.4000 43.1000 ;
	    RECT 36.1000 41.1000 36.5000 44.8000 ;
	    RECT 38.2000 41.1000 38.6000 45.4000 ;
	    RECT 39.8000 41.1000 40.2000 47.9000 ;
	    RECT 41.4000 46.8000 41.8000 47.6000 ;
	    RECT 40.6000 44.4000 41.0000 45.2000 ;
	    RECT 42.2000 41.1000 42.6000 47.9000 ;
	    RECT 43.8000 46.8000 44.2000 47.6000 ;
	    RECT 43.8000 44.1000 44.2000 44.2000 ;
	    RECT 44.6000 44.1000 45.0000 47.9000 ;
	    RECT 46.2000 47.1000 46.6000 49.9000 ;
	    RECT 45.4000 46.8000 46.6000 47.1000 ;
	    RECT 45.4000 46.2000 45.7000 46.8000 ;
	    RECT 45.4000 45.8000 45.8000 46.2000 ;
	    RECT 45.4000 44.4000 45.8000 45.2000 ;
	    RECT 43.8000 43.8000 45.0000 44.1000 ;
	    RECT 44.6000 41.1000 45.0000 43.8000 ;
	    RECT 46.2000 41.1000 46.6000 46.8000 ;
	    RECT 47.0000 45.8000 47.4000 46.2000 ;
	    RECT 47.0000 45.1000 47.3000 45.8000 ;
	    RECT 47.8000 45.1000 48.2000 49.9000 ;
	    RECT 47.0000 44.8000 48.2000 45.1000 ;
	    RECT 47.8000 41.1000 48.2000 44.8000 ;
	    RECT 50.2000 45.1000 50.6000 49.9000 ;
	    RECT 51.3000 48.2000 51.7000 49.9000 ;
	    RECT 54.2000 48.9000 54.6000 49.9000 ;
	    RECT 51.3000 47.9000 52.2000 48.2000 ;
	    RECT 51.0000 45.1000 51.4000 45.2000 ;
	    RECT 50.2000 44.8000 51.4000 45.1000 ;
	    RECT 50.2000 41.1000 50.6000 44.8000 ;
	    RECT 51.0000 44.4000 51.4000 44.8000 ;
	    RECT 51.8000 41.1000 52.2000 47.9000 ;
	    RECT 54.3000 47.8000 54.6000 48.9000 ;
	    RECT 55.8000 47.9000 56.2000 49.9000 ;
	    RECT 52.6000 47.1000 53.0000 47.6000 ;
	    RECT 54.3000 47.5000 55.5000 47.8000 ;
	    RECT 53.4000 47.1000 53.8000 47.2000 ;
	    RECT 54.2000 47.1000 54.7000 47.2000 ;
	    RECT 52.6000 46.8000 54.7000 47.1000 ;
	    RECT 54.4000 46.4000 54.8000 46.8000 ;
	    RECT 55.2000 46.0000 55.5000 47.5000 ;
	    RECT 55.9000 46.2000 56.2000 47.9000 ;
	    RECT 57.2000 47.1000 57.6000 49.9000 ;
	    RECT 62.2000 48.9000 62.6000 49.9000 ;
	    RECT 61.4000 47.8000 61.8000 48.6000 ;
	    RECT 62.3000 47.8000 62.6000 48.9000 ;
	    RECT 63.8000 47.9000 64.2000 49.9000 ;
	    RECT 62.3000 47.5000 63.5000 47.8000 ;
	    RECT 55.1000 45.7000 55.5000 46.0000 ;
	    RECT 55.8000 45.8000 56.2000 46.2000 ;
	    RECT 53.4000 45.6000 55.5000 45.7000 ;
	    RECT 53.4000 45.4000 55.4000 45.6000 ;
	    RECT 53.4000 41.1000 53.8000 45.4000 ;
	    RECT 55.9000 45.2000 56.2000 45.8000 ;
	    RECT 56.7000 46.9000 57.6000 47.1000 ;
	    RECT 56.7000 46.8000 57.5000 46.9000 ;
	    RECT 56.7000 45.2000 57.0000 46.8000 ;
	    RECT 57.8000 45.8000 58.6000 46.2000 ;
	    RECT 63.2000 46.0000 63.5000 47.5000 ;
	    RECT 63.9000 47.2000 64.2000 47.9000 ;
	    RECT 63.8000 46.8000 64.2000 47.2000 ;
	    RECT 65.2000 47.1000 65.6000 49.9000 ;
	    RECT 63.9000 46.2000 64.2000 46.8000 ;
	    RECT 63.1000 45.7000 63.5000 46.0000 ;
	    RECT 63.8000 45.8000 64.2000 46.2000 ;
	    RECT 61.4000 45.6000 63.5000 45.7000 ;
	    RECT 55.8000 45.1000 56.2000 45.2000 ;
	    RECT 55.5000 44.8000 56.2000 45.1000 ;
	    RECT 56.6000 44.8000 57.0000 45.2000 ;
	    RECT 59.0000 44.8000 59.4000 45.6000 ;
	    RECT 61.4000 45.4000 63.4000 45.6000 ;
	    RECT 55.5000 41.1000 55.9000 44.8000 ;
	    RECT 56.7000 43.5000 57.0000 44.8000 ;
	    RECT 57.4000 43.8000 57.8000 44.6000 ;
	    RECT 60.6000 44.1000 61.0000 44.2000 ;
	    RECT 58.2000 43.8000 61.0000 44.1000 ;
	    RECT 58.2000 43.5000 58.5000 43.8000 ;
	    RECT 56.7000 43.2000 58.5000 43.5000 ;
	    RECT 56.7000 43.1000 57.0000 43.2000 ;
	    RECT 56.6000 41.1000 57.0000 43.1000 ;
	    RECT 58.2000 43.1000 58.5000 43.2000 ;
	    RECT 58.2000 41.1000 58.6000 43.1000 ;
	    RECT 61.4000 41.1000 61.8000 45.4000 ;
	    RECT 63.9000 45.1000 64.2000 45.8000 ;
	    RECT 64.7000 46.9000 65.6000 47.1000 ;
	    RECT 69.6000 49.2000 70.0000 49.9000 ;
	    RECT 69.6000 48.8000 70.6000 49.2000 ;
	    RECT 69.6000 47.1000 70.0000 48.8000 ;
	    RECT 72.8000 47.1000 73.2000 49.9000 ;
	    RECT 74.2000 47.9000 74.6000 49.9000 ;
	    RECT 75.8000 48.9000 76.2000 49.9000 ;
	    RECT 74.2000 47.2000 74.5000 47.9000 ;
	    RECT 75.8000 47.8000 76.1000 48.9000 ;
	    RECT 74.9000 47.5000 76.1000 47.8000 ;
	    RECT 76.6000 47.8000 77.0000 48.6000 ;
	    RECT 78.7000 48.2000 79.1000 49.9000 ;
	    RECT 78.2000 47.9000 79.1000 48.2000 ;
	    RECT 69.6000 46.9000 70.5000 47.1000 ;
	    RECT 72.8000 46.9000 73.7000 47.1000 ;
	    RECT 64.7000 46.8000 65.5000 46.9000 ;
	    RECT 69.7000 46.8000 70.5000 46.9000 ;
	    RECT 72.9000 46.8000 73.7000 46.9000 ;
	    RECT 64.7000 45.2000 65.0000 46.8000 ;
	    RECT 65.8000 45.8000 66.6000 46.2000 ;
	    RECT 68.6000 45.8000 69.4000 46.2000 ;
	    RECT 63.5000 44.8000 64.2000 45.1000 ;
	    RECT 64.6000 44.8000 65.0000 45.2000 ;
	    RECT 67.0000 44.8000 67.4000 45.6000 ;
	    RECT 67.8000 45.1000 68.2000 45.6000 ;
	    RECT 70.2000 45.2000 70.5000 46.8000 ;
	    RECT 71.8000 45.8000 72.6000 46.2000 ;
	    RECT 73.4000 45.2000 73.7000 46.8000 ;
	    RECT 74.2000 46.8000 74.6000 47.2000 ;
	    RECT 74.2000 46.2000 74.5000 46.8000 ;
	    RECT 74.2000 45.8000 74.6000 46.2000 ;
	    RECT 74.9000 46.0000 75.2000 47.5000 ;
	    RECT 76.6000 47.1000 76.9000 47.8000 ;
	    RECT 77.4000 47.1000 77.8000 47.6000 ;
	    RECT 76.6000 46.8000 77.8000 47.1000 ;
	    RECT 68.6000 45.1000 69.0000 45.2000 ;
	    RECT 67.8000 44.8000 69.0000 45.1000 ;
	    RECT 70.2000 44.8000 70.6000 45.2000 ;
	    RECT 73.4000 44.8000 73.8000 45.2000 ;
	    RECT 74.2000 45.1000 74.5000 45.8000 ;
	    RECT 74.9000 45.7000 75.3000 46.0000 ;
	    RECT 74.9000 45.6000 77.0000 45.7000 ;
	    RECT 75.0000 45.4000 77.0000 45.6000 ;
	    RECT 74.2000 44.8000 74.9000 45.1000 ;
	    RECT 63.5000 41.1000 63.9000 44.8000 ;
	    RECT 64.7000 43.5000 65.0000 44.8000 ;
	    RECT 65.4000 43.8000 65.8000 44.6000 ;
	    RECT 69.4000 43.8000 69.8000 44.6000 ;
	    RECT 70.2000 43.5000 70.5000 44.8000 ;
	    RECT 72.6000 43.8000 73.0000 44.6000 ;
	    RECT 73.4000 43.5000 73.7000 44.8000 ;
	    RECT 64.7000 43.2000 66.5000 43.5000 ;
	    RECT 64.7000 43.1000 65.0000 43.2000 ;
	    RECT 64.6000 41.1000 65.0000 43.1000 ;
	    RECT 66.2000 43.1000 66.5000 43.2000 ;
	    RECT 68.7000 43.2000 70.5000 43.5000 ;
	    RECT 68.7000 43.1000 69.0000 43.2000 ;
	    RECT 66.2000 41.1000 66.6000 43.1000 ;
	    RECT 68.6000 41.1000 69.0000 43.1000 ;
	    RECT 70.2000 43.1000 70.5000 43.2000 ;
	    RECT 71.9000 43.2000 73.7000 43.5000 ;
	    RECT 71.9000 43.1000 72.2000 43.2000 ;
	    RECT 70.2000 41.1000 70.6000 43.1000 ;
	    RECT 71.8000 41.1000 72.2000 43.1000 ;
	    RECT 73.4000 43.1000 73.7000 43.2000 ;
	    RECT 73.4000 41.1000 73.8000 43.1000 ;
	    RECT 74.5000 41.1000 74.9000 44.8000 ;
	    RECT 76.6000 41.1000 77.0000 45.4000 ;
	    RECT 78.2000 41.1000 78.6000 47.9000 ;
	    RECT 79.0000 45.1000 79.4000 45.2000 ;
	    RECT 80.6000 45.1000 81.0000 49.9000 ;
	    RECT 81.7000 48.2000 82.1000 49.9000 ;
	    RECT 81.7000 47.9000 82.6000 48.2000 ;
	    RECT 79.0000 44.8000 81.0000 45.1000 ;
	    RECT 79.0000 44.4000 79.4000 44.8000 ;
	    RECT 80.6000 41.1000 81.0000 44.8000 ;
	    RECT 82.2000 41.1000 82.6000 47.9000 ;
	    RECT 83.0000 46.8000 83.4000 47.6000 ;
	    RECT 85.6000 47.1000 86.0000 49.9000 ;
	    RECT 87.0000 47.9000 87.4000 49.9000 ;
	    RECT 88.6000 48.9000 89.0000 49.9000 ;
	    RECT 85.6000 46.9000 86.5000 47.1000 ;
	    RECT 85.7000 46.8000 86.5000 46.9000 ;
	    RECT 84.6000 45.8000 85.8000 46.2000 ;
	    RECT 86.2000 45.2000 86.5000 46.8000 ;
	    RECT 87.0000 46.2000 87.3000 47.9000 ;
	    RECT 88.6000 47.8000 88.9000 48.9000 ;
	    RECT 89.4000 47.8000 89.8000 48.6000 ;
	    RECT 91.5000 48.2000 91.9000 49.9000 ;
	    RECT 91.0000 47.9000 91.9000 48.2000 ;
	    RECT 87.7000 47.5000 88.9000 47.8000 ;
	    RECT 87.0000 45.8000 87.4000 46.2000 ;
	    RECT 87.7000 46.0000 88.0000 47.5000 ;
	    RECT 89.4000 47.1000 89.8000 47.2000 ;
	    RECT 90.2000 47.1000 90.6000 47.6000 ;
	    RECT 89.4000 46.8000 90.6000 47.1000 ;
	    RECT 86.2000 44.8000 86.6000 45.2000 ;
	    RECT 87.0000 45.1000 87.3000 45.8000 ;
	    RECT 87.7000 45.7000 88.1000 46.0000 ;
	    RECT 87.7000 45.6000 89.8000 45.7000 ;
	    RECT 87.8000 45.4000 89.8000 45.6000 ;
	    RECT 87.0000 44.8000 87.7000 45.1000 ;
	    RECT 85.4000 43.8000 85.8000 44.6000 ;
	    RECT 86.2000 43.5000 86.5000 44.8000 ;
	    RECT 84.7000 43.2000 86.5000 43.5000 ;
	    RECT 84.6000 41.1000 85.0000 43.2000 ;
	    RECT 86.2000 43.1000 86.5000 43.2000 ;
	    RECT 86.2000 41.1000 86.6000 43.1000 ;
	    RECT 87.3000 41.1000 87.7000 44.8000 ;
	    RECT 89.4000 41.1000 89.8000 45.4000 ;
	    RECT 90.2000 44.8000 90.6000 45.2000 ;
	    RECT 90.2000 44.1000 90.5000 44.8000 ;
	    RECT 91.0000 44.1000 91.4000 47.9000 ;
	    RECT 92.6000 47.1000 93.0000 49.9000 ;
	    RECT 91.8000 46.8000 93.0000 47.1000 ;
	    RECT 91.8000 46.2000 92.1000 46.8000 ;
	    RECT 91.8000 45.8000 92.2000 46.2000 ;
	    RECT 91.8000 44.4000 92.2000 45.2000 ;
	    RECT 90.2000 43.8000 91.4000 44.1000 ;
	    RECT 91.0000 41.1000 91.4000 43.8000 ;
	    RECT 92.6000 41.1000 93.0000 46.8000 ;
	    RECT 93.4000 45.8000 93.8000 46.2000 ;
	    RECT 93.4000 45.1000 93.7000 45.8000 ;
	    RECT 94.2000 45.1000 94.6000 49.9000 ;
	    RECT 96.4000 47.1000 96.8000 49.9000 ;
	    RECT 95.9000 46.9000 96.8000 47.1000 ;
	    RECT 100.8000 49.2000 101.2000 49.9000 ;
	    RECT 100.8000 48.8000 101.8000 49.2000 ;
	    RECT 100.8000 47.1000 101.2000 48.8000 ;
	    RECT 102.5000 48.2000 102.9000 49.9000 ;
	    RECT 105.9000 48.2000 106.3000 49.9000 ;
	    RECT 102.5000 47.9000 103.4000 48.2000 ;
	    RECT 103.0000 47.1000 103.4000 47.9000 ;
	    RECT 105.4000 47.9000 106.3000 48.2000 ;
	    RECT 107.0000 47.9000 107.4000 49.9000 ;
	    RECT 107.8000 48.0000 108.2000 49.9000 ;
	    RECT 109.4000 48.0000 109.8000 49.9000 ;
	    RECT 107.8000 47.9000 109.8000 48.0000 ;
	    RECT 100.8000 46.9000 101.7000 47.1000 ;
	    RECT 95.9000 46.8000 96.7000 46.9000 ;
	    RECT 100.9000 46.8000 101.7000 46.9000 ;
	    RECT 95.9000 45.2000 96.2000 46.8000 ;
	    RECT 97.0000 45.8000 97.8000 46.2000 ;
	    RECT 99.8000 45.8000 100.6000 46.2000 ;
	    RECT 93.4000 44.8000 94.6000 45.1000 ;
	    RECT 95.8000 44.8000 96.2000 45.2000 ;
	    RECT 98.2000 44.8000 98.6000 45.6000 ;
	    RECT 101.4000 45.2000 101.7000 46.8000 ;
	    RECT 102.2000 46.8000 103.4000 47.1000 ;
	    RECT 104.6000 46.8000 105.0000 47.6000 ;
	    RECT 102.2000 46.2000 102.5000 46.8000 ;
	    RECT 102.2000 45.8000 102.6000 46.2000 ;
	    RECT 101.4000 44.8000 101.8000 45.2000 ;
	    RECT 94.2000 41.1000 94.6000 44.8000 ;
	    RECT 95.9000 43.5000 96.2000 44.8000 ;
	    RECT 96.6000 43.8000 97.0000 44.6000 ;
	    RECT 100.6000 44.1000 101.0000 44.6000 ;
	    RECT 97.4000 43.8000 101.0000 44.1000 ;
	    RECT 97.4000 43.5000 97.7000 43.8000 ;
	    RECT 101.4000 43.5000 101.7000 44.8000 ;
	    RECT 102.2000 44.4000 102.6000 45.2000 ;
	    RECT 95.9000 43.2000 97.7000 43.5000 ;
	    RECT 95.9000 43.1000 96.2000 43.2000 ;
	    RECT 95.8000 41.1000 96.2000 43.1000 ;
	    RECT 97.4000 43.1000 97.7000 43.2000 ;
	    RECT 99.9000 43.2000 101.7000 43.5000 ;
	    RECT 99.9000 43.1000 100.2000 43.2000 ;
	    RECT 97.4000 41.1000 97.8000 43.1000 ;
	    RECT 99.8000 41.1000 100.2000 43.1000 ;
	    RECT 101.4000 43.1000 101.7000 43.2000 ;
	    RECT 101.4000 41.1000 101.8000 43.1000 ;
	    RECT 103.0000 41.1000 103.4000 46.8000 ;
	    RECT 105.4000 46.1000 105.8000 47.9000 ;
	    RECT 107.1000 47.2000 107.4000 47.9000 ;
	    RECT 107.9000 47.7000 109.7000 47.9000 ;
	    RECT 109.0000 47.2000 109.4000 47.4000 ;
	    RECT 107.0000 46.8000 108.3000 47.2000 ;
	    RECT 109.0000 47.1000 109.8000 47.2000 ;
	    RECT 110.2000 47.1000 110.6000 49.9000 ;
	    RECT 109.0000 46.9000 110.6000 47.1000 ;
	    RECT 109.4000 46.8000 110.6000 46.9000 ;
	    RECT 105.4000 45.8000 107.3000 46.1000 ;
	    RECT 105.4000 41.1000 105.8000 45.8000 ;
	    RECT 107.0000 45.2000 107.3000 45.8000 ;
	    RECT 107.0000 45.1000 107.4000 45.2000 ;
	    RECT 108.0000 45.1000 108.3000 46.8000 ;
	    RECT 108.6000 45.8000 109.0000 46.6000 ;
	    RECT 107.0000 44.8000 107.7000 45.1000 ;
	    RECT 108.0000 44.8000 108.5000 45.1000 ;
	    RECT 107.4000 44.2000 107.7000 44.8000 ;
	    RECT 108.1000 44.2000 108.5000 44.8000 ;
	    RECT 107.4000 43.8000 107.8000 44.2000 ;
	    RECT 108.1000 43.8000 109.0000 44.2000 ;
	    RECT 108.1000 41.1000 108.5000 43.8000 ;
	    RECT 110.2000 41.1000 110.6000 46.8000 ;
	    RECT 114.2000 41.1000 114.6000 49.9000 ;
	    RECT 117.6000 47.1000 118.0000 49.9000 ;
	    RECT 119.0000 47.9000 119.4000 49.9000 ;
	    RECT 120.6000 48.9000 121.0000 49.9000 ;
	    RECT 123.0000 49.1000 123.4000 49.2000 ;
	    RECT 124.0000 49.1000 124.4000 49.9000 ;
	    RECT 117.6000 46.9000 118.5000 47.1000 ;
	    RECT 117.7000 46.8000 118.5000 46.9000 ;
	    RECT 116.6000 45.8000 117.4000 46.2000 ;
	    RECT 118.2000 45.2000 118.5000 46.8000 ;
	    RECT 119.0000 46.2000 119.3000 47.9000 ;
	    RECT 120.6000 47.8000 120.9000 48.9000 ;
	    RECT 123.0000 48.8000 124.4000 49.1000 ;
	    RECT 121.4000 47.8000 121.8000 48.6000 ;
	    RECT 119.7000 47.5000 120.9000 47.8000 ;
	    RECT 119.0000 45.8000 119.4000 46.2000 ;
	    RECT 119.7000 46.0000 120.0000 47.5000 ;
	    RECT 124.0000 47.1000 124.4000 48.8000 ;
	    RECT 127.2000 47.1000 127.6000 49.9000 ;
	    RECT 130.4000 47.1000 130.8000 49.9000 ;
	    RECT 131.8000 47.9000 132.2000 49.9000 ;
	    RECT 133.4000 48.9000 133.8000 49.9000 ;
	    RECT 135.8000 48.9000 136.2000 49.9000 ;
	    RECT 124.0000 46.9000 124.9000 47.1000 ;
	    RECT 127.2000 46.9000 128.1000 47.1000 ;
	    RECT 130.4000 46.9000 131.3000 47.1000 ;
	    RECT 124.1000 46.8000 124.9000 46.9000 ;
	    RECT 127.3000 46.8000 128.1000 46.9000 ;
	    RECT 130.5000 46.8000 131.3000 46.9000 ;
	    RECT 118.2000 44.8000 118.6000 45.2000 ;
	    RECT 119.0000 45.1000 119.3000 45.8000 ;
	    RECT 119.7000 45.7000 120.1000 46.0000 ;
	    RECT 123.0000 45.8000 123.8000 46.2000 ;
	    RECT 119.7000 45.6000 121.8000 45.7000 ;
	    RECT 119.8000 45.4000 121.8000 45.6000 ;
	    RECT 119.0000 44.8000 119.7000 45.1000 ;
	    RECT 117.4000 43.8000 117.8000 44.6000 ;
	    RECT 118.2000 43.5000 118.5000 44.8000 ;
	    RECT 116.7000 43.2000 118.5000 43.5000 ;
	    RECT 116.7000 43.1000 117.0000 43.2000 ;
	    RECT 116.6000 41.1000 117.0000 43.1000 ;
	    RECT 118.2000 43.1000 118.5000 43.2000 ;
	    RECT 118.2000 41.1000 118.6000 43.1000 ;
	    RECT 119.3000 41.1000 119.7000 44.8000 ;
	    RECT 121.4000 41.1000 121.8000 45.4000 ;
	    RECT 124.6000 45.2000 124.9000 46.8000 ;
	    RECT 126.2000 45.8000 127.0000 46.2000 ;
	    RECT 127.8000 45.2000 128.1000 46.8000 ;
	    RECT 129.4000 45.8000 130.2000 46.2000 ;
	    RECT 124.6000 44.8000 125.0000 45.2000 ;
	    RECT 127.8000 44.8000 128.2000 45.2000 ;
	    RECT 128.6000 44.8000 129.0000 45.6000 ;
	    RECT 131.0000 45.2000 131.3000 46.8000 ;
	    RECT 131.8000 46.2000 132.1000 47.9000 ;
	    RECT 133.4000 47.8000 133.7000 48.9000 ;
	    RECT 134.2000 48.1000 134.6000 48.6000 ;
	    RECT 135.0000 48.1000 135.4000 48.6000 ;
	    RECT 134.2000 47.8000 135.4000 48.1000 ;
	    RECT 135.9000 47.8000 136.2000 48.9000 ;
	    RECT 137.4000 47.9000 137.8000 49.9000 ;
	    RECT 139.0000 48.9000 139.4000 49.9000 ;
	    RECT 132.5000 47.5000 133.7000 47.8000 ;
	    RECT 135.9000 47.5000 137.1000 47.8000 ;
	    RECT 131.8000 45.8000 132.2000 46.2000 ;
	    RECT 132.5000 46.0000 132.8000 47.5000 ;
	    RECT 136.8000 46.0000 137.1000 47.5000 ;
	    RECT 137.5000 46.2000 137.8000 47.9000 ;
	    RECT 139.1000 47.8000 139.4000 48.9000 ;
	    RECT 140.6000 47.9000 141.0000 49.9000 ;
	    RECT 142.2000 49.1000 142.6000 49.2000 ;
	    RECT 143.2000 49.1000 143.6000 49.9000 ;
	    RECT 142.2000 48.8000 143.6000 49.1000 ;
	    RECT 139.1000 47.5000 140.3000 47.8000 ;
	    RECT 139.0000 46.8000 139.5000 47.2000 ;
	    RECT 139.2000 46.4000 139.6000 46.8000 ;
	    RECT 131.8000 45.2000 132.1000 45.8000 ;
	    RECT 132.5000 45.7000 132.9000 46.0000 ;
	    RECT 136.7000 45.7000 137.1000 46.0000 ;
	    RECT 137.4000 45.8000 137.8000 46.2000 ;
	    RECT 140.0000 46.0000 140.3000 47.5000 ;
	    RECT 140.7000 47.2000 141.0000 47.9000 ;
	    RECT 140.6000 46.8000 141.0000 47.2000 ;
	    RECT 143.2000 47.1000 143.6000 48.8000 ;
	    RECT 144.9000 48.2000 145.3000 49.9000 ;
	    RECT 148.8000 49.2000 149.2000 49.9000 ;
	    RECT 148.6000 48.8000 149.2000 49.2000 ;
	    RECT 144.9000 47.9000 145.8000 48.2000 ;
	    RECT 143.2000 46.9000 144.1000 47.1000 ;
	    RECT 143.3000 46.8000 144.1000 46.9000 ;
	    RECT 140.7000 46.2000 141.0000 46.8000 ;
	    RECT 132.5000 45.6000 134.6000 45.7000 ;
	    RECT 132.6000 45.4000 134.6000 45.6000 ;
	    RECT 131.0000 44.8000 131.4000 45.2000 ;
	    RECT 131.8000 45.1000 132.2000 45.2000 ;
	    RECT 131.8000 44.8000 132.5000 45.1000 ;
	    RECT 123.8000 43.8000 124.2000 44.6000 ;
	    RECT 124.6000 43.5000 124.9000 44.8000 ;
	    RECT 127.0000 43.8000 127.4000 44.6000 ;
	    RECT 127.8000 43.5000 128.1000 44.8000 ;
	    RECT 130.2000 43.8000 130.6000 44.6000 ;
	    RECT 131.0000 43.5000 131.3000 44.8000 ;
	    RECT 123.1000 43.2000 124.9000 43.5000 ;
	    RECT 126.3000 43.2000 128.1000 43.5000 ;
	    RECT 123.1000 43.1000 123.4000 43.2000 ;
	    RECT 123.0000 41.1000 123.4000 43.1000 ;
	    RECT 124.6000 43.1000 124.9000 43.2000 ;
	    RECT 124.6000 41.1000 125.0000 43.1000 ;
	    RECT 126.2000 41.1000 126.6000 43.2000 ;
	    RECT 127.8000 43.1000 128.1000 43.2000 ;
	    RECT 129.5000 43.2000 131.3000 43.5000 ;
	    RECT 129.5000 43.1000 129.8000 43.2000 ;
	    RECT 127.8000 41.1000 128.2000 43.1000 ;
	    RECT 129.4000 41.1000 129.8000 43.1000 ;
	    RECT 131.0000 43.1000 131.3000 43.2000 ;
	    RECT 131.0000 41.1000 131.4000 43.1000 ;
	    RECT 132.1000 41.1000 132.5000 44.8000 ;
	    RECT 134.2000 41.1000 134.6000 45.4000 ;
	    RECT 135.0000 45.6000 137.1000 45.7000 ;
	    RECT 135.0000 45.4000 137.0000 45.6000 ;
	    RECT 135.0000 41.1000 135.4000 45.4000 ;
	    RECT 137.5000 45.1000 137.8000 45.8000 ;
	    RECT 139.9000 45.7000 140.3000 46.0000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 142.2000 45.8000 143.0000 46.2000 ;
	    RECT 137.1000 44.8000 137.8000 45.1000 ;
	    RECT 138.2000 45.6000 140.3000 45.7000 ;
	    RECT 138.2000 45.4000 140.2000 45.6000 ;
	    RECT 137.1000 41.1000 137.5000 44.8000 ;
	    RECT 138.2000 41.1000 138.6000 45.4000 ;
	    RECT 140.7000 45.1000 141.0000 45.8000 ;
	    RECT 140.3000 44.8000 141.0000 45.1000 ;
	    RECT 141.4000 44.8000 141.8000 45.6000 ;
	    RECT 143.8000 45.2000 144.1000 46.8000 ;
	    RECT 143.8000 44.8000 144.2000 45.2000 ;
	    RECT 140.3000 41.1000 140.7000 44.8000 ;
	    RECT 143.0000 43.8000 143.4000 44.6000 ;
	    RECT 143.8000 43.5000 144.1000 44.8000 ;
	    RECT 144.6000 44.4000 145.0000 45.2000 ;
	    RECT 142.3000 43.2000 144.1000 43.5000 ;
	    RECT 142.3000 43.1000 142.6000 43.2000 ;
	    RECT 142.2000 41.1000 142.6000 43.1000 ;
	    RECT 143.8000 43.1000 144.1000 43.2000 ;
	    RECT 143.8000 41.1000 144.2000 43.1000 ;
	    RECT 145.4000 41.1000 145.8000 47.9000 ;
	    RECT 146.2000 46.8000 146.6000 47.6000 ;
	    RECT 148.8000 47.1000 149.2000 48.8000 ;
	    RECT 152.0000 47.1000 152.4000 49.9000 ;
	    RECT 154.2000 48.9000 154.6000 49.9000 ;
	    RECT 153.4000 47.8000 153.8000 48.6000 ;
	    RECT 154.3000 47.8000 154.6000 48.9000 ;
	    RECT 155.8000 47.9000 156.2000 49.9000 ;
	    RECT 154.3000 47.5000 155.5000 47.8000 ;
	    RECT 148.8000 46.9000 149.7000 47.1000 ;
	    RECT 152.0000 46.9000 152.9000 47.1000 ;
	    RECT 148.9000 46.8000 149.7000 46.9000 ;
	    RECT 152.1000 46.8000 152.9000 46.9000 ;
	    RECT 147.8000 45.8000 148.6000 46.2000 ;
	    RECT 149.4000 45.2000 149.7000 46.8000 ;
	    RECT 151.0000 45.8000 151.8000 46.2000 ;
	    RECT 149.4000 44.8000 149.8000 45.2000 ;
	    RECT 150.2000 44.8000 150.6000 45.6000 ;
	    RECT 152.6000 45.2000 152.9000 46.8000 ;
	    RECT 155.2000 46.0000 155.5000 47.5000 ;
	    RECT 155.9000 46.2000 156.2000 47.9000 ;
	    RECT 157.2000 47.1000 157.6000 49.9000 ;
	    RECT 161.1000 49.2000 161.5000 49.9000 ;
	    RECT 161.1000 48.8000 161.8000 49.2000 ;
	    RECT 161.1000 48.2000 161.5000 48.8000 ;
	    RECT 158.2000 47.8000 158.6000 48.2000 ;
	    RECT 160.6000 47.9000 161.5000 48.2000 ;
	    RECT 158.2000 47.1000 158.5000 47.8000 ;
	    RECT 155.1000 45.7000 155.5000 46.0000 ;
	    RECT 155.8000 45.8000 156.2000 46.2000 ;
	    RECT 153.4000 45.6000 155.5000 45.7000 ;
	    RECT 153.4000 45.4000 155.4000 45.6000 ;
	    RECT 152.6000 44.8000 153.0000 45.2000 ;
	    RECT 148.6000 43.8000 149.0000 44.6000 ;
	    RECT 149.4000 43.5000 149.7000 44.8000 ;
	    RECT 150.2000 44.1000 150.6000 44.2000 ;
	    RECT 150.2000 43.8000 151.3000 44.1000 ;
	    RECT 151.8000 43.8000 152.2000 44.6000 ;
	    RECT 147.9000 43.2000 149.7000 43.5000 ;
	    RECT 147.9000 43.1000 148.2000 43.2000 ;
	    RECT 147.8000 41.1000 148.2000 43.1000 ;
	    RECT 149.4000 43.1000 149.7000 43.2000 ;
	    RECT 151.0000 43.5000 151.3000 43.8000 ;
	    RECT 152.6000 43.5000 152.9000 44.8000 ;
	    RECT 151.0000 43.2000 152.9000 43.5000 ;
	    RECT 149.4000 41.1000 149.8000 43.1000 ;
	    RECT 151.0000 41.1000 151.4000 43.2000 ;
	    RECT 152.6000 43.1000 152.9000 43.2000 ;
	    RECT 152.6000 41.1000 153.0000 43.1000 ;
	    RECT 153.4000 41.1000 153.8000 45.4000 ;
	    RECT 155.9000 45.1000 156.2000 45.8000 ;
	    RECT 156.7000 46.8000 158.5000 47.1000 ;
	    RECT 159.8000 46.8000 160.2000 47.6000 ;
	    RECT 156.7000 45.2000 157.0000 46.8000 ;
	    RECT 157.8000 45.8000 158.6000 46.2000 ;
	    RECT 155.5000 44.8000 156.2000 45.1000 ;
	    RECT 156.6000 44.8000 157.0000 45.2000 ;
	    RECT 159.0000 44.8000 159.4000 45.6000 ;
	    RECT 155.5000 41.1000 155.9000 44.8000 ;
	    RECT 156.7000 43.5000 157.0000 44.8000 ;
	    RECT 157.4000 43.8000 157.8000 44.6000 ;
	    RECT 156.7000 43.2000 158.5000 43.5000 ;
	    RECT 156.7000 43.1000 157.0000 43.2000 ;
	    RECT 156.6000 41.1000 157.0000 43.1000 ;
	    RECT 158.2000 43.1000 158.5000 43.2000 ;
	    RECT 158.2000 41.1000 158.6000 43.1000 ;
	    RECT 160.6000 41.1000 161.0000 47.9000 ;
	    RECT 164.0000 47.1000 164.4000 49.9000 ;
	    RECT 166.0000 47.1000 166.4000 49.9000 ;
	    RECT 164.0000 46.9000 164.9000 47.1000 ;
	    RECT 164.1000 46.8000 164.9000 46.9000 ;
	    RECT 163.0000 45.8000 163.8000 46.2000 ;
	    RECT 164.6000 45.2000 164.9000 46.8000 ;
	    RECT 165.5000 46.9000 166.4000 47.1000 ;
	    RECT 168.6000 47.9000 169.0000 49.9000 ;
	    RECT 170.2000 48.9000 170.6000 49.9000 ;
	    RECT 165.5000 46.8000 166.3000 46.9000 ;
	    RECT 165.5000 45.2000 165.8000 46.8000 ;
	    RECT 168.6000 46.2000 168.9000 47.9000 ;
	    RECT 170.2000 47.8000 170.5000 48.9000 ;
	    RECT 171.0000 47.8000 171.4000 48.6000 ;
	    RECT 169.3000 47.5000 170.5000 47.8000 ;
	    RECT 166.6000 45.8000 167.4000 46.2000 ;
	    RECT 168.6000 45.8000 169.0000 46.2000 ;
	    RECT 169.3000 46.0000 169.6000 47.5000 ;
	    RECT 164.6000 44.8000 165.0000 45.2000 ;
	    RECT 165.4000 44.8000 165.8000 45.2000 ;
	    RECT 168.6000 45.2000 168.9000 45.8000 ;
	    RECT 169.3000 45.7000 169.7000 46.0000 ;
	    RECT 169.3000 45.6000 171.4000 45.7000 ;
	    RECT 169.4000 45.4000 171.4000 45.6000 ;
	    RECT 168.6000 45.1000 169.0000 45.2000 ;
	    RECT 168.6000 44.8000 169.3000 45.1000 ;
	    RECT 163.8000 43.8000 164.2000 44.6000 ;
	    RECT 164.6000 43.5000 164.9000 44.8000 ;
	    RECT 163.1000 43.2000 164.9000 43.5000 ;
	    RECT 163.1000 43.1000 163.4000 43.2000 ;
	    RECT 163.0000 41.1000 163.4000 43.1000 ;
	    RECT 164.6000 43.1000 164.9000 43.2000 ;
	    RECT 165.5000 43.5000 165.8000 44.8000 ;
	    RECT 166.2000 43.8000 166.6000 44.6000 ;
	    RECT 165.5000 43.2000 167.3000 43.5000 ;
	    RECT 165.5000 43.1000 165.8000 43.2000 ;
	    RECT 164.6000 41.1000 165.0000 43.1000 ;
	    RECT 165.4000 41.1000 165.8000 43.1000 ;
	    RECT 167.0000 43.1000 167.3000 43.2000 ;
	    RECT 167.0000 41.1000 167.4000 43.1000 ;
	    RECT 168.9000 41.1000 169.3000 44.8000 ;
	    RECT 171.0000 41.1000 171.4000 45.4000 ;
	    RECT 0.6000 37.9000 1.0000 39.9000 ;
	    RECT 0.7000 37.8000 1.0000 37.9000 ;
	    RECT 2.2000 37.9000 2.6000 39.9000 ;
	    RECT 3.8000 37.9000 4.2000 39.9000 ;
	    RECT 2.2000 37.8000 2.5000 37.9000 ;
	    RECT 0.7000 37.5000 2.5000 37.8000 ;
	    RECT 3.9000 37.8000 4.2000 37.9000 ;
	    RECT 5.4000 37.9000 5.8000 39.9000 ;
	    RECT 7.8000 37.9000 8.2000 39.9000 ;
	    RECT 5.4000 37.8000 5.7000 37.9000 ;
	    RECT 3.9000 37.5000 5.7000 37.8000 ;
	    RECT 7.9000 37.8000 8.2000 37.9000 ;
	    RECT 9.4000 37.9000 9.8000 39.9000 ;
	    RECT 10.2000 37.9000 10.6000 39.9000 ;
	    RECT 9.4000 37.8000 9.7000 37.9000 ;
	    RECT 7.9000 37.5000 9.7000 37.8000 ;
	    RECT 0.7000 36.2000 1.0000 37.5000 ;
	    RECT 1.4000 36.4000 1.8000 37.2000 ;
	    RECT 3.9000 36.2000 4.2000 37.5000 ;
	    RECT 4.6000 36.4000 5.0000 37.2000 ;
	    RECT 8.6000 36.4000 9.0000 37.2000 ;
	    RECT 9.4000 36.2000 9.7000 37.5000 ;
	    RECT 10.3000 37.8000 10.6000 37.9000 ;
	    RECT 11.8000 37.9000 12.2000 39.9000 ;
	    RECT 13.4000 37.9000 13.8000 39.9000 ;
	    RECT 11.8000 37.8000 12.1000 37.9000 ;
	    RECT 10.3000 37.5000 12.1000 37.8000 ;
	    RECT 13.5000 37.8000 13.8000 37.9000 ;
	    RECT 15.0000 37.9000 15.4000 39.9000 ;
	    RECT 15.0000 37.8000 15.3000 37.9000 ;
	    RECT 13.5000 37.5000 15.3000 37.8000 ;
	    RECT 17.4000 37.8000 17.8000 39.9000 ;
	    RECT 19.0000 37.9000 19.4000 39.9000 ;
	    RECT 19.0000 37.8000 19.3000 37.9000 ;
	    RECT 17.4000 37.5000 19.3000 37.8000 ;
	    RECT 10.3000 36.2000 10.6000 37.5000 ;
	    RECT 11.0000 36.4000 11.4000 37.2000 ;
	    RECT 13.5000 36.2000 13.8000 37.5000 ;
	    RECT 14.2000 37.1000 14.6000 37.2000 ;
	    RECT 17.4000 37.1000 17.7000 37.5000 ;
	    RECT 14.2000 36.8000 17.7000 37.1000 ;
	    RECT 14.2000 36.4000 14.6000 36.8000 ;
	    RECT 18.2000 36.4000 18.6000 37.2000 ;
	    RECT 19.0000 36.2000 19.3000 37.5000 ;
	    RECT 19.8000 36.8000 20.2000 37.2000 ;
	    RECT 0.6000 35.8000 1.0000 36.2000 ;
	    RECT 0.7000 34.2000 1.0000 35.8000 ;
	    RECT 3.0000 35.4000 3.4000 36.2000 ;
	    RECT 3.8000 35.8000 4.2000 36.2000 ;
	    RECT 1.8000 34.8000 2.6000 35.2000 ;
	    RECT 3.9000 34.2000 4.2000 35.8000 ;
	    RECT 6.2000 35.4000 6.6000 36.2000 ;
	    RECT 9.4000 35.8000 9.8000 36.2000 ;
	    RECT 10.2000 35.8000 10.6000 36.2000 ;
	    RECT 13.4000 35.8000 13.8000 36.2000 ;
	    RECT 5.0000 34.8000 5.8000 35.2000 ;
	    RECT 7.8000 34.8000 8.6000 35.2000 ;
	    RECT 9.4000 34.2000 9.7000 35.8000 ;
	    RECT 0.7000 33.9000 1.8000 34.2000 ;
	    RECT 3.9000 33.9000 5.0000 34.2000 ;
	    RECT 8.9000 34.1000 9.7000 34.2000 ;
	    RECT 1.2000 33.8000 1.8000 33.9000 ;
	    RECT 4.4000 33.8000 5.0000 33.9000 ;
	    RECT 8.8000 33.9000 9.7000 34.1000 ;
	    RECT 10.3000 34.2000 10.6000 35.8000 ;
	    RECT 11.4000 34.8000 12.2000 35.2000 ;
	    RECT 13.5000 34.2000 13.8000 35.8000 ;
	    RECT 14.6000 34.8000 15.4000 35.2000 ;
	    RECT 16.6000 34.8000 17.0000 36.2000 ;
	    RECT 19.0000 35.8000 19.4000 36.2000 ;
	    RECT 19.8000 36.1000 20.1000 36.8000 ;
	    RECT 20.6000 36.1000 21.0000 39.9000 ;
	    RECT 23.0000 37.8000 23.4000 39.9000 ;
	    RECT 24.6000 37.9000 25.0000 39.9000 ;
	    RECT 24.6000 37.8000 24.9000 37.9000 ;
	    RECT 23.0000 37.5000 24.9000 37.8000 ;
	    RECT 23.0000 37.2000 23.3000 37.5000 ;
	    RECT 23.0000 36.8000 23.4000 37.2000 ;
	    RECT 19.8000 35.8000 21.0000 36.1000 ;
	    RECT 21.4000 35.8000 21.8000 36.6000 ;
	    RECT 23.8000 36.4000 24.2000 37.2000 ;
	    RECT 24.6000 36.2000 24.9000 37.5000 ;
	    RECT 25.7000 36.2000 26.1000 39.9000 ;
	    RECT 17.4000 34.8000 18.2000 35.2000 ;
	    RECT 19.0000 34.2000 19.3000 35.8000 ;
	    RECT 10.3000 34.1000 11.1000 34.2000 ;
	    RECT 13.5000 34.1000 14.3000 34.2000 ;
	    RECT 18.5000 34.1000 19.3000 34.2000 ;
	    RECT 10.3000 33.9000 11.2000 34.1000 ;
	    RECT 13.5000 33.9000 14.4000 34.1000 ;
	    RECT 1.2000 31.1000 1.6000 33.8000 ;
	    RECT 4.4000 31.1000 4.8000 33.8000 ;
	    RECT 8.8000 31.1000 9.2000 33.9000 ;
	    RECT 10.8000 31.1000 11.2000 33.9000 ;
	    RECT 14.0000 31.1000 14.4000 33.9000 ;
	    RECT 18.4000 33.9000 19.3000 34.1000 ;
	    RECT 18.4000 31.1000 18.8000 33.9000 ;
	    RECT 20.6000 33.1000 21.0000 35.8000 ;
	    RECT 22.2000 35.4000 22.6000 36.2000 ;
	    RECT 24.6000 35.8000 25.0000 36.2000 ;
	    RECT 25.4000 35.9000 26.1000 36.2000 ;
	    RECT 23.0000 34.8000 23.8000 35.2000 ;
	    RECT 24.6000 34.2000 24.9000 35.8000 ;
	    RECT 24.1000 34.1000 24.9000 34.2000 ;
	    RECT 24.0000 33.9000 24.9000 34.1000 ;
	    RECT 25.4000 35.2000 25.7000 35.9000 ;
	    RECT 27.8000 35.6000 28.2000 39.9000 ;
	    RECT 29.4000 37.9000 29.8000 39.9000 ;
	    RECT 29.5000 37.8000 29.8000 37.9000 ;
	    RECT 31.0000 37.9000 31.4000 39.9000 ;
	    RECT 31.0000 37.8000 31.3000 37.9000 ;
	    RECT 29.5000 37.5000 31.3000 37.8000 ;
	    RECT 30.2000 36.4000 30.6000 37.2000 ;
	    RECT 31.0000 36.2000 31.3000 37.5000 ;
	    RECT 32.1000 36.2000 32.5000 39.9000 ;
	    RECT 26.2000 35.4000 28.2000 35.6000 ;
	    RECT 28.6000 36.1000 29.0000 36.2000 ;
	    RECT 29.4000 36.1000 29.8000 36.2000 ;
	    RECT 28.6000 35.8000 29.8000 36.1000 ;
	    RECT 31.0000 35.8000 31.4000 36.2000 ;
	    RECT 31.8000 35.9000 32.5000 36.2000 ;
	    RECT 28.6000 35.4000 29.0000 35.8000 ;
	    RECT 26.1000 35.3000 28.2000 35.4000 ;
	    RECT 25.4000 34.8000 25.8000 35.2000 ;
	    RECT 26.1000 35.0000 26.5000 35.3000 ;
	    RECT 20.6000 32.8000 21.5000 33.1000 ;
	    RECT 21.1000 31.1000 21.5000 32.8000 ;
	    RECT 24.0000 31.1000 24.4000 33.9000 ;
	    RECT 25.4000 33.1000 25.7000 34.8000 ;
	    RECT 26.1000 33.5000 26.4000 35.0000 ;
	    RECT 29.4000 34.8000 30.2000 35.2000 ;
	    RECT 31.0000 34.2000 31.3000 35.8000 ;
	    RECT 30.5000 34.1000 31.3000 34.2000 ;
	    RECT 30.4000 33.9000 31.3000 34.1000 ;
	    RECT 31.8000 35.2000 32.1000 35.9000 ;
	    RECT 34.2000 35.6000 34.6000 39.9000 ;
	    RECT 32.6000 35.4000 34.6000 35.6000 ;
	    RECT 32.5000 35.3000 34.6000 35.4000 ;
	    RECT 31.8000 34.8000 32.2000 35.2000 ;
	    RECT 32.5000 35.0000 32.9000 35.3000 ;
	    RECT 26.1000 33.2000 27.3000 33.5000 ;
	    RECT 25.4000 31.1000 25.8000 33.1000 ;
	    RECT 27.0000 32.1000 27.3000 33.2000 ;
	    RECT 27.8000 32.4000 28.2000 33.2000 ;
	    RECT 27.0000 31.1000 27.4000 32.1000 ;
	    RECT 30.4000 31.1000 30.8000 33.9000 ;
	    RECT 31.8000 33.1000 32.1000 34.8000 ;
	    RECT 32.5000 33.5000 32.8000 35.0000 ;
	    RECT 35.0000 34.1000 35.4000 34.2000 ;
	    RECT 34.2000 33.8000 35.4000 34.1000 ;
	    RECT 32.5000 33.2000 33.7000 33.5000 ;
	    RECT 31.8000 31.1000 32.2000 33.1000 ;
	    RECT 33.4000 32.1000 33.7000 33.2000 ;
	    RECT 34.2000 33.2000 34.5000 33.8000 ;
	    RECT 35.0000 33.4000 35.4000 33.8000 ;
	    RECT 34.2000 32.4000 34.6000 33.2000 ;
	    RECT 35.8000 33.1000 36.2000 39.9000 ;
	    RECT 36.6000 36.1000 37.0000 36.6000 ;
	    RECT 37.4000 36.1000 37.8000 39.9000 ;
	    RECT 39.4000 36.8000 39.8000 37.2000 ;
	    RECT 39.4000 36.2000 39.7000 36.8000 ;
	    RECT 40.1000 36.2000 40.5000 39.9000 ;
	    RECT 36.6000 35.8000 37.8000 36.1000 ;
	    RECT 39.0000 35.9000 39.7000 36.2000 ;
	    RECT 40.0000 35.9000 40.5000 36.2000 ;
	    RECT 39.0000 35.8000 39.4000 35.9000 ;
	    RECT 35.8000 32.8000 36.7000 33.1000 ;
	    RECT 33.4000 31.1000 33.8000 32.1000 ;
	    RECT 36.3000 31.1000 36.7000 32.8000 ;
	    RECT 37.4000 31.1000 37.8000 35.8000 ;
	    RECT 39.0000 34.8000 39.4000 35.2000 ;
	    RECT 39.0000 34.2000 39.3000 34.8000 ;
	    RECT 40.0000 34.2000 40.3000 35.9000 ;
	    RECT 40.6000 34.4000 41.0000 35.2000 ;
	    RECT 39.0000 33.8000 40.3000 34.2000 ;
	    RECT 41.4000 34.1000 41.8000 34.2000 ;
	    RECT 42.2000 34.1000 42.6000 39.9000 ;
	    RECT 43.8000 35.6000 44.2000 39.9000 ;
	    RECT 45.9000 36.2000 46.3000 39.9000 ;
	    RECT 47.0000 37.9000 47.4000 39.9000 ;
	    RECT 47.1000 37.8000 47.4000 37.9000 ;
	    RECT 48.6000 37.9000 49.0000 39.9000 ;
	    RECT 48.6000 37.8000 48.9000 37.9000 ;
	    RECT 47.1000 37.5000 48.9000 37.8000 ;
	    RECT 47.1000 36.2000 47.4000 37.5000 ;
	    RECT 47.8000 36.4000 48.2000 37.2000 ;
	    RECT 45.9000 35.9000 46.6000 36.2000 ;
	    RECT 43.8000 35.4000 45.8000 35.6000 ;
	    RECT 43.8000 35.3000 45.9000 35.4000 ;
	    RECT 45.5000 35.0000 45.9000 35.3000 ;
	    RECT 46.3000 35.2000 46.6000 35.9000 ;
	    RECT 47.0000 35.8000 47.4000 36.2000 ;
	    RECT 41.0000 33.8000 42.6000 34.1000 ;
	    RECT 39.1000 33.1000 39.4000 33.8000 ;
	    RECT 41.0000 33.6000 41.4000 33.8000 ;
	    RECT 39.9000 33.1000 41.7000 33.3000 ;
	    RECT 39.0000 31.1000 39.4000 33.1000 ;
	    RECT 39.8000 33.0000 41.8000 33.1000 ;
	    RECT 39.8000 31.1000 40.2000 33.0000 ;
	    RECT 41.4000 31.1000 41.8000 33.0000 ;
	    RECT 42.2000 31.1000 42.6000 33.8000 ;
	    RECT 45.6000 33.5000 45.9000 35.0000 ;
	    RECT 46.2000 34.8000 46.6000 35.2000 ;
	    RECT 44.7000 33.2000 45.9000 33.5000 ;
	    RECT 43.8000 32.4000 44.2000 33.2000 ;
	    RECT 44.7000 32.1000 45.0000 33.2000 ;
	    RECT 46.3000 33.1000 46.6000 34.8000 ;
	    RECT 47.1000 34.2000 47.4000 35.8000 ;
	    RECT 49.4000 35.4000 49.8000 36.2000 ;
	    RECT 51.0000 36.1000 51.4000 39.9000 ;
	    RECT 51.8000 36.1000 52.2000 36.6000 ;
	    RECT 51.0000 35.8000 52.2000 36.1000 ;
	    RECT 48.2000 34.8000 49.0000 35.2000 ;
	    RECT 47.1000 34.1000 47.9000 34.2000 ;
	    RECT 47.1000 33.9000 48.9000 34.1000 ;
	    RECT 44.6000 31.1000 45.0000 32.1000 ;
	    RECT 46.2000 31.1000 46.6000 33.1000 ;
	    RECT 47.6000 33.8000 48.9000 33.9000 ;
	    RECT 47.6000 31.1000 48.0000 33.8000 ;
	    RECT 48.6000 33.2000 48.9000 33.8000 ;
	    RECT 48.6000 32.8000 49.0000 33.2000 ;
	    RECT 51.0000 31.1000 51.4000 35.8000 ;
	    RECT 52.6000 33.1000 53.0000 39.9000 ;
	    RECT 54.2000 37.9000 54.6000 39.9000 ;
	    RECT 54.3000 37.8000 54.6000 37.9000 ;
	    RECT 55.8000 37.9000 56.2000 39.9000 ;
	    RECT 55.8000 37.8000 56.1000 37.9000 ;
	    RECT 54.3000 37.5000 56.1000 37.8000 ;
	    RECT 54.3000 36.2000 54.6000 37.5000 ;
	    RECT 55.0000 36.4000 55.4000 37.2000 ;
	    RECT 54.2000 35.8000 54.6000 36.2000 ;
	    RECT 54.3000 34.2000 54.6000 35.8000 ;
	    RECT 56.6000 35.4000 57.0000 36.2000 ;
	    RECT 57.4000 35.8000 57.8000 36.6000 ;
	    RECT 55.4000 34.8000 56.2000 35.2000 ;
	    RECT 53.4000 33.4000 53.8000 34.2000 ;
	    RECT 54.3000 34.1000 55.1000 34.2000 ;
	    RECT 54.3000 33.9000 55.2000 34.1000 ;
	    RECT 52.1000 32.8000 53.0000 33.1000 ;
	    RECT 52.1000 31.1000 52.5000 32.8000 ;
	    RECT 54.8000 31.1000 55.2000 33.9000 ;
	    RECT 58.2000 33.2000 58.6000 39.9000 ;
	    RECT 57.4000 32.8000 58.6000 33.2000 ;
	    RECT 57.7000 31.1000 58.1000 32.8000 ;
	    RECT 62.2000 31.1000 62.6000 39.9000 ;
	    RECT 63.0000 37.9000 63.4000 39.9000 ;
	    RECT 63.1000 37.8000 63.4000 37.9000 ;
	    RECT 64.6000 37.9000 65.0000 39.9000 ;
	    RECT 66.2000 37.9000 66.6000 39.9000 ;
	    RECT 64.6000 37.8000 64.9000 37.9000 ;
	    RECT 63.1000 37.5000 64.9000 37.8000 ;
	    RECT 66.3000 37.8000 66.6000 37.9000 ;
	    RECT 67.8000 37.9000 68.2000 39.9000 ;
	    RECT 70.2000 37.9000 70.6000 39.9000 ;
	    RECT 67.8000 37.8000 68.1000 37.9000 ;
	    RECT 66.3000 37.5000 68.1000 37.8000 ;
	    RECT 70.3000 37.8000 70.6000 37.9000 ;
	    RECT 71.8000 37.8000 72.2000 39.9000 ;
	    RECT 72.6000 37.9000 73.0000 39.9000 ;
	    RECT 72.7000 37.8000 73.0000 37.9000 ;
	    RECT 74.2000 37.9000 74.6000 39.9000 ;
	    RECT 74.2000 37.8000 74.5000 37.9000 ;
	    RECT 70.3000 37.5000 72.1000 37.8000 ;
	    RECT 63.1000 36.2000 63.4000 37.5000 ;
	    RECT 63.8000 36.4000 64.2000 37.2000 ;
	    RECT 66.3000 36.2000 66.6000 37.5000 ;
	    RECT 67.0000 36.4000 67.4000 37.2000 ;
	    RECT 71.0000 36.4000 71.4000 37.2000 ;
	    RECT 71.8000 36.2000 72.1000 37.5000 ;
	    RECT 72.7000 37.5000 74.5000 37.8000 ;
	    RECT 72.7000 36.2000 73.0000 37.5000 ;
	    RECT 73.4000 36.4000 73.8000 37.2000 ;
	    RECT 76.2000 36.8000 76.6000 37.2000 ;
	    RECT 76.2000 36.2000 76.5000 36.8000 ;
	    RECT 76.9000 36.2000 77.3000 39.9000 ;
	    RECT 63.0000 35.8000 63.4000 36.2000 ;
	    RECT 63.1000 34.2000 63.4000 35.8000 ;
	    RECT 65.4000 35.4000 65.8000 36.2000 ;
	    RECT 66.2000 35.8000 66.6000 36.2000 ;
	    RECT 64.2000 34.8000 65.0000 35.2000 ;
	    RECT 66.3000 34.2000 66.6000 35.8000 ;
	    RECT 68.6000 35.4000 69.0000 36.2000 ;
	    RECT 71.8000 35.8000 72.2000 36.2000 ;
	    RECT 72.6000 35.8000 73.0000 36.2000 ;
	    RECT 75.8000 35.9000 76.5000 36.2000 ;
	    RECT 76.8000 35.9000 77.3000 36.2000 ;
	    RECT 75.8000 35.8000 76.2000 35.9000 ;
	    RECT 67.4000 34.8000 68.2000 35.2000 ;
	    RECT 70.2000 34.8000 71.0000 35.2000 ;
	    RECT 71.8000 34.2000 72.1000 35.8000 ;
	    RECT 63.1000 34.1000 63.9000 34.2000 ;
	    RECT 66.3000 34.1000 67.1000 34.2000 ;
	    RECT 71.3000 34.1000 72.1000 34.2000 ;
	    RECT 63.1000 33.9000 64.0000 34.1000 ;
	    RECT 66.3000 33.9000 67.2000 34.1000 ;
	    RECT 63.6000 31.1000 64.0000 33.9000 ;
	    RECT 66.8000 31.1000 67.2000 33.9000 ;
	    RECT 71.2000 33.9000 72.1000 34.1000 ;
	    RECT 72.7000 34.2000 73.0000 35.8000 ;
	    RECT 73.8000 34.8000 74.6000 35.2000 ;
	    RECT 75.8000 35.1000 76.2000 35.2000 ;
	    RECT 76.8000 35.1000 77.1000 35.9000 ;
	    RECT 75.8000 34.8000 77.1000 35.1000 ;
	    RECT 76.8000 34.2000 77.1000 34.8000 ;
	    RECT 77.4000 34.4000 77.8000 35.2000 ;
	    RECT 72.7000 34.1000 73.5000 34.2000 ;
	    RECT 72.7000 33.9000 73.6000 34.1000 ;
	    RECT 71.2000 31.1000 71.6000 33.9000 ;
	    RECT 73.2000 31.1000 73.6000 33.9000 ;
	    RECT 75.8000 33.8000 77.1000 34.2000 ;
	    RECT 78.2000 34.1000 78.6000 34.2000 ;
	    RECT 79.0000 34.1000 79.4000 39.9000 ;
	    RECT 77.8000 33.8000 79.4000 34.1000 ;
	    RECT 75.9000 33.1000 76.2000 33.8000 ;
	    RECT 77.8000 33.6000 78.2000 33.8000 ;
	    RECT 76.7000 33.1000 78.5000 33.3000 ;
	    RECT 75.8000 31.1000 76.2000 33.1000 ;
	    RECT 76.6000 33.0000 78.6000 33.1000 ;
	    RECT 76.6000 31.1000 77.0000 33.0000 ;
	    RECT 78.2000 31.1000 78.6000 33.0000 ;
	    RECT 79.0000 31.1000 79.4000 33.8000 ;
	    RECT 81.4000 31.1000 81.8000 39.9000 ;
	    RECT 83.8000 36.1000 84.2000 39.9000 ;
	    RECT 84.6000 36.1000 85.0000 36.6000 ;
	    RECT 83.8000 35.8000 85.0000 36.1000 ;
	    RECT 83.8000 31.1000 84.2000 35.8000 ;
	    RECT 85.4000 33.1000 85.8000 39.9000 ;
	    RECT 87.8000 36.1000 88.2000 39.9000 ;
	    RECT 88.6000 36.8000 89.0000 37.2000 ;
	    RECT 88.6000 36.1000 88.9000 36.8000 ;
	    RECT 87.8000 35.8000 88.9000 36.1000 ;
	    RECT 86.2000 33.4000 86.6000 34.2000 ;
	    RECT 84.9000 32.8000 85.8000 33.1000 ;
	    RECT 84.9000 31.1000 85.3000 32.8000 ;
	    RECT 87.8000 31.1000 88.2000 35.8000 ;
	    RECT 88.6000 33.4000 89.0000 34.2000 ;
	    RECT 89.4000 33.1000 89.8000 39.9000 ;
	    RECT 90.2000 35.8000 90.6000 36.6000 ;
	    RECT 91.0000 35.6000 91.4000 39.9000 ;
	    RECT 93.1000 36.2000 93.5000 39.9000 ;
	    RECT 94.2000 37.9000 94.6000 39.9000 ;
	    RECT 94.3000 37.8000 94.6000 37.9000 ;
	    RECT 95.8000 37.9000 96.2000 39.9000 ;
	    RECT 97.4000 37.9000 97.8000 39.9000 ;
	    RECT 95.8000 37.8000 96.1000 37.9000 ;
	    RECT 94.3000 37.5000 96.1000 37.8000 ;
	    RECT 97.5000 37.8000 97.8000 37.9000 ;
	    RECT 99.0000 37.9000 99.4000 39.9000 ;
	    RECT 99.0000 37.8000 99.3000 37.9000 ;
	    RECT 97.5000 37.5000 99.3000 37.8000 ;
	    RECT 94.3000 36.2000 94.6000 37.5000 ;
	    RECT 95.0000 36.4000 95.4000 37.2000 ;
	    RECT 97.5000 36.2000 97.8000 37.5000 ;
	    RECT 98.2000 36.4000 98.6000 37.2000 ;
	    RECT 100.9000 36.2000 101.3000 39.9000 ;
	    RECT 93.1000 35.9000 93.8000 36.2000 ;
	    RECT 91.0000 35.4000 93.0000 35.6000 ;
	    RECT 91.0000 35.3000 93.1000 35.4000 ;
	    RECT 92.7000 35.0000 93.1000 35.3000 ;
	    RECT 93.5000 35.2000 93.8000 35.9000 ;
	    RECT 94.2000 35.8000 94.6000 36.2000 ;
	    RECT 92.8000 33.5000 93.1000 35.0000 ;
	    RECT 93.4000 34.8000 93.8000 35.2000 ;
	    RECT 91.9000 33.2000 93.1000 33.5000 ;
	    RECT 89.4000 32.8000 90.3000 33.1000 ;
	    RECT 89.9000 31.1000 90.3000 32.8000 ;
	    RECT 91.0000 32.4000 91.4000 33.2000 ;
	    RECT 91.9000 32.1000 92.2000 33.2000 ;
	    RECT 93.5000 33.1000 93.8000 34.8000 ;
	    RECT 94.3000 34.2000 94.6000 35.8000 ;
	    RECT 96.6000 35.4000 97.0000 36.2000 ;
	    RECT 97.4000 35.8000 97.8000 36.2000 ;
	    RECT 95.4000 34.8000 96.2000 35.2000 ;
	    RECT 97.5000 34.2000 97.8000 35.8000 ;
	    RECT 99.8000 35.4000 100.2000 36.2000 ;
	    RECT 100.6000 35.9000 101.3000 36.2000 ;
	    RECT 100.6000 35.2000 100.9000 35.9000 ;
	    RECT 103.0000 35.6000 103.4000 39.9000 ;
	    RECT 101.4000 35.4000 103.4000 35.6000 ;
	    RECT 101.3000 35.3000 103.4000 35.4000 ;
	    RECT 98.6000 34.8000 99.4000 35.2000 ;
	    RECT 100.6000 34.8000 101.0000 35.2000 ;
	    RECT 101.3000 35.0000 101.7000 35.3000 ;
	    RECT 103.8000 35.1000 104.2000 35.2000 ;
	    RECT 104.6000 35.1000 105.0000 39.9000 ;
	    RECT 105.4000 37.9000 105.8000 39.9000 ;
	    RECT 105.5000 37.8000 105.8000 37.9000 ;
	    RECT 107.0000 37.9000 107.4000 39.9000 ;
	    RECT 109.4000 37.9000 109.8000 39.9000 ;
	    RECT 107.0000 37.8000 107.3000 37.9000 ;
	    RECT 105.5000 37.5000 107.3000 37.8000 ;
	    RECT 109.5000 37.8000 109.8000 37.9000 ;
	    RECT 111.0000 37.9000 111.4000 39.9000 ;
	    RECT 111.0000 37.8000 111.3000 37.9000 ;
	    RECT 109.5000 37.5000 111.3000 37.8000 ;
	    RECT 105.5000 36.2000 105.8000 37.5000 ;
	    RECT 106.2000 36.4000 106.6000 37.2000 ;
	    RECT 110.2000 36.4000 110.6000 37.2000 ;
	    RECT 111.0000 36.2000 111.3000 37.5000 ;
	    RECT 105.4000 35.8000 105.8000 36.2000 ;
	    RECT 94.3000 34.1000 95.1000 34.2000 ;
	    RECT 94.3000 33.9000 95.2000 34.1000 ;
	    RECT 97.5000 33.9000 98.6000 34.2000 ;
	    RECT 91.8000 31.1000 92.2000 32.1000 ;
	    RECT 93.4000 31.1000 93.8000 33.1000 ;
	    RECT 94.8000 31.1000 95.2000 33.9000 ;
	    RECT 98.0000 33.8000 98.6000 33.9000 ;
	    RECT 98.0000 31.1000 98.4000 33.8000 ;
	    RECT 100.6000 33.1000 100.9000 34.8000 ;
	    RECT 101.3000 33.5000 101.6000 35.0000 ;
	    RECT 103.8000 34.8000 105.0000 35.1000 ;
	    RECT 102.0000 34.2000 102.4000 34.6000 ;
	    RECT 102.1000 33.8000 102.6000 34.2000 ;
	    RECT 101.3000 33.2000 102.5000 33.5000 ;
	    RECT 100.6000 31.1000 101.0000 33.1000 ;
	    RECT 102.2000 32.1000 102.5000 33.2000 ;
	    RECT 102.2000 31.1000 102.6000 32.1000 ;
	    RECT 104.6000 31.1000 105.0000 34.8000 ;
	    RECT 105.5000 34.2000 105.8000 35.8000 ;
	    RECT 108.6000 36.1000 109.0000 36.2000 ;
	    RECT 109.4000 36.1000 109.8000 36.2000 ;
	    RECT 108.6000 35.8000 109.8000 36.1000 ;
	    RECT 111.0000 35.8000 111.4000 36.2000 ;
	    RECT 108.6000 35.4000 109.0000 35.8000 ;
	    RECT 106.6000 34.8000 107.4000 35.2000 ;
	    RECT 109.4000 34.8000 110.2000 35.2000 ;
	    RECT 111.0000 34.2000 111.3000 35.8000 ;
	    RECT 113.4000 35.6000 113.8000 39.9000 ;
	    RECT 115.5000 36.2000 115.9000 39.9000 ;
	    RECT 116.6000 37.9000 117.0000 39.9000 ;
	    RECT 116.7000 37.8000 117.0000 37.9000 ;
	    RECT 118.2000 37.9000 118.6000 39.9000 ;
	    RECT 120.6000 37.9000 121.0000 39.9000 ;
	    RECT 118.2000 37.8000 118.5000 37.9000 ;
	    RECT 116.7000 37.5000 118.5000 37.8000 ;
	    RECT 120.7000 37.8000 121.0000 37.9000 ;
	    RECT 122.2000 37.9000 122.6000 39.9000 ;
	    RECT 122.2000 37.8000 122.5000 37.9000 ;
	    RECT 120.7000 37.5000 122.5000 37.8000 ;
	    RECT 116.7000 36.2000 117.0000 37.5000 ;
	    RECT 117.4000 36.4000 117.8000 37.2000 ;
	    RECT 121.4000 36.4000 121.8000 37.2000 ;
	    RECT 122.2000 36.2000 122.5000 37.5000 ;
	    RECT 115.5000 35.9000 116.2000 36.2000 ;
	    RECT 113.4000 35.4000 115.4000 35.6000 ;
	    RECT 113.4000 35.3000 115.5000 35.4000 ;
	    RECT 115.1000 35.0000 115.5000 35.3000 ;
	    RECT 115.9000 35.2000 116.2000 35.9000 ;
	    RECT 116.6000 35.8000 117.0000 36.2000 ;
	    RECT 105.5000 34.1000 106.3000 34.2000 ;
	    RECT 110.5000 34.1000 111.3000 34.2000 ;
	    RECT 105.5000 33.9000 106.4000 34.1000 ;
	    RECT 106.0000 31.1000 106.4000 33.9000 ;
	    RECT 110.4000 33.9000 111.3000 34.1000 ;
	    RECT 110.4000 31.1000 110.8000 33.9000 ;
	    RECT 115.2000 33.5000 115.5000 35.0000 ;
	    RECT 115.8000 34.8000 116.2000 35.2000 ;
	    RECT 115.9000 34.2000 116.2000 34.8000 ;
	    RECT 115.8000 33.8000 116.2000 34.2000 ;
	    RECT 116.7000 34.2000 117.0000 35.8000 ;
	    RECT 119.0000 35.4000 119.4000 36.2000 ;
	    RECT 119.8000 35.4000 120.2000 36.2000 ;
	    RECT 122.2000 35.8000 122.6000 36.2000 ;
	    RECT 123.8000 36.1000 124.2000 39.9000 ;
	    RECT 125.4000 37.9000 125.8000 39.9000 ;
	    RECT 125.5000 37.8000 125.8000 37.9000 ;
	    RECT 127.0000 37.9000 127.4000 39.9000 ;
	    RECT 127.0000 37.8000 127.3000 37.9000 ;
	    RECT 125.5000 37.5000 127.3000 37.8000 ;
	    RECT 126.2000 36.4000 126.6000 37.2000 ;
	    RECT 127.0000 36.2000 127.3000 37.5000 ;
	    RECT 124.6000 36.1000 125.0000 36.2000 ;
	    RECT 123.8000 35.8000 125.0000 36.1000 ;
	    RECT 117.8000 34.8000 118.6000 35.2000 ;
	    RECT 120.6000 34.8000 121.4000 35.2000 ;
	    RECT 122.2000 34.2000 122.5000 35.8000 ;
	    RECT 116.7000 34.1000 117.5000 34.2000 ;
	    RECT 121.7000 34.1000 122.5000 34.2000 ;
	    RECT 116.7000 33.9000 117.6000 34.1000 ;
	    RECT 114.3000 33.2000 115.5000 33.5000 ;
	    RECT 112.6000 33.1000 113.0000 33.2000 ;
	    RECT 113.4000 33.1000 113.8000 33.2000 ;
	    RECT 112.6000 32.8000 113.8000 33.1000 ;
	    RECT 113.4000 32.4000 113.8000 32.8000 ;
	    RECT 114.3000 32.1000 114.6000 33.2000 ;
	    RECT 115.9000 33.1000 116.2000 33.8000 ;
	    RECT 114.2000 31.1000 114.6000 32.1000 ;
	    RECT 115.8000 31.1000 116.2000 33.1000 ;
	    RECT 117.2000 33.1000 117.6000 33.9000 ;
	    RECT 121.6000 33.9000 122.5000 34.1000 ;
	    RECT 118.2000 33.1000 118.6000 33.2000 ;
	    RECT 117.2000 32.8000 118.6000 33.1000 ;
	    RECT 117.2000 31.1000 117.6000 32.8000 ;
	    RECT 121.6000 31.1000 122.0000 33.9000 ;
	    RECT 123.8000 31.1000 124.2000 35.8000 ;
	    RECT 124.6000 35.4000 125.0000 35.8000 ;
	    RECT 127.0000 35.8000 127.4000 36.2000 ;
	    RECT 125.4000 34.8000 126.2000 35.2000 ;
	    RECT 127.0000 34.2000 127.3000 35.8000 ;
	    RECT 126.5000 34.1000 127.3000 34.2000 ;
	    RECT 126.4000 33.9000 127.3000 34.1000 ;
	    RECT 126.4000 31.1000 126.8000 33.9000 ;
	    RECT 128.6000 31.1000 129.0000 39.9000 ;
	    RECT 129.4000 35.6000 129.8000 39.9000 ;
	    RECT 131.5000 36.2000 131.9000 39.9000 ;
	    RECT 132.6000 37.1000 133.0000 37.2000 ;
	    RECT 133.4000 37.1000 133.8000 39.9000 ;
	    RECT 132.6000 36.8000 133.8000 37.1000 ;
	    RECT 131.5000 35.9000 132.2000 36.2000 ;
	    RECT 129.4000 35.4000 131.4000 35.6000 ;
	    RECT 129.4000 35.3000 131.5000 35.4000 ;
	    RECT 131.1000 35.0000 131.5000 35.3000 ;
	    RECT 131.9000 35.2000 132.2000 35.9000 ;
	    RECT 131.2000 33.5000 131.5000 35.0000 ;
	    RECT 131.8000 34.8000 132.2000 35.2000 ;
	    RECT 131.9000 34.1000 132.2000 34.8000 ;
	    RECT 132.6000 34.8000 133.0000 35.2000 ;
	    RECT 132.6000 34.1000 132.9000 34.8000 ;
	    RECT 131.8000 33.8000 132.9000 34.1000 ;
	    RECT 130.3000 33.2000 131.5000 33.5000 ;
	    RECT 129.4000 32.4000 129.8000 33.2000 ;
	    RECT 130.3000 32.1000 130.6000 33.2000 ;
	    RECT 131.9000 33.1000 132.2000 33.8000 ;
	    RECT 130.2000 31.1000 130.6000 32.1000 ;
	    RECT 131.8000 31.1000 132.2000 33.1000 ;
	    RECT 133.4000 31.1000 133.8000 36.8000 ;
	    RECT 134.2000 35.8000 134.6000 36.6000 ;
	    RECT 135.0000 33.1000 135.4000 39.9000 ;
	    RECT 137.4000 37.9000 137.8000 39.9000 ;
	    RECT 137.5000 37.8000 137.8000 37.9000 ;
	    RECT 139.0000 37.9000 139.4000 39.9000 ;
	    RECT 139.0000 37.8000 139.3000 37.9000 ;
	    RECT 137.5000 37.5000 139.3000 37.8000 ;
	    RECT 138.2000 36.4000 138.6000 37.2000 ;
	    RECT 139.0000 36.2000 139.3000 37.5000 ;
	    RECT 140.6000 37.1000 141.0000 39.9000 ;
	    RECT 142.2000 37.9000 142.6000 39.9000 ;
	    RECT 142.3000 37.8000 142.6000 37.9000 ;
	    RECT 143.8000 37.9000 144.2000 39.9000 ;
	    RECT 146.2000 37.9000 146.6000 39.9000 ;
	    RECT 143.8000 37.8000 144.1000 37.9000 ;
	    RECT 142.3000 37.5000 144.1000 37.8000 ;
	    RECT 146.3000 37.8000 146.6000 37.9000 ;
	    RECT 147.8000 37.9000 148.2000 39.9000 ;
	    RECT 148.6000 37.9000 149.0000 39.9000 ;
	    RECT 147.8000 37.8000 148.1000 37.9000 ;
	    RECT 146.3000 37.5000 148.1000 37.8000 ;
	    RECT 140.6000 36.8000 141.7000 37.1000 ;
	    RECT 139.0000 35.8000 139.4000 36.2000 ;
	    RECT 139.8000 35.8000 140.2000 36.6000 ;
	    RECT 137.4000 34.8000 138.2000 35.2000 ;
	    RECT 139.0000 34.2000 139.3000 35.8000 ;
	    RECT 135.8000 33.4000 136.2000 34.2000 ;
	    RECT 138.5000 34.1000 139.3000 34.2000 ;
	    RECT 138.4000 33.9000 139.3000 34.1000 ;
	    RECT 134.5000 32.8000 135.4000 33.1000 ;
	    RECT 134.5000 32.2000 134.9000 32.8000 ;
	    RECT 134.5000 31.8000 135.4000 32.2000 ;
	    RECT 134.5000 31.1000 134.9000 31.8000 ;
	    RECT 138.4000 31.1000 138.8000 33.9000 ;
	    RECT 140.6000 33.1000 141.0000 36.8000 ;
	    RECT 141.4000 36.2000 141.7000 36.8000 ;
	    RECT 142.3000 36.2000 142.6000 37.5000 ;
	    RECT 143.0000 36.4000 143.4000 37.2000 ;
	    RECT 143.8000 37.1000 144.1000 37.5000 ;
	    RECT 147.8000 37.2000 148.1000 37.5000 ;
	    RECT 148.7000 37.8000 149.0000 37.9000 ;
	    RECT 150.2000 37.9000 150.6000 39.9000 ;
	    RECT 150.2000 37.8000 150.5000 37.9000 ;
	    RECT 148.7000 37.5000 150.5000 37.8000 ;
	    RECT 146.2000 37.1000 146.6000 37.2000 ;
	    RECT 143.8000 36.8000 146.6000 37.1000 ;
	    RECT 147.0000 36.4000 147.4000 37.2000 ;
	    RECT 147.8000 36.8000 148.2000 37.2000 ;
	    RECT 147.8000 36.2000 148.1000 36.8000 ;
	    RECT 148.7000 36.2000 149.0000 37.5000 ;
	    RECT 149.4000 36.4000 149.8000 37.2000 ;
	    RECT 141.4000 35.8000 141.8000 36.2000 ;
	    RECT 142.2000 35.8000 142.6000 36.2000 ;
	    RECT 142.3000 34.2000 142.6000 35.8000 ;
	    RECT 144.6000 35.4000 145.0000 36.2000 ;
	    RECT 145.4000 35.4000 145.8000 36.2000 ;
	    RECT 147.8000 35.8000 148.2000 36.2000 ;
	    RECT 148.6000 35.8000 149.0000 36.2000 ;
	    RECT 143.0000 34.8000 144.2000 35.2000 ;
	    RECT 146.2000 34.8000 147.0000 35.2000 ;
	    RECT 147.8000 34.2000 148.1000 35.8000 ;
	    RECT 141.4000 33.4000 141.8000 34.2000 ;
	    RECT 142.3000 34.1000 143.1000 34.2000 ;
	    RECT 147.3000 34.1000 148.1000 34.2000 ;
	    RECT 142.3000 33.9000 143.2000 34.1000 ;
	    RECT 140.1000 32.8000 141.0000 33.1000 ;
	    RECT 140.1000 31.1000 140.5000 32.8000 ;
	    RECT 142.8000 31.1000 143.2000 33.9000 ;
	    RECT 147.2000 33.9000 148.1000 34.1000 ;
	    RECT 148.7000 34.2000 149.0000 35.8000 ;
	    RECT 149.8000 34.8000 150.6000 35.2000 ;
	    RECT 151.8000 35.1000 152.2000 39.9000 ;
	    RECT 154.2000 37.9000 154.6000 39.9000 ;
	    RECT 154.3000 37.8000 154.6000 37.9000 ;
	    RECT 155.8000 37.9000 156.2000 39.9000 ;
	    RECT 155.8000 37.8000 156.1000 37.9000 ;
	    RECT 154.3000 37.5000 156.1000 37.8000 ;
	    RECT 155.8000 37.2000 156.1000 37.5000 ;
	    RECT 155.0000 36.4000 155.4000 37.2000 ;
	    RECT 155.8000 36.8000 156.2000 37.2000 ;
	    RECT 155.8000 36.2000 156.1000 36.8000 ;
	    RECT 153.4000 35.1000 153.8000 36.2000 ;
	    RECT 155.8000 35.8000 156.2000 36.2000 ;
	    RECT 156.6000 35.9000 157.0000 39.9000 ;
	    RECT 158.2000 36.2000 158.6000 39.9000 ;
	    RECT 157.5000 35.9000 158.6000 36.2000 ;
	    RECT 159.0000 35.9000 159.4000 39.9000 ;
	    RECT 160.6000 36.2000 161.0000 39.9000 ;
	    RECT 162.2000 37.9000 162.6000 39.9000 ;
	    RECT 162.3000 37.8000 162.6000 37.9000 ;
	    RECT 163.8000 37.9000 164.2000 39.9000 ;
	    RECT 165.4000 37.9000 165.8000 39.9000 ;
	    RECT 163.8000 37.8000 164.1000 37.9000 ;
	    RECT 162.3000 37.5000 164.1000 37.8000 ;
	    RECT 165.5000 37.8000 165.8000 37.9000 ;
	    RECT 167.0000 37.9000 167.4000 39.9000 ;
	    RECT 167.0000 37.8000 167.3000 37.9000 ;
	    RECT 165.5000 37.5000 167.3000 37.8000 ;
	    RECT 163.0000 36.4000 163.4000 37.2000 ;
	    RECT 159.9000 35.9000 161.0000 36.2000 ;
	    RECT 163.8000 36.2000 164.1000 37.5000 ;
	    RECT 166.2000 36.4000 166.6000 37.2000 ;
	    RECT 167.0000 36.2000 167.3000 37.5000 ;
	    RECT 151.8000 34.8000 153.8000 35.1000 ;
	    RECT 154.2000 34.8000 155.0000 35.2000 ;
	    RECT 148.7000 34.1000 149.5000 34.2000 ;
	    RECT 148.7000 33.9000 149.6000 34.1000 ;
	    RECT 147.2000 31.1000 147.6000 33.9000 ;
	    RECT 149.2000 31.1000 149.6000 33.9000 ;
	    RECT 151.8000 31.1000 152.2000 34.8000 ;
	    RECT 155.8000 34.2000 156.1000 35.8000 ;
	    RECT 155.3000 34.1000 156.1000 34.2000 ;
	    RECT 155.2000 33.9000 156.1000 34.1000 ;
	    RECT 156.6000 34.8000 156.9000 35.9000 ;
	    RECT 157.5000 35.6000 157.8000 35.9000 ;
	    RECT 157.2000 35.2000 157.8000 35.6000 ;
	    RECT 155.2000 31.1000 155.6000 33.9000 ;
	    RECT 156.6000 31.1000 157.0000 34.8000 ;
	    RECT 157.5000 33.7000 157.8000 35.2000 ;
	    RECT 159.0000 34.8000 159.3000 35.9000 ;
	    RECT 159.9000 35.6000 160.2000 35.9000 ;
	    RECT 159.6000 35.2000 160.2000 35.6000 ;
	    RECT 163.8000 35.8000 164.2000 36.2000 ;
	    RECT 157.5000 33.4000 158.6000 33.7000 ;
	    RECT 158.2000 31.1000 158.6000 33.4000 ;
	    RECT 159.0000 31.1000 159.4000 34.8000 ;
	    RECT 159.9000 33.7000 160.2000 35.2000 ;
	    RECT 162.2000 34.8000 163.0000 35.2000 ;
	    RECT 163.8000 34.2000 164.1000 35.8000 ;
	    RECT 164.6000 35.4000 165.0000 36.2000 ;
	    RECT 167.0000 35.8000 167.4000 36.2000 ;
	    RECT 168.6000 36.1000 169.0000 39.9000 ;
	    RECT 169.4000 36.1000 169.8000 36.6000 ;
	    RECT 168.6000 35.8000 169.8000 36.1000 ;
	    RECT 170.2000 36.1000 170.6000 39.9000 ;
	    RECT 171.0000 36.1000 171.4000 36.2000 ;
	    RECT 170.2000 35.8000 171.4000 36.1000 ;
	    RECT 165.4000 34.8000 166.2000 35.2000 ;
	    RECT 167.0000 34.2000 167.3000 35.8000 ;
	    RECT 163.3000 34.1000 164.1000 34.2000 ;
	    RECT 166.5000 34.1000 167.3000 34.2000 ;
	    RECT 163.2000 33.9000 164.1000 34.1000 ;
	    RECT 166.4000 33.9000 167.3000 34.1000 ;
	    RECT 159.9000 33.4000 161.0000 33.7000 ;
	    RECT 160.6000 31.1000 161.0000 33.4000 ;
	    RECT 163.2000 31.1000 163.6000 33.9000 ;
	    RECT 166.4000 31.1000 166.8000 33.9000 ;
	    RECT 168.6000 31.1000 169.0000 35.8000 ;
	    RECT 170.2000 33.1000 170.6000 35.8000 ;
	    RECT 171.0000 33.4000 171.4000 34.2000 ;
	    RECT 169.7000 32.8000 170.6000 33.1000 ;
	    RECT 169.7000 31.1000 170.1000 32.8000 ;
	    RECT 1.4000 25.1000 1.8000 29.9000 ;
	    RECT 2.5000 29.2000 2.9000 29.9000 ;
	    RECT 2.2000 28.8000 2.9000 29.2000 ;
	    RECT 2.5000 28.2000 2.9000 28.8000 ;
	    RECT 2.5000 27.9000 3.4000 28.2000 ;
	    RECT 2.2000 25.1000 2.6000 25.2000 ;
	    RECT 1.4000 24.8000 2.6000 25.1000 ;
	    RECT 1.4000 21.1000 1.8000 24.8000 ;
	    RECT 2.2000 24.4000 2.6000 24.8000 ;
	    RECT 3.0000 21.1000 3.4000 27.9000 ;
	    RECT 4.6000 27.9000 5.0000 29.9000 ;
	    RECT 6.2000 28.9000 6.6000 29.9000 ;
	    RECT 8.4000 29.2000 8.8000 29.9000 ;
	    RECT 3.8000 26.8000 4.2000 27.6000 ;
	    RECT 4.6000 26.2000 4.9000 27.9000 ;
	    RECT 6.2000 27.8000 6.5000 28.9000 ;
	    RECT 5.3000 27.5000 6.5000 27.8000 ;
	    RECT 8.4000 28.8000 9.0000 29.2000 ;
	    RECT 4.6000 25.8000 5.0000 26.2000 ;
	    RECT 5.3000 26.0000 5.6000 27.5000 ;
	    RECT 6.1000 26.8000 6.6000 27.2000 ;
	    RECT 8.4000 27.1000 8.8000 28.8000 ;
	    RECT 7.9000 26.9000 8.8000 27.1000 ;
	    RECT 7.9000 26.8000 8.7000 26.9000 ;
	    RECT 6.0000 26.4000 6.4000 26.8000 ;
	    RECT 4.6000 25.1000 4.9000 25.8000 ;
	    RECT 5.3000 25.7000 5.7000 26.0000 ;
	    RECT 5.3000 25.6000 7.4000 25.7000 ;
	    RECT 5.4000 25.4000 7.4000 25.6000 ;
	    RECT 4.6000 24.8000 5.3000 25.1000 ;
	    RECT 4.9000 21.1000 5.3000 24.8000 ;
	    RECT 7.0000 21.1000 7.4000 25.4000 ;
	    RECT 7.9000 25.2000 8.2000 26.8000 ;
	    RECT 11.0000 26.2000 11.4000 29.9000 ;
	    RECT 12.6000 27.6000 13.0000 29.9000 ;
	    RECT 15.2000 29.2000 15.6000 29.9000 ;
	    RECT 18.4000 29.2000 18.8000 29.9000 ;
	    RECT 15.0000 28.8000 15.6000 29.2000 ;
	    RECT 18.2000 28.8000 18.8000 29.2000 ;
	    RECT 11.9000 27.3000 13.0000 27.6000 ;
	    RECT 9.0000 25.8000 9.8000 26.2000 ;
	    RECT 7.8000 24.8000 8.2000 25.2000 ;
	    RECT 7.9000 23.5000 8.2000 24.8000 ;
	    RECT 11.0000 25.1000 11.3000 26.2000 ;
	    RECT 11.9000 25.8000 12.2000 27.3000 ;
	    RECT 15.2000 27.1000 15.6000 28.8000 ;
	    RECT 18.4000 27.1000 18.8000 28.8000 ;
	    RECT 19.8000 27.6000 20.2000 29.9000 ;
	    RECT 19.8000 27.3000 20.9000 27.6000 ;
	    RECT 15.2000 26.9000 16.1000 27.1000 ;
	    RECT 18.4000 26.9000 19.3000 27.1000 ;
	    RECT 15.3000 26.8000 16.1000 26.9000 ;
	    RECT 18.5000 26.8000 19.3000 26.9000 ;
	    RECT 14.2000 25.8000 15.0000 26.2000 ;
	    RECT 11.6000 25.4000 12.2000 25.8000 ;
	    RECT 11.9000 25.1000 12.2000 25.4000 ;
	    RECT 15.8000 25.2000 16.1000 26.8000 ;
	    RECT 17.4000 25.8000 18.2000 26.2000 ;
	    RECT 19.0000 25.2000 19.3000 26.8000 ;
	    RECT 20.6000 25.8000 20.9000 27.3000 ;
	    RECT 21.4000 26.2000 21.8000 29.9000 ;
	    RECT 24.0000 27.1000 24.4000 29.9000 ;
	    RECT 25.4000 27.9000 25.8000 29.9000 ;
	    RECT 27.0000 28.9000 27.4000 29.9000 ;
	    RECT 24.0000 26.9000 24.9000 27.1000 ;
	    RECT 24.1000 26.8000 24.9000 26.9000 ;
	    RECT 20.6000 25.4000 21.2000 25.8000 ;
	    RECT 8.6000 23.8000 9.0000 24.6000 ;
	    RECT 7.9000 23.2000 9.7000 23.5000 ;
	    RECT 7.9000 23.1000 8.2000 23.2000 ;
	    RECT 7.8000 21.1000 8.2000 23.1000 ;
	    RECT 9.4000 23.1000 9.7000 23.2000 ;
	    RECT 9.4000 21.1000 9.8000 23.1000 ;
	    RECT 11.0000 21.1000 11.4000 25.1000 ;
	    RECT 11.9000 24.8000 13.0000 25.1000 ;
	    RECT 12.6000 21.1000 13.0000 24.8000 ;
	    RECT 15.8000 24.8000 16.2000 25.2000 ;
	    RECT 19.0000 24.8000 19.4000 25.2000 ;
	    RECT 20.6000 25.1000 20.9000 25.4000 ;
	    RECT 21.5000 25.1000 21.8000 26.2000 ;
	    RECT 23.0000 25.8000 24.2000 26.2000 ;
	    RECT 19.8000 24.8000 20.9000 25.1000 ;
	    RECT 15.0000 23.8000 15.4000 24.6000 ;
	    RECT 15.8000 23.5000 16.1000 24.8000 ;
	    RECT 18.2000 23.8000 18.6000 24.6000 ;
	    RECT 19.0000 23.5000 19.3000 24.8000 ;
	    RECT 14.3000 23.2000 16.1000 23.5000 ;
	    RECT 14.3000 23.1000 14.6000 23.2000 ;
	    RECT 14.2000 21.1000 14.6000 23.1000 ;
	    RECT 15.8000 23.1000 16.1000 23.2000 ;
	    RECT 17.5000 23.2000 19.3000 23.5000 ;
	    RECT 17.5000 23.1000 17.8000 23.2000 ;
	    RECT 15.8000 21.1000 16.2000 23.1000 ;
	    RECT 17.4000 21.1000 17.8000 23.1000 ;
	    RECT 19.0000 23.1000 19.3000 23.2000 ;
	    RECT 19.0000 21.1000 19.4000 23.1000 ;
	    RECT 19.8000 21.1000 20.2000 24.8000 ;
	    RECT 21.4000 21.1000 21.8000 25.1000 ;
	    RECT 22.2000 24.8000 22.6000 25.6000 ;
	    RECT 24.6000 25.2000 24.9000 26.8000 ;
	    RECT 25.4000 26.2000 25.7000 27.9000 ;
	    RECT 27.0000 27.8000 27.3000 28.9000 ;
	    RECT 27.8000 27.8000 28.2000 28.6000 ;
	    RECT 26.1000 27.5000 27.3000 27.8000 ;
	    RECT 28.6000 27.6000 29.0000 29.9000 ;
	    RECT 25.4000 25.8000 25.8000 26.2000 ;
	    RECT 26.1000 26.0000 26.4000 27.5000 ;
	    RECT 28.6000 27.3000 29.7000 27.6000 ;
	    RECT 24.6000 24.8000 25.0000 25.2000 ;
	    RECT 25.4000 25.1000 25.7000 25.8000 ;
	    RECT 26.1000 25.7000 26.5000 26.0000 ;
	    RECT 29.4000 25.8000 29.7000 27.3000 ;
	    RECT 30.2000 27.1000 30.6000 29.9000 ;
	    RECT 32.3000 28.2000 32.7000 29.9000 ;
	    RECT 31.8000 27.9000 32.7000 28.2000 ;
	    RECT 31.0000 27.1000 31.4000 27.6000 ;
	    RECT 30.2000 26.8000 31.4000 27.1000 ;
	    RECT 30.2000 26.2000 30.6000 26.8000 ;
	    RECT 26.1000 25.6000 28.2000 25.7000 ;
	    RECT 26.2000 25.4000 28.2000 25.6000 ;
	    RECT 25.4000 24.8000 26.1000 25.1000 ;
	    RECT 23.0000 24.1000 23.4000 24.2000 ;
	    RECT 23.8000 24.1000 24.2000 24.6000 ;
	    RECT 23.0000 23.8000 24.2000 24.1000 ;
	    RECT 24.6000 23.5000 24.9000 24.8000 ;
	    RECT 23.1000 23.2000 24.9000 23.5000 ;
	    RECT 23.0000 21.1000 23.4000 23.2000 ;
	    RECT 24.6000 23.1000 24.9000 23.2000 ;
	    RECT 24.6000 21.1000 25.0000 23.1000 ;
	    RECT 25.7000 21.1000 26.1000 24.8000 ;
	    RECT 27.8000 21.1000 28.2000 25.4000 ;
	    RECT 29.4000 25.4000 30.0000 25.8000 ;
	    RECT 29.4000 25.1000 29.7000 25.4000 ;
	    RECT 30.3000 25.1000 30.6000 26.2000 ;
	    RECT 28.6000 24.8000 29.7000 25.1000 ;
	    RECT 28.6000 21.1000 29.0000 24.8000 ;
	    RECT 30.2000 21.1000 30.6000 25.1000 ;
	    RECT 31.0000 24.8000 31.4000 25.2000 ;
	    RECT 31.0000 24.1000 31.3000 24.8000 ;
	    RECT 31.8000 24.1000 32.2000 27.9000 ;
	    RECT 35.2000 27.1000 35.6000 29.9000 ;
	    RECT 36.6000 27.9000 37.0000 29.9000 ;
	    RECT 38.2000 28.9000 38.6000 29.9000 ;
	    RECT 35.2000 26.9000 36.1000 27.1000 ;
	    RECT 35.3000 26.8000 36.1000 26.9000 ;
	    RECT 34.2000 25.8000 35.0000 26.2000 ;
	    RECT 32.6000 24.4000 33.0000 25.2000 ;
	    RECT 33.4000 24.8000 33.8000 25.6000 ;
	    RECT 35.8000 25.2000 36.1000 26.8000 ;
	    RECT 36.6000 26.2000 36.9000 27.9000 ;
	    RECT 38.2000 27.8000 38.5000 28.9000 ;
	    RECT 39.0000 27.8000 39.4000 28.6000 ;
	    RECT 37.3000 27.5000 38.5000 27.8000 ;
	    RECT 36.6000 25.8000 37.0000 26.2000 ;
	    RECT 37.3000 26.0000 37.6000 27.5000 ;
	    RECT 35.8000 24.8000 36.2000 25.2000 ;
	    RECT 36.6000 25.1000 36.9000 25.8000 ;
	    RECT 37.3000 25.7000 37.7000 26.0000 ;
	    RECT 37.3000 25.6000 39.4000 25.7000 ;
	    RECT 37.4000 25.4000 39.4000 25.6000 ;
	    RECT 36.6000 24.8000 37.3000 25.1000 ;
	    RECT 31.0000 23.8000 32.2000 24.1000 ;
	    RECT 31.8000 21.1000 32.2000 23.8000 ;
	    RECT 34.2000 23.8000 34.6000 24.2000 ;
	    RECT 35.0000 23.8000 35.4000 24.6000 ;
	    RECT 34.2000 23.5000 34.5000 23.8000 ;
	    RECT 35.8000 23.5000 36.1000 24.8000 ;
	    RECT 34.2000 23.2000 36.1000 23.5000 ;
	    RECT 34.2000 21.1000 34.6000 23.2000 ;
	    RECT 35.8000 23.1000 36.1000 23.2000 ;
	    RECT 35.8000 21.1000 36.2000 23.1000 ;
	    RECT 36.9000 21.1000 37.3000 24.8000 ;
	    RECT 39.0000 21.1000 39.4000 25.4000 ;
	    RECT 39.8000 21.1000 40.2000 29.9000 ;
	    RECT 42.2000 25.1000 42.6000 29.9000 ;
	    RECT 43.3000 28.2000 43.7000 29.9000 ;
	    RECT 43.3000 27.9000 44.2000 28.2000 ;
	    RECT 43.0000 25.1000 43.4000 25.2000 ;
	    RECT 42.2000 24.8000 43.4000 25.1000 ;
	    RECT 42.2000 21.1000 42.6000 24.8000 ;
	    RECT 43.0000 24.4000 43.4000 24.8000 ;
	    RECT 43.8000 25.1000 44.2000 27.9000 ;
	    RECT 44.6000 26.8000 45.0000 27.6000 ;
	    RECT 44.6000 25.1000 45.0000 25.2000 ;
	    RECT 43.8000 24.8000 45.0000 25.1000 ;
	    RECT 46.2000 25.1000 46.6000 29.9000 ;
	    RECT 47.3000 29.2000 47.7000 29.9000 ;
	    RECT 47.0000 28.8000 47.7000 29.2000 ;
	    RECT 50.2000 28.9000 50.6000 29.9000 ;
	    RECT 47.3000 28.2000 47.7000 28.8000 ;
	    RECT 47.3000 27.9000 48.2000 28.2000 ;
	    RECT 47.0000 25.1000 47.4000 25.2000 ;
	    RECT 46.2000 24.8000 47.4000 25.1000 ;
	    RECT 43.8000 21.1000 44.2000 24.8000 ;
	    RECT 46.2000 21.1000 46.6000 24.8000 ;
	    RECT 47.0000 24.4000 47.4000 24.8000 ;
	    RECT 47.8000 21.1000 48.2000 27.9000 ;
	    RECT 49.4000 27.8000 49.8000 28.6000 ;
	    RECT 50.3000 27.8000 50.6000 28.9000 ;
	    RECT 51.8000 27.9000 52.2000 29.9000 ;
	    RECT 48.6000 27.1000 49.0000 27.6000 ;
	    RECT 49.4000 27.1000 49.7000 27.8000 ;
	    RECT 50.3000 27.5000 51.5000 27.8000 ;
	    RECT 48.6000 26.8000 49.7000 27.1000 ;
	    RECT 51.2000 26.0000 51.5000 27.5000 ;
	    RECT 51.9000 26.2000 52.2000 27.9000 ;
	    RECT 53.2000 27.1000 53.6000 29.9000 ;
	    RECT 56.4000 29.2000 56.8000 29.9000 ;
	    RECT 56.4000 28.8000 57.0000 29.2000 ;
	    RECT 56.4000 27.1000 56.8000 28.8000 ;
	    RECT 51.1000 25.7000 51.5000 26.0000 ;
	    RECT 51.8000 25.8000 52.2000 26.2000 ;
	    RECT 49.4000 25.6000 51.5000 25.7000 ;
	    RECT 49.4000 25.4000 51.4000 25.6000 ;
	    RECT 49.4000 21.1000 49.8000 25.4000 ;
	    RECT 51.9000 25.1000 52.2000 25.8000 ;
	    RECT 52.7000 26.9000 53.6000 27.1000 ;
	    RECT 55.9000 26.9000 56.8000 27.1000 ;
	    RECT 52.7000 26.8000 53.5000 26.9000 ;
	    RECT 55.9000 26.8000 56.7000 26.9000 ;
	    RECT 52.7000 25.2000 53.0000 26.8000 ;
	    RECT 53.8000 25.8000 54.6000 26.2000 ;
	    RECT 55.9000 25.2000 56.2000 26.8000 ;
	    RECT 59.0000 26.2000 59.4000 29.9000 ;
	    RECT 60.6000 27.6000 61.0000 29.9000 ;
	    RECT 63.3000 29.2000 63.7000 29.9000 ;
	    RECT 65.7000 29.2000 66.1000 29.9000 ;
	    RECT 63.3000 28.8000 64.2000 29.2000 ;
	    RECT 65.7000 28.8000 66.6000 29.2000 ;
	    RECT 63.3000 28.2000 63.7000 28.8000 ;
	    RECT 65.7000 28.2000 66.1000 28.8000 ;
	    RECT 63.3000 27.9000 64.2000 28.2000 ;
	    RECT 65.7000 27.9000 66.6000 28.2000 ;
	    RECT 59.9000 27.3000 61.0000 27.6000 ;
	    RECT 57.0000 25.8000 57.8000 26.2000 ;
	    RECT 51.5000 24.8000 52.2000 25.1000 ;
	    RECT 52.6000 24.8000 53.0000 25.2000 ;
	    RECT 55.8000 24.8000 56.2000 25.2000 ;
	    RECT 51.5000 21.1000 51.9000 24.8000 ;
	    RECT 52.7000 23.5000 53.0000 24.8000 ;
	    RECT 53.4000 23.8000 53.8000 24.6000 ;
	    RECT 54.2000 23.8000 54.6000 24.2000 ;
	    RECT 54.2000 23.5000 54.5000 23.8000 ;
	    RECT 52.7000 23.2000 54.5000 23.5000 ;
	    RECT 52.7000 23.1000 53.0000 23.2000 ;
	    RECT 52.6000 21.1000 53.0000 23.1000 ;
	    RECT 54.2000 23.1000 54.5000 23.2000 ;
	    RECT 55.9000 23.5000 56.2000 24.8000 ;
	    RECT 59.0000 25.1000 59.3000 26.2000 ;
	    RECT 59.9000 25.8000 60.2000 27.3000 ;
	    RECT 59.6000 25.4000 60.2000 25.8000 ;
	    RECT 59.9000 25.1000 60.2000 25.4000 ;
	    RECT 61.4000 25.1000 61.8000 25.2000 ;
	    RECT 63.0000 25.1000 63.4000 25.2000 ;
	    RECT 56.6000 23.8000 57.0000 24.6000 ;
	    RECT 55.9000 23.2000 57.7000 23.5000 ;
	    RECT 55.9000 23.1000 56.2000 23.2000 ;
	    RECT 54.2000 21.1000 54.6000 23.1000 ;
	    RECT 55.8000 21.1000 56.2000 23.1000 ;
	    RECT 57.4000 23.1000 57.7000 23.2000 ;
	    RECT 57.4000 21.1000 57.8000 23.1000 ;
	    RECT 59.0000 21.1000 59.4000 25.1000 ;
	    RECT 59.9000 24.8000 61.0000 25.1000 ;
	    RECT 61.4000 24.8000 63.4000 25.1000 ;
	    RECT 60.6000 21.1000 61.0000 24.8000 ;
	    RECT 63.0000 24.4000 63.4000 24.8000 ;
	    RECT 63.8000 21.1000 64.2000 27.9000 ;
	    RECT 65.4000 24.4000 65.8000 25.2000 ;
	    RECT 66.2000 21.1000 66.6000 27.9000 ;
	    RECT 67.8000 26.2000 68.2000 29.9000 ;
	    RECT 69.4000 27.6000 69.8000 29.9000 ;
	    RECT 71.0000 28.9000 71.4000 29.9000 ;
	    RECT 70.2000 27.8000 70.6000 28.6000 ;
	    RECT 71.1000 27.8000 71.4000 28.9000 ;
	    RECT 72.6000 27.9000 73.0000 29.9000 ;
	    RECT 75.2000 29.2000 75.6000 29.9000 ;
	    RECT 76.9000 29.2000 77.3000 29.9000 ;
	    RECT 75.0000 28.8000 75.6000 29.2000 ;
	    RECT 76.6000 28.8000 77.3000 29.2000 ;
	    RECT 68.7000 27.3000 69.8000 27.6000 ;
	    RECT 71.1000 27.5000 72.3000 27.8000 ;
	    RECT 67.8000 25.1000 68.1000 26.2000 ;
	    RECT 68.7000 25.8000 69.0000 27.3000 ;
	    RECT 72.0000 26.0000 72.3000 27.5000 ;
	    RECT 72.7000 26.2000 73.0000 27.9000 ;
	    RECT 75.2000 27.1000 75.6000 28.8000 ;
	    RECT 76.9000 28.2000 77.3000 28.8000 ;
	    RECT 76.9000 27.9000 77.8000 28.2000 ;
	    RECT 75.2000 26.9000 76.1000 27.1000 ;
	    RECT 75.3000 26.8000 76.1000 26.9000 ;
	    RECT 68.4000 25.4000 69.0000 25.8000 ;
	    RECT 71.9000 25.7000 72.3000 26.0000 ;
	    RECT 72.6000 25.8000 73.0000 26.2000 ;
	    RECT 74.2000 25.8000 75.0000 26.2000 ;
	    RECT 68.7000 25.1000 69.0000 25.4000 ;
	    RECT 70.2000 25.6000 72.3000 25.7000 ;
	    RECT 70.2000 25.4000 72.2000 25.6000 ;
	    RECT 67.8000 21.1000 68.2000 25.1000 ;
	    RECT 68.7000 24.8000 69.8000 25.1000 ;
	    RECT 69.4000 21.1000 69.8000 24.8000 ;
	    RECT 70.2000 21.1000 70.6000 25.4000 ;
	    RECT 72.7000 25.1000 73.0000 25.8000 ;
	    RECT 72.3000 24.8000 73.0000 25.1000 ;
	    RECT 73.4000 24.8000 73.8000 25.6000 ;
	    RECT 75.8000 25.2000 76.1000 26.8000 ;
	    RECT 75.8000 24.8000 76.2000 25.2000 ;
	    RECT 72.3000 24.1000 72.7000 24.8000 ;
	    RECT 74.2000 24.1000 74.6000 24.2000 ;
	    RECT 72.3000 23.8000 74.6000 24.1000 ;
	    RECT 75.0000 23.8000 75.4000 24.6000 ;
	    RECT 72.3000 21.1000 72.7000 23.8000 ;
	    RECT 75.8000 23.5000 76.1000 24.8000 ;
	    RECT 76.6000 24.4000 77.0000 25.2000 ;
	    RECT 74.3000 23.2000 76.1000 23.5000 ;
	    RECT 74.3000 23.1000 74.6000 23.2000 ;
	    RECT 74.2000 21.1000 74.6000 23.1000 ;
	    RECT 75.8000 23.1000 76.1000 23.2000 ;
	    RECT 75.8000 21.1000 76.2000 23.1000 ;
	    RECT 77.4000 21.1000 77.8000 27.9000 ;
	    RECT 79.0000 26.2000 79.4000 29.9000 ;
	    RECT 80.6000 27.6000 81.0000 29.9000 ;
	    RECT 82.2000 29.1000 82.6000 29.2000 ;
	    RECT 83.2000 29.1000 83.6000 29.9000 ;
	    RECT 82.2000 28.8000 83.6000 29.1000 ;
	    RECT 85.4000 28.9000 85.8000 29.9000 ;
	    RECT 79.9000 27.3000 81.0000 27.6000 ;
	    RECT 79.0000 25.1000 79.3000 26.2000 ;
	    RECT 79.9000 25.8000 80.2000 27.3000 ;
	    RECT 83.2000 27.1000 83.6000 28.8000 ;
	    RECT 84.6000 27.8000 85.0000 28.6000 ;
	    RECT 85.5000 27.8000 85.8000 28.9000 ;
	    RECT 87.0000 27.9000 87.4000 29.9000 ;
	    RECT 85.5000 27.5000 86.7000 27.8000 ;
	    RECT 83.2000 26.9000 84.1000 27.1000 ;
	    RECT 83.3000 26.8000 84.1000 26.9000 ;
	    RECT 82.2000 25.8000 83.0000 26.2000 ;
	    RECT 79.6000 25.4000 80.2000 25.8000 ;
	    RECT 79.9000 25.1000 80.2000 25.4000 ;
	    RECT 83.8000 25.2000 84.1000 26.8000 ;
	    RECT 86.4000 26.0000 86.7000 27.5000 ;
	    RECT 87.1000 26.2000 87.4000 27.9000 ;
	    RECT 86.3000 25.7000 86.7000 26.0000 ;
	    RECT 87.0000 25.8000 87.4000 26.2000 ;
	    RECT 84.6000 25.6000 86.7000 25.7000 ;
	    RECT 84.6000 25.4000 86.6000 25.6000 ;
	    RECT 79.0000 21.1000 79.4000 25.1000 ;
	    RECT 79.9000 24.8000 81.0000 25.1000 ;
	    RECT 80.6000 21.1000 81.0000 24.8000 ;
	    RECT 83.8000 24.8000 84.2000 25.2000 ;
	    RECT 83.0000 23.8000 83.4000 24.6000 ;
	    RECT 83.8000 23.5000 84.1000 24.8000 ;
	    RECT 82.3000 23.2000 84.1000 23.5000 ;
	    RECT 82.3000 23.1000 82.6000 23.2000 ;
	    RECT 82.2000 21.1000 82.6000 23.1000 ;
	    RECT 83.8000 23.1000 84.1000 23.2000 ;
	    RECT 83.8000 21.1000 84.2000 23.1000 ;
	    RECT 84.6000 21.1000 85.0000 25.4000 ;
	    RECT 87.1000 25.2000 87.4000 25.8000 ;
	    RECT 87.0000 25.1000 87.4000 25.2000 ;
	    RECT 86.7000 24.8000 87.4000 25.1000 ;
	    RECT 86.7000 21.1000 87.1000 24.8000 ;
	    RECT 88.6000 21.1000 89.0000 29.9000 ;
	    RECT 90.7000 28.2000 91.1000 29.9000 ;
	    RECT 90.2000 27.9000 91.1000 28.2000 ;
	    RECT 89.4000 26.8000 89.8000 27.6000 ;
	    RECT 90.2000 21.1000 90.6000 27.9000 ;
	    RECT 91.0000 25.1000 91.4000 25.2000 ;
	    RECT 91.8000 25.1000 92.2000 29.9000 ;
	    RECT 94.0000 27.1000 94.4000 29.9000 ;
	    RECT 97.2000 29.1000 97.6000 29.9000 ;
	    RECT 101.6000 29.2000 102.0000 29.9000 ;
	    RECT 98.2000 29.1000 98.6000 29.2000 ;
	    RECT 97.2000 28.8000 98.6000 29.1000 ;
	    RECT 101.4000 28.8000 102.0000 29.2000 ;
	    RECT 95.0000 27.8000 95.4000 28.2000 ;
	    RECT 95.0000 27.1000 95.3000 27.8000 ;
	    RECT 97.2000 27.1000 97.6000 28.8000 ;
	    RECT 93.5000 26.8000 95.3000 27.1000 ;
	    RECT 96.7000 26.9000 97.6000 27.1000 ;
	    RECT 101.6000 27.1000 102.0000 28.8000 ;
	    RECT 101.6000 26.9000 102.5000 27.1000 ;
	    RECT 96.7000 26.8000 97.5000 26.9000 ;
	    RECT 101.7000 26.8000 102.5000 26.9000 ;
	    RECT 93.5000 25.2000 93.8000 26.8000 ;
	    RECT 94.6000 25.8000 95.4000 26.2000 ;
	    RECT 91.0000 24.8000 92.2000 25.1000 ;
	    RECT 93.4000 24.8000 93.8000 25.2000 ;
	    RECT 95.8000 24.8000 96.2000 25.6000 ;
	    RECT 96.7000 25.2000 97.0000 26.8000 ;
	    RECT 97.8000 25.8000 98.6000 26.2000 ;
	    RECT 100.6000 25.8000 101.4000 26.2000 ;
	    RECT 96.6000 24.8000 97.0000 25.2000 ;
	    RECT 91.0000 24.4000 91.4000 24.8000 ;
	    RECT 91.8000 21.1000 92.2000 24.8000 ;
	    RECT 93.5000 23.5000 93.8000 24.8000 ;
	    RECT 94.2000 23.8000 94.6000 24.6000 ;
	    RECT 96.7000 23.5000 97.0000 24.8000 ;
	    RECT 102.2000 25.2000 102.5000 26.8000 ;
	    RECT 102.2000 24.8000 102.6000 25.2000 ;
	    RECT 103.8000 25.1000 104.2000 29.9000 ;
	    RECT 104.9000 29.2000 105.3000 29.9000 ;
	    RECT 104.9000 28.8000 105.8000 29.2000 ;
	    RECT 107.8000 29.1000 108.2000 29.2000 ;
	    RECT 108.8000 29.1000 109.2000 29.9000 ;
	    RECT 107.8000 28.8000 109.2000 29.1000 ;
	    RECT 104.9000 28.2000 105.3000 28.8000 ;
	    RECT 104.9000 27.9000 105.8000 28.2000 ;
	    RECT 104.6000 25.1000 105.0000 25.2000 ;
	    RECT 103.8000 24.8000 105.0000 25.1000 ;
	    RECT 97.4000 24.1000 97.8000 24.6000 ;
	    RECT 99.8000 24.1000 100.2000 24.2000 ;
	    RECT 97.4000 23.8000 100.2000 24.1000 ;
	    RECT 101.4000 23.8000 101.8000 24.6000 ;
	    RECT 102.2000 23.5000 102.5000 24.8000 ;
	    RECT 93.5000 23.2000 95.3000 23.5000 ;
	    RECT 93.5000 23.1000 93.8000 23.2000 ;
	    RECT 93.4000 21.1000 93.8000 23.1000 ;
	    RECT 95.0000 23.1000 95.3000 23.2000 ;
	    RECT 96.7000 23.2000 98.5000 23.5000 ;
	    RECT 96.7000 23.1000 97.0000 23.2000 ;
	    RECT 95.0000 21.1000 95.4000 23.1000 ;
	    RECT 96.6000 21.1000 97.0000 23.1000 ;
	    RECT 98.2000 23.1000 98.5000 23.2000 ;
	    RECT 100.7000 23.2000 102.5000 23.5000 ;
	    RECT 100.7000 23.1000 101.0000 23.2000 ;
	    RECT 98.2000 21.1000 98.6000 23.1000 ;
	    RECT 100.6000 21.1000 101.0000 23.1000 ;
	    RECT 102.2000 23.1000 102.5000 23.2000 ;
	    RECT 102.2000 21.1000 102.6000 23.1000 ;
	    RECT 103.8000 21.1000 104.2000 24.8000 ;
	    RECT 104.6000 24.4000 105.0000 24.8000 ;
	    RECT 105.4000 21.1000 105.8000 27.9000 ;
	    RECT 106.2000 26.8000 106.6000 27.6000 ;
	    RECT 108.8000 27.1000 109.2000 28.8000 ;
	    RECT 108.8000 26.9000 109.7000 27.1000 ;
	    RECT 108.9000 26.8000 109.7000 26.9000 ;
	    RECT 107.8000 25.8000 109.0000 26.2000 ;
	    RECT 109.4000 25.2000 109.7000 26.8000 ;
	    RECT 110.2000 26.2000 110.6000 29.9000 ;
	    RECT 111.8000 27.6000 112.2000 29.9000 ;
	    RECT 114.5000 28.2000 114.9000 29.9000 ;
	    RECT 116.9000 29.2000 117.3000 29.9000 ;
	    RECT 116.9000 28.8000 117.8000 29.2000 ;
	    RECT 119.8000 28.9000 120.2000 29.9000 ;
	    RECT 116.9000 28.2000 117.3000 28.8000 ;
	    RECT 114.5000 27.9000 115.4000 28.2000 ;
	    RECT 116.9000 27.9000 117.8000 28.2000 ;
	    RECT 111.1000 27.3000 112.2000 27.6000 ;
	    RECT 109.4000 24.8000 109.8000 25.2000 ;
	    RECT 110.2000 25.1000 110.5000 26.2000 ;
	    RECT 111.1000 25.8000 111.4000 27.3000 ;
	    RECT 110.8000 25.4000 111.4000 25.8000 ;
	    RECT 111.1000 25.1000 111.4000 25.4000 ;
	    RECT 108.6000 23.8000 109.0000 24.6000 ;
	    RECT 109.4000 23.5000 109.7000 24.8000 ;
	    RECT 107.9000 23.2000 109.7000 23.5000 ;
	    RECT 107.9000 23.1000 108.2000 23.2000 ;
	    RECT 107.8000 21.1000 108.2000 23.1000 ;
	    RECT 109.4000 23.1000 109.7000 23.2000 ;
	    RECT 109.4000 21.1000 109.8000 23.1000 ;
	    RECT 110.2000 21.1000 110.6000 25.1000 ;
	    RECT 111.1000 24.8000 112.2000 25.1000 ;
	    RECT 111.8000 21.1000 112.2000 24.8000 ;
	    RECT 114.2000 24.4000 114.6000 25.2000 ;
	    RECT 115.0000 25.1000 115.4000 27.9000 ;
	    RECT 115.8000 26.8000 116.2000 27.6000 ;
	    RECT 115.8000 25.8000 116.2000 26.2000 ;
	    RECT 115.8000 25.1000 116.1000 25.8000 ;
	    RECT 115.0000 24.8000 116.1000 25.1000 ;
	    RECT 115.0000 21.1000 115.4000 24.8000 ;
	    RECT 116.6000 24.4000 117.0000 25.2000 ;
	    RECT 117.4000 21.1000 117.8000 27.9000 ;
	    RECT 119.0000 27.8000 119.4000 28.6000 ;
	    RECT 119.9000 27.8000 120.2000 28.9000 ;
	    RECT 121.4000 27.9000 121.8000 29.9000 ;
	    RECT 119.9000 27.5000 121.1000 27.8000 ;
	    RECT 120.8000 26.0000 121.1000 27.5000 ;
	    RECT 121.5000 26.2000 121.8000 27.9000 ;
	    RECT 122.8000 27.1000 123.2000 29.9000 ;
	    RECT 126.7000 29.2000 127.1000 29.9000 ;
	    RECT 126.2000 28.8000 127.1000 29.2000 ;
	    RECT 128.6000 28.9000 129.0000 29.9000 ;
	    RECT 126.7000 28.2000 127.1000 28.8000 ;
	    RECT 120.7000 25.7000 121.1000 26.0000 ;
	    RECT 121.4000 25.8000 121.8000 26.2000 ;
	    RECT 119.0000 25.6000 121.1000 25.7000 ;
	    RECT 119.0000 25.4000 121.0000 25.6000 ;
	    RECT 119.0000 21.1000 119.4000 25.4000 ;
	    RECT 121.5000 25.1000 121.8000 25.8000 ;
	    RECT 122.3000 26.9000 123.2000 27.1000 ;
	    RECT 126.2000 27.9000 127.1000 28.2000 ;
	    RECT 122.3000 26.8000 123.1000 26.9000 ;
	    RECT 122.3000 25.2000 122.6000 26.8000 ;
	    RECT 123.4000 25.8000 124.2000 26.2000 ;
	    RECT 121.1000 24.8000 121.8000 25.1000 ;
	    RECT 122.2000 24.8000 122.6000 25.2000 ;
	    RECT 121.1000 21.1000 121.5000 24.8000 ;
	    RECT 122.3000 23.5000 122.6000 24.8000 ;
	    RECT 123.0000 23.8000 123.4000 24.6000 ;
	    RECT 122.3000 23.2000 124.1000 23.5000 ;
	    RECT 122.3000 23.1000 122.6000 23.2000 ;
	    RECT 122.2000 21.1000 122.6000 23.1000 ;
	    RECT 123.8000 21.1000 124.2000 23.2000 ;
	    RECT 126.2000 21.1000 126.6000 27.9000 ;
	    RECT 127.8000 27.8000 128.2000 28.6000 ;
	    RECT 128.7000 27.8000 129.0000 28.9000 ;
	    RECT 130.2000 27.9000 130.6000 29.9000 ;
	    RECT 128.7000 27.5000 129.9000 27.8000 ;
	    RECT 129.6000 26.0000 129.9000 27.5000 ;
	    RECT 130.3000 26.2000 130.6000 27.9000 ;
	    RECT 131.6000 27.1000 132.0000 29.9000 ;
	    RECT 129.5000 25.7000 129.9000 26.0000 ;
	    RECT 130.2000 25.8000 130.6000 26.2000 ;
	    RECT 127.8000 25.6000 129.9000 25.7000 ;
	    RECT 127.8000 25.4000 129.8000 25.6000 ;
	    RECT 127.0000 24.4000 127.4000 25.2000 ;
	    RECT 127.8000 21.1000 128.2000 25.4000 ;
	    RECT 130.3000 25.1000 130.6000 25.8000 ;
	    RECT 131.1000 26.9000 132.0000 27.1000 ;
	    RECT 136.0000 29.2000 136.4000 29.9000 ;
	    RECT 138.7000 29.2000 139.1000 29.9000 ;
	    RECT 136.0000 28.8000 137.0000 29.2000 ;
	    RECT 138.2000 28.8000 139.1000 29.2000 ;
	    RECT 140.6000 28.9000 141.0000 29.9000 ;
	    RECT 136.0000 27.1000 136.4000 28.8000 ;
	    RECT 138.7000 28.2000 139.1000 28.8000 ;
	    RECT 138.2000 27.9000 139.1000 28.2000 ;
	    RECT 136.0000 26.9000 136.9000 27.1000 ;
	    RECT 131.1000 26.8000 131.9000 26.9000 ;
	    RECT 136.1000 26.8000 136.9000 26.9000 ;
	    RECT 131.1000 25.2000 131.4000 26.8000 ;
	    RECT 132.2000 25.8000 133.0000 26.2000 ;
	    RECT 135.0000 25.8000 135.8000 26.2000 ;
	    RECT 129.9000 24.8000 130.6000 25.1000 ;
	    RECT 131.0000 24.8000 131.4000 25.2000 ;
	    RECT 133.4000 24.8000 133.8000 25.6000 ;
	    RECT 136.6000 25.2000 136.9000 26.8000 ;
	    RECT 136.6000 24.8000 137.0000 25.2000 ;
	    RECT 129.9000 21.1000 130.3000 24.8000 ;
	    RECT 131.1000 23.5000 131.4000 24.8000 ;
	    RECT 131.8000 23.8000 132.2000 24.6000 ;
	    RECT 135.8000 23.8000 136.2000 24.6000 ;
	    RECT 136.6000 23.5000 136.9000 24.8000 ;
	    RECT 131.1000 23.2000 132.9000 23.5000 ;
	    RECT 135.1000 23.2000 136.9000 23.5000 ;
	    RECT 131.1000 23.1000 131.4000 23.2000 ;
	    RECT 131.0000 21.1000 131.4000 23.1000 ;
	    RECT 132.6000 21.1000 133.0000 23.2000 ;
	    RECT 135.1000 23.1000 135.4000 23.2000 ;
	    RECT 135.0000 21.1000 135.4000 23.1000 ;
	    RECT 136.6000 23.1000 136.9000 23.2000 ;
	    RECT 136.6000 21.1000 137.0000 23.1000 ;
	    RECT 138.2000 21.1000 138.6000 27.9000 ;
	    RECT 139.8000 27.8000 140.2000 28.6000 ;
	    RECT 140.7000 27.8000 141.0000 28.9000 ;
	    RECT 142.2000 27.9000 142.6000 29.9000 ;
	    RECT 140.7000 27.5000 141.9000 27.8000 ;
	    RECT 141.6000 26.0000 141.9000 27.5000 ;
	    RECT 142.3000 26.2000 142.6000 27.9000 ;
	    RECT 143.6000 29.2000 144.0000 29.9000 ;
	    RECT 143.6000 28.8000 144.2000 29.2000 ;
	    RECT 143.6000 27.1000 144.0000 28.8000 ;
	    RECT 141.5000 25.7000 141.9000 26.0000 ;
	    RECT 142.2000 25.8000 142.6000 26.2000 ;
	    RECT 139.8000 25.6000 141.9000 25.7000 ;
	    RECT 139.8000 25.4000 141.8000 25.6000 ;
	    RECT 139.0000 24.4000 139.4000 25.2000 ;
	    RECT 139.8000 21.1000 140.2000 25.4000 ;
	    RECT 142.3000 25.1000 142.6000 25.8000 ;
	    RECT 143.1000 26.9000 144.0000 27.1000 ;
	    RECT 143.1000 26.8000 143.9000 26.9000 ;
	    RECT 143.1000 25.2000 143.4000 26.8000 ;
	    RECT 144.2000 25.8000 145.0000 26.2000 ;
	    RECT 147.0000 26.1000 147.4000 29.9000 ;
	    RECT 149.9000 29.2000 150.3000 29.9000 ;
	    RECT 149.4000 28.8000 150.3000 29.2000 ;
	    RECT 151.8000 29.1000 152.2000 29.2000 ;
	    RECT 152.8000 29.1000 153.2000 29.9000 ;
	    RECT 155.5000 29.2000 155.9000 29.9000 ;
	    RECT 151.8000 28.8000 153.2000 29.1000 ;
	    RECT 155.0000 28.8000 155.9000 29.2000 ;
	    RECT 149.9000 28.2000 150.3000 28.8000 ;
	    RECT 145.4000 25.8000 147.4000 26.1000 ;
	    RECT 141.9000 24.8000 142.6000 25.1000 ;
	    RECT 143.0000 24.8000 143.4000 25.2000 ;
	    RECT 145.4000 24.8000 145.8000 25.8000 ;
	    RECT 141.9000 21.1000 142.3000 24.8000 ;
	    RECT 143.1000 23.5000 143.4000 24.8000 ;
	    RECT 143.8000 24.1000 144.2000 24.6000 ;
	    RECT 144.6000 24.1000 145.0000 24.2000 ;
	    RECT 143.8000 23.8000 145.0000 24.1000 ;
	    RECT 143.1000 23.2000 144.9000 23.5000 ;
	    RECT 143.1000 23.1000 143.4000 23.2000 ;
	    RECT 143.0000 21.1000 143.4000 23.1000 ;
	    RECT 144.6000 23.1000 144.9000 23.2000 ;
	    RECT 144.6000 21.1000 145.0000 23.1000 ;
	    RECT 147.0000 21.1000 147.4000 25.8000 ;
	    RECT 149.4000 27.9000 150.3000 28.2000 ;
	    RECT 149.4000 21.1000 149.8000 27.9000 ;
	    RECT 152.8000 27.1000 153.2000 28.8000 ;
	    RECT 155.5000 28.2000 155.9000 28.8000 ;
	    RECT 155.0000 27.9000 155.9000 28.2000 ;
	    RECT 152.8000 26.9000 153.7000 27.1000 ;
	    RECT 152.9000 26.8000 153.7000 26.9000 ;
	    RECT 151.8000 25.8000 152.6000 26.2000 ;
	    RECT 153.4000 25.2000 153.7000 26.8000 ;
	    RECT 150.2000 24.4000 150.6000 25.2000 ;
	    RECT 153.4000 24.8000 153.8000 25.2000 ;
	    RECT 152.6000 23.8000 153.0000 24.6000 ;
	    RECT 153.4000 23.5000 153.7000 24.8000 ;
	    RECT 151.9000 23.2000 153.7000 23.5000 ;
	    RECT 151.9000 23.1000 152.2000 23.2000 ;
	    RECT 151.8000 21.1000 152.2000 23.1000 ;
	    RECT 153.4000 23.1000 153.7000 23.2000 ;
	    RECT 153.4000 21.1000 153.8000 23.1000 ;
	    RECT 155.0000 21.1000 155.4000 27.9000 ;
	    RECT 156.6000 26.2000 157.0000 29.9000 ;
	    RECT 158.2000 27.6000 158.6000 29.9000 ;
	    RECT 157.5000 27.3000 158.6000 27.6000 ;
	    RECT 159.0000 27.5000 159.4000 29.9000 ;
	    RECT 161.2000 29.2000 161.6000 29.9000 ;
	    RECT 160.6000 28.9000 161.6000 29.2000 ;
	    RECT 163.4000 28.9000 163.8000 29.9000 ;
	    RECT 165.5000 29.2000 166.1000 29.9000 ;
	    RECT 165.4000 28.9000 166.1000 29.2000 ;
	    RECT 160.6000 28.5000 161.0000 28.9000 ;
	    RECT 163.4000 28.6000 163.7000 28.9000 ;
	    RECT 161.4000 28.2000 161.8000 28.6000 ;
	    RECT 162.3000 28.3000 163.7000 28.6000 ;
	    RECT 165.4000 28.5000 165.8000 28.9000 ;
	    RECT 162.3000 28.2000 162.7000 28.3000 ;
	    RECT 155.8000 24.4000 156.2000 25.2000 ;
	    RECT 156.6000 25.1000 156.9000 26.2000 ;
	    RECT 157.5000 25.8000 157.8000 27.3000 ;
	    RECT 161.5000 27.2000 161.8000 28.2000 ;
	    RECT 166.3000 27.7000 166.7000 27.8000 ;
	    RECT 167.8000 27.7000 168.2000 29.9000 ;
	    RECT 169.4000 28.9000 169.8000 29.9000 ;
	    RECT 168.6000 27.8000 169.0000 28.6000 ;
	    RECT 169.5000 27.8000 169.8000 28.9000 ;
	    RECT 171.0000 29.1000 171.4000 29.9000 ;
	    RECT 171.8000 29.1000 172.2000 29.2000 ;
	    RECT 171.0000 28.8000 172.2000 29.1000 ;
	    RECT 171.0000 27.9000 171.4000 28.8000 ;
	    RECT 166.3000 27.4000 168.2000 27.7000 ;
	    RECT 169.5000 27.5000 170.7000 27.8000 ;
	    RECT 159.4000 27.1000 160.2000 27.2000 ;
	    RECT 161.4000 27.1000 161.8000 27.2000 ;
	    RECT 164.3000 27.1000 164.7000 27.2000 ;
	    RECT 159.4000 26.8000 164.9000 27.1000 ;
	    RECT 160.9000 26.7000 161.3000 26.8000 ;
	    RECT 160.1000 26.2000 160.5000 26.3000 ;
	    RECT 160.1000 25.9000 162.6000 26.2000 ;
	    RECT 162.2000 25.8000 162.6000 25.9000 ;
	    RECT 157.2000 25.4000 157.8000 25.8000 ;
	    RECT 157.5000 25.1000 157.8000 25.4000 ;
	    RECT 159.0000 25.5000 161.8000 25.6000 ;
	    RECT 159.0000 25.4000 161.9000 25.5000 ;
	    RECT 159.0000 25.3000 163.9000 25.4000 ;
	    RECT 156.6000 21.1000 157.0000 25.1000 ;
	    RECT 157.5000 24.8000 158.6000 25.1000 ;
	    RECT 158.2000 21.1000 158.6000 24.8000 ;
	    RECT 159.0000 21.1000 159.4000 25.3000 ;
	    RECT 161.5000 25.1000 163.9000 25.3000 ;
	    RECT 160.6000 24.5000 163.3000 24.8000 ;
	    RECT 160.6000 24.4000 161.0000 24.5000 ;
	    RECT 162.9000 24.4000 163.3000 24.5000 ;
	    RECT 163.6000 24.5000 163.9000 25.1000 ;
	    RECT 164.6000 25.2000 164.9000 26.8000 ;
	    RECT 165.4000 26.4000 165.8000 26.5000 ;
	    RECT 165.4000 26.1000 167.3000 26.4000 ;
	    RECT 166.9000 26.0000 167.3000 26.1000 ;
	    RECT 166.1000 25.7000 166.5000 25.8000 ;
	    RECT 167.8000 25.7000 168.2000 27.4000 ;
	    RECT 170.4000 26.0000 170.7000 27.5000 ;
	    RECT 171.1000 26.2000 171.4000 27.9000 ;
	    RECT 170.3000 25.7000 170.7000 26.0000 ;
	    RECT 171.0000 25.8000 171.4000 26.2000 ;
	    RECT 166.1000 25.4000 168.2000 25.7000 ;
	    RECT 164.6000 24.9000 165.8000 25.2000 ;
	    RECT 164.3000 24.5000 164.7000 24.6000 ;
	    RECT 163.6000 24.2000 164.7000 24.5000 ;
	    RECT 165.5000 24.4000 165.8000 24.9000 ;
	    RECT 165.5000 24.0000 166.2000 24.4000 ;
	    RECT 162.3000 23.7000 162.7000 23.8000 ;
	    RECT 163.7000 23.7000 164.1000 23.8000 ;
	    RECT 160.6000 23.1000 161.0000 23.5000 ;
	    RECT 162.3000 23.4000 164.1000 23.7000 ;
	    RECT 163.4000 23.1000 163.7000 23.4000 ;
	    RECT 165.4000 23.1000 165.8000 23.5000 ;
	    RECT 160.6000 22.8000 161.6000 23.1000 ;
	    RECT 161.2000 21.1000 161.6000 22.8000 ;
	    RECT 163.4000 21.1000 163.8000 23.1000 ;
	    RECT 165.5000 21.1000 166.1000 23.1000 ;
	    RECT 167.8000 21.1000 168.2000 25.4000 ;
	    RECT 168.6000 25.6000 170.7000 25.7000 ;
	    RECT 168.6000 25.4000 170.6000 25.6000 ;
	    RECT 168.6000 21.1000 169.0000 25.4000 ;
	    RECT 171.1000 25.1000 171.4000 25.8000 ;
	    RECT 170.7000 24.8000 171.4000 25.1000 ;
	    RECT 170.7000 21.1000 171.1000 24.8000 ;
	    RECT 1.4000 11.1000 1.8000 19.9000 ;
	    RECT 3.0000 17.9000 3.4000 19.9000 ;
	    RECT 3.1000 17.8000 3.4000 17.9000 ;
	    RECT 4.6000 17.9000 5.0000 19.9000 ;
	    RECT 4.6000 17.8000 4.9000 17.9000 ;
	    RECT 3.1000 17.5000 4.9000 17.8000 ;
	    RECT 3.1000 16.2000 3.4000 17.5000 ;
	    RECT 3.8000 16.4000 4.2000 17.2000 ;
	    RECT 6.5000 16.2000 6.9000 19.9000 ;
	    RECT 3.0000 15.8000 3.4000 16.2000 ;
	    RECT 3.1000 14.2000 3.4000 15.8000 ;
	    RECT 5.4000 15.4000 5.8000 16.2000 ;
	    RECT 6.2000 15.9000 6.9000 16.2000 ;
	    RECT 6.2000 15.2000 6.5000 15.9000 ;
	    RECT 8.6000 15.6000 9.0000 19.9000 ;
	    RECT 9.4000 17.9000 9.8000 19.9000 ;
	    RECT 9.5000 17.8000 9.8000 17.9000 ;
	    RECT 11.0000 17.9000 11.4000 19.9000 ;
	    RECT 11.0000 17.8000 11.3000 17.9000 ;
	    RECT 9.5000 17.5000 11.3000 17.8000 ;
	    RECT 9.5000 16.2000 9.8000 17.5000 ;
	    RECT 10.2000 16.4000 10.6000 17.2000 ;
	    RECT 9.4000 15.8000 9.8000 16.2000 ;
	    RECT 7.0000 15.4000 9.0000 15.6000 ;
	    RECT 6.9000 15.3000 9.0000 15.4000 ;
	    RECT 4.2000 14.8000 5.0000 15.2000 ;
	    RECT 6.2000 14.8000 6.6000 15.2000 ;
	    RECT 6.9000 15.0000 7.3000 15.3000 ;
	    RECT 3.1000 14.1000 3.9000 14.2000 ;
	    RECT 3.1000 13.9000 4.9000 14.1000 ;
	    RECT 3.6000 13.8000 4.9000 13.9000 ;
	    RECT 3.6000 11.1000 4.0000 13.8000 ;
	    RECT 4.6000 13.2000 4.9000 13.8000 ;
	    RECT 4.6000 12.8000 5.0000 13.2000 ;
	    RECT 6.2000 13.1000 6.5000 14.8000 ;
	    RECT 6.9000 13.5000 7.2000 15.0000 ;
	    RECT 9.5000 14.2000 9.8000 15.8000 ;
	    RECT 11.8000 16.1000 12.2000 16.2000 ;
	    RECT 12.6000 16.1000 13.0000 19.9000 ;
	    RECT 15.0000 17.9000 15.4000 19.9000 ;
	    RECT 15.1000 17.8000 15.4000 17.9000 ;
	    RECT 16.6000 17.9000 17.0000 19.9000 ;
	    RECT 18.2000 17.9000 18.6000 19.9000 ;
	    RECT 16.6000 17.8000 16.9000 17.9000 ;
	    RECT 15.1000 17.5000 16.9000 17.8000 ;
	    RECT 18.3000 17.8000 18.6000 17.9000 ;
	    RECT 19.8000 17.9000 20.2000 19.9000 ;
	    RECT 19.8000 17.8000 20.1000 17.9000 ;
	    RECT 18.3000 17.5000 20.1000 17.8000 ;
	    RECT 15.8000 16.4000 16.2000 17.2000 ;
	    RECT 11.8000 15.8000 13.0000 16.1000 ;
	    RECT 11.8000 15.4000 12.2000 15.8000 ;
	    RECT 10.6000 14.8000 11.4000 15.2000 ;
	    RECT 9.5000 14.1000 10.3000 14.2000 ;
	    RECT 9.5000 13.9000 10.4000 14.1000 ;
	    RECT 6.9000 13.2000 8.1000 13.5000 ;
	    RECT 6.2000 11.1000 6.6000 13.1000 ;
	    RECT 7.8000 12.1000 8.1000 13.2000 ;
	    RECT 8.6000 12.4000 9.0000 13.2000 ;
	    RECT 7.8000 11.1000 8.2000 12.1000 ;
	    RECT 10.0000 11.1000 10.4000 13.9000 ;
	    RECT 12.6000 11.1000 13.0000 15.8000 ;
	    RECT 16.6000 16.2000 16.9000 17.5000 ;
	    RECT 19.0000 16.4000 19.4000 17.2000 ;
	    RECT 19.8000 16.2000 20.1000 17.5000 ;
	    RECT 16.6000 15.8000 17.0000 16.2000 ;
	    RECT 17.4000 16.1000 17.8000 16.2000 ;
	    RECT 18.2000 16.1000 18.6000 16.2000 ;
	    RECT 17.4000 15.8000 18.6000 16.1000 ;
	    RECT 19.8000 15.8000 20.2000 16.2000 ;
	    RECT 15.0000 14.8000 15.8000 15.2000 ;
	    RECT 16.6000 14.2000 16.9000 15.8000 ;
	    RECT 17.4000 15.4000 17.8000 15.8000 ;
	    RECT 18.2000 14.8000 19.0000 15.2000 ;
	    RECT 19.8000 14.2000 20.1000 15.8000 ;
	    RECT 16.1000 14.1000 16.9000 14.2000 ;
	    RECT 19.3000 14.1000 20.1000 14.2000 ;
	    RECT 16.0000 13.9000 16.9000 14.1000 ;
	    RECT 19.2000 13.9000 20.1000 14.1000 ;
	    RECT 16.0000 11.1000 16.4000 13.9000 ;
	    RECT 19.2000 11.1000 19.6000 13.9000 ;
	    RECT 21.4000 13.1000 21.8000 19.9000 ;
	    RECT 23.8000 17.9000 24.2000 19.9000 ;
	    RECT 23.9000 17.8000 24.2000 17.9000 ;
	    RECT 25.4000 17.9000 25.8000 19.9000 ;
	    RECT 27.0000 17.9000 27.4000 19.9000 ;
	    RECT 25.4000 17.8000 25.7000 17.9000 ;
	    RECT 23.9000 17.5000 25.7000 17.8000 ;
	    RECT 27.1000 17.8000 27.4000 17.9000 ;
	    RECT 28.6000 17.9000 29.0000 19.9000 ;
	    RECT 28.6000 17.8000 28.9000 17.9000 ;
	    RECT 27.1000 17.5000 28.9000 17.8000 ;
	    RECT 22.2000 15.8000 22.6000 16.6000 ;
	    RECT 24.6000 16.4000 25.0000 17.2000 ;
	    RECT 25.4000 16.2000 25.7000 17.5000 ;
	    RECT 27.8000 16.4000 28.2000 17.2000 ;
	    RECT 28.6000 16.2000 28.9000 17.5000 ;
	    RECT 29.4000 16.2000 29.8000 19.9000 ;
	    RECT 25.4000 15.8000 25.8000 16.2000 ;
	    RECT 23.8000 14.8000 24.6000 15.2000 ;
	    RECT 25.4000 14.2000 25.7000 15.8000 ;
	    RECT 26.2000 15.4000 26.6000 16.2000 ;
	    RECT 28.6000 15.8000 29.0000 16.2000 ;
	    RECT 29.4000 15.9000 30.5000 16.2000 ;
	    RECT 31.0000 15.9000 31.4000 19.9000 ;
	    RECT 32.6000 17.9000 33.0000 19.9000 ;
	    RECT 32.7000 17.8000 33.0000 17.9000 ;
	    RECT 34.2000 17.9000 34.6000 19.9000 ;
	    RECT 34.2000 17.8000 34.5000 17.9000 ;
	    RECT 32.7000 17.5000 34.5000 17.8000 ;
	    RECT 33.4000 16.4000 33.8000 17.2000 ;
	    RECT 34.2000 16.2000 34.5000 17.5000 ;
	    RECT 35.3000 16.2000 35.7000 19.9000 ;
	    RECT 27.0000 14.8000 27.8000 15.2000 ;
	    RECT 28.6000 14.2000 28.9000 15.8000 ;
	    RECT 24.9000 14.1000 25.7000 14.2000 ;
	    RECT 28.1000 14.1000 28.9000 14.2000 ;
	    RECT 24.8000 13.9000 25.7000 14.1000 ;
	    RECT 28.0000 13.9000 28.9000 14.1000 ;
	    RECT 30.2000 15.6000 30.5000 15.9000 ;
	    RECT 30.2000 15.2000 30.8000 15.6000 ;
	    RECT 21.4000 12.8000 22.3000 13.1000 ;
	    RECT 21.9000 11.1000 22.3000 12.8000 ;
	    RECT 24.8000 11.1000 25.2000 13.9000 ;
	    RECT 28.0000 11.1000 28.4000 13.9000 ;
	    RECT 30.2000 13.7000 30.5000 15.2000 ;
	    RECT 31.1000 14.8000 31.4000 15.9000 ;
	    RECT 31.8000 15.4000 32.2000 16.2000 ;
	    RECT 34.2000 15.8000 34.6000 16.2000 ;
	    RECT 35.0000 15.9000 35.7000 16.2000 ;
	    RECT 32.6000 14.8000 33.4000 15.2000 ;
	    RECT 29.4000 13.4000 30.5000 13.7000 ;
	    RECT 29.4000 11.1000 29.8000 13.4000 ;
	    RECT 31.0000 11.1000 31.4000 14.8000 ;
	    RECT 34.2000 14.2000 34.5000 15.8000 ;
	    RECT 33.7000 14.1000 34.5000 14.2000 ;
	    RECT 33.6000 13.9000 34.5000 14.1000 ;
	    RECT 35.0000 15.2000 35.3000 15.9000 ;
	    RECT 37.4000 15.6000 37.8000 19.9000 ;
	    RECT 38.5000 16.2000 38.9000 19.9000 ;
	    RECT 35.8000 15.4000 37.8000 15.6000 ;
	    RECT 35.7000 15.3000 37.8000 15.4000 ;
	    RECT 38.2000 15.9000 38.9000 16.2000 ;
	    RECT 35.0000 14.8000 35.4000 15.2000 ;
	    RECT 35.7000 15.0000 36.1000 15.3000 ;
	    RECT 38.2000 15.2000 38.5000 15.9000 ;
	    RECT 40.6000 15.6000 41.0000 19.9000 ;
	    RECT 41.7000 16.2000 42.1000 19.9000 ;
	    RECT 39.0000 15.4000 41.0000 15.6000 ;
	    RECT 38.9000 15.3000 41.0000 15.4000 ;
	    RECT 41.4000 15.9000 42.1000 16.2000 ;
	    RECT 33.6000 11.1000 34.0000 13.9000 ;
	    RECT 35.0000 13.1000 35.3000 14.8000 ;
	    RECT 35.7000 13.5000 36.0000 15.0000 ;
	    RECT 38.2000 14.8000 38.6000 15.2000 ;
	    RECT 38.9000 15.0000 39.3000 15.3000 ;
	    RECT 41.4000 15.2000 41.7000 15.9000 ;
	    RECT 43.8000 15.6000 44.2000 19.9000 ;
	    RECT 45.9000 17.2000 46.3000 19.9000 ;
	    RECT 45.4000 16.8000 46.3000 17.2000 ;
	    RECT 46.6000 16.8000 47.0000 17.2000 ;
	    RECT 45.9000 16.2000 46.3000 16.8000 ;
	    RECT 46.7000 16.2000 47.0000 16.8000 ;
	    RECT 45.9000 15.9000 46.4000 16.2000 ;
	    RECT 46.7000 15.9000 47.4000 16.2000 ;
	    RECT 42.2000 15.4000 44.2000 15.6000 ;
	    RECT 42.1000 15.3000 44.2000 15.4000 ;
	    RECT 35.7000 13.2000 36.9000 13.5000 ;
	    RECT 35.0000 11.1000 35.4000 13.1000 ;
	    RECT 36.6000 12.1000 36.9000 13.2000 ;
	    RECT 37.4000 12.4000 37.8000 13.2000 ;
	    RECT 38.2000 13.1000 38.5000 14.8000 ;
	    RECT 38.9000 13.5000 39.2000 15.0000 ;
	    RECT 41.4000 14.8000 41.8000 15.2000 ;
	    RECT 42.1000 15.0000 42.5000 15.3000 ;
	    RECT 38.9000 13.2000 40.1000 13.5000 ;
	    RECT 36.6000 11.1000 37.0000 12.1000 ;
	    RECT 38.2000 11.1000 38.6000 13.1000 ;
	    RECT 39.8000 12.1000 40.1000 13.2000 ;
	    RECT 40.6000 12.4000 41.0000 13.2000 ;
	    RECT 41.4000 13.1000 41.7000 14.8000 ;
	    RECT 42.1000 13.5000 42.4000 15.0000 ;
	    RECT 45.4000 14.4000 45.8000 15.2000 ;
	    RECT 46.1000 14.2000 46.4000 15.9000 ;
	    RECT 47.0000 15.8000 47.4000 15.9000 ;
	    RECT 44.6000 14.1000 45.0000 14.2000 ;
	    RECT 44.6000 13.8000 45.4000 14.1000 ;
	    RECT 46.1000 13.8000 47.4000 14.2000 ;
	    RECT 45.0000 13.6000 45.4000 13.8000 ;
	    RECT 42.1000 13.2000 43.3000 13.5000 ;
	    RECT 39.8000 11.1000 40.2000 12.1000 ;
	    RECT 41.4000 11.1000 41.8000 13.1000 ;
	    RECT 43.0000 12.1000 43.3000 13.2000 ;
	    RECT 43.8000 12.4000 44.2000 13.2000 ;
	    RECT 44.7000 13.1000 46.5000 13.3000 ;
	    RECT 47.0000 13.1000 47.3000 13.8000 ;
	    RECT 44.6000 13.0000 46.6000 13.1000 ;
	    RECT 43.0000 11.1000 43.4000 12.1000 ;
	    RECT 44.6000 11.1000 45.0000 13.0000 ;
	    RECT 46.2000 11.1000 46.6000 13.0000 ;
	    RECT 47.0000 11.1000 47.4000 13.1000 ;
	    RECT 47.8000 11.1000 48.2000 19.9000 ;
	    RECT 49.4000 17.9000 49.8000 19.9000 ;
	    RECT 49.5000 17.8000 49.8000 17.9000 ;
	    RECT 51.0000 17.9000 51.4000 19.9000 ;
	    RECT 51.0000 17.8000 51.3000 17.9000 ;
	    RECT 49.5000 17.5000 51.3000 17.8000 ;
	    RECT 49.5000 16.2000 49.8000 17.5000 ;
	    RECT 50.2000 16.4000 50.6000 17.2000 ;
	    RECT 52.9000 16.2000 53.3000 19.9000 ;
	    RECT 49.4000 15.8000 49.8000 16.2000 ;
	    RECT 51.0000 16.1000 51.4000 16.2000 ;
	    RECT 51.8000 16.1000 52.2000 16.2000 ;
	    RECT 51.0000 15.8000 52.2000 16.1000 ;
	    RECT 49.5000 14.2000 49.8000 15.8000 ;
	    RECT 51.8000 15.4000 52.2000 15.8000 ;
	    RECT 52.6000 15.9000 53.3000 16.2000 ;
	    RECT 52.6000 15.2000 52.9000 15.9000 ;
	    RECT 55.0000 15.6000 55.4000 19.9000 ;
	    RECT 56.9000 19.2000 57.3000 19.9000 ;
	    RECT 56.9000 18.8000 57.8000 19.2000 ;
	    RECT 56.2000 16.8000 56.6000 17.2000 ;
	    RECT 56.2000 16.2000 56.5000 16.8000 ;
	    RECT 56.9000 16.2000 57.3000 18.8000 ;
	    RECT 55.8000 15.9000 56.5000 16.2000 ;
	    RECT 56.8000 15.9000 57.3000 16.2000 ;
	    RECT 55.8000 15.8000 56.2000 15.9000 ;
	    RECT 53.4000 15.4000 55.4000 15.6000 ;
	    RECT 53.3000 15.3000 55.4000 15.4000 ;
	    RECT 50.6000 14.8000 51.4000 15.2000 ;
	    RECT 52.6000 14.8000 53.0000 15.2000 ;
	    RECT 53.3000 15.0000 53.7000 15.3000 ;
	    RECT 49.5000 14.1000 50.3000 14.2000 ;
	    RECT 49.5000 13.9000 50.4000 14.1000 ;
	    RECT 50.0000 11.1000 50.4000 13.9000 ;
	    RECT 52.6000 13.1000 52.9000 14.8000 ;
	    RECT 53.3000 13.5000 53.6000 15.0000 ;
	    RECT 56.8000 14.2000 57.1000 15.9000 ;
	    RECT 57.4000 15.1000 57.8000 15.2000 ;
	    RECT 58.2000 15.1000 58.6000 15.2000 ;
	    RECT 57.4000 14.8000 58.6000 15.1000 ;
	    RECT 57.4000 14.4000 57.8000 14.8000 ;
	    RECT 55.8000 13.8000 57.1000 14.2000 ;
	    RECT 58.2000 14.1000 58.6000 14.2000 ;
	    RECT 59.0000 14.1000 59.4000 19.9000 ;
	    RECT 57.8000 13.8000 59.4000 14.1000 ;
	    RECT 53.3000 13.2000 54.5000 13.5000 ;
	    RECT 52.6000 11.1000 53.0000 13.1000 ;
	    RECT 54.2000 12.1000 54.5000 13.2000 ;
	    RECT 55.0000 12.4000 55.4000 13.2000 ;
	    RECT 55.9000 13.1000 56.2000 13.8000 ;
	    RECT 57.8000 13.6000 58.2000 13.8000 ;
	    RECT 56.7000 13.1000 58.5000 13.3000 ;
	    RECT 54.2000 11.1000 54.6000 12.1000 ;
	    RECT 55.8000 11.1000 56.2000 13.1000 ;
	    RECT 56.6000 13.0000 58.6000 13.1000 ;
	    RECT 56.6000 11.1000 57.0000 13.0000 ;
	    RECT 58.2000 11.1000 58.6000 13.0000 ;
	    RECT 59.0000 11.1000 59.4000 13.8000 ;
	    RECT 63.0000 14.1000 63.4000 19.9000 ;
	    RECT 65.1000 16.2000 65.5000 19.9000 ;
	    RECT 67.0000 17.9000 67.4000 19.9000 ;
	    RECT 67.1000 17.8000 67.4000 17.9000 ;
	    RECT 68.6000 17.9000 69.0000 19.9000 ;
	    RECT 68.6000 17.8000 68.9000 17.9000 ;
	    RECT 67.1000 17.5000 68.9000 17.8000 ;
	    RECT 65.8000 16.8000 66.2000 17.2000 ;
	    RECT 65.9000 16.2000 66.2000 16.8000 ;
	    RECT 67.1000 16.2000 67.4000 17.5000 ;
	    RECT 67.8000 16.4000 68.2000 17.2000 ;
	    RECT 65.1000 15.9000 65.6000 16.2000 ;
	    RECT 65.9000 15.9000 66.6000 16.2000 ;
	    RECT 65.3000 15.2000 65.6000 15.9000 ;
	    RECT 66.2000 15.8000 66.6000 15.9000 ;
	    RECT 67.0000 15.8000 67.4000 16.2000 ;
	    RECT 63.8000 15.1000 64.2000 15.2000 ;
	    RECT 64.6000 15.1000 65.0000 15.2000 ;
	    RECT 63.8000 14.8000 65.0000 15.1000 ;
	    RECT 64.6000 14.4000 65.0000 14.8000 ;
	    RECT 65.3000 14.8000 65.8000 15.2000 ;
	    RECT 65.3000 14.2000 65.6000 14.8000 ;
	    RECT 67.1000 14.2000 67.4000 15.8000 ;
	    RECT 69.4000 15.4000 69.8000 16.2000 ;
	    RECT 70.2000 15.6000 70.6000 19.9000 ;
	    RECT 72.3000 17.2000 72.7000 19.9000 ;
	    RECT 74.5000 19.2000 74.9000 19.9000 ;
	    RECT 74.5000 18.8000 75.4000 19.2000 ;
	    RECT 72.3000 16.8000 73.0000 17.2000 ;
	    RECT 73.8000 16.8000 74.2000 17.2000 ;
	    RECT 72.3000 16.2000 72.7000 16.8000 ;
	    RECT 73.8000 16.2000 74.1000 16.8000 ;
	    RECT 74.5000 16.2000 74.9000 18.8000 ;
	    RECT 72.3000 15.9000 73.0000 16.2000 ;
	    RECT 70.2000 15.4000 72.2000 15.6000 ;
	    RECT 70.2000 15.3000 72.3000 15.4000 ;
	    RECT 68.2000 14.8000 69.0000 15.2000 ;
	    RECT 71.9000 15.0000 72.3000 15.3000 ;
	    RECT 72.7000 15.2000 73.0000 15.9000 ;
	    RECT 73.4000 15.9000 74.1000 16.2000 ;
	    RECT 74.4000 15.9000 74.9000 16.2000 ;
	    RECT 73.4000 15.8000 73.8000 15.9000 ;
	    RECT 63.8000 14.1000 64.2000 14.2000 ;
	    RECT 63.0000 13.8000 64.6000 14.1000 ;
	    RECT 65.3000 13.8000 66.6000 14.2000 ;
	    RECT 67.1000 14.1000 67.9000 14.2000 ;
	    RECT 67.1000 13.9000 68.0000 14.1000 ;
	    RECT 63.0000 11.1000 63.4000 13.8000 ;
	    RECT 64.2000 13.6000 64.6000 13.8000 ;
	    RECT 63.9000 13.1000 65.7000 13.3000 ;
	    RECT 66.2000 13.1000 66.5000 13.8000 ;
	    RECT 63.8000 13.0000 65.8000 13.1000 ;
	    RECT 63.8000 11.1000 64.2000 13.0000 ;
	    RECT 65.4000 11.1000 65.8000 13.0000 ;
	    RECT 66.2000 11.1000 66.6000 13.1000 ;
	    RECT 67.6000 11.1000 68.0000 13.9000 ;
	    RECT 72.0000 13.5000 72.3000 15.0000 ;
	    RECT 72.6000 14.8000 73.0000 15.2000 ;
	    RECT 71.1000 13.2000 72.3000 13.5000 ;
	    RECT 70.2000 12.4000 70.6000 13.2000 ;
	    RECT 71.1000 12.1000 71.4000 13.2000 ;
	    RECT 72.7000 13.1000 73.0000 14.8000 ;
	    RECT 74.4000 14.2000 74.7000 15.9000 ;
	    RECT 75.0000 15.1000 75.4000 15.2000 ;
	    RECT 75.8000 15.1000 76.2000 15.2000 ;
	    RECT 75.0000 14.8000 76.2000 15.1000 ;
	    RECT 75.0000 14.4000 75.4000 14.8000 ;
	    RECT 73.4000 13.8000 74.7000 14.2000 ;
	    RECT 75.8000 14.1000 76.2000 14.2000 ;
	    RECT 76.6000 14.1000 77.0000 19.9000 ;
	    RECT 78.2000 15.6000 78.6000 19.9000 ;
	    RECT 80.3000 16.2000 80.7000 19.9000 ;
	    RECT 82.2000 17.9000 82.6000 19.9000 ;
	    RECT 82.3000 17.8000 82.6000 17.9000 ;
	    RECT 83.8000 17.9000 84.2000 19.9000 ;
	    RECT 85.4000 17.9000 85.8000 19.9000 ;
	    RECT 83.8000 17.8000 84.1000 17.9000 ;
	    RECT 82.3000 17.5000 84.1000 17.8000 ;
	    RECT 85.5000 17.8000 85.8000 17.9000 ;
	    RECT 87.0000 17.9000 87.4000 19.9000 ;
	    RECT 87.0000 17.8000 87.3000 17.9000 ;
	    RECT 85.5000 17.5000 87.3000 17.8000 ;
	    RECT 83.0000 16.4000 83.4000 17.2000 ;
	    RECT 83.8000 16.2000 84.1000 17.5000 ;
	    RECT 86.2000 16.4000 86.6000 17.2000 ;
	    RECT 87.0000 16.2000 87.3000 17.5000 ;
	    RECT 88.1000 16.2000 88.5000 19.9000 ;
	    RECT 80.3000 15.9000 81.0000 16.2000 ;
	    RECT 80.6000 15.8000 81.0000 15.9000 ;
	    RECT 78.2000 15.4000 80.2000 15.6000 ;
	    RECT 78.2000 15.3000 80.3000 15.4000 ;
	    RECT 79.9000 15.0000 80.3000 15.3000 ;
	    RECT 80.7000 15.2000 81.0000 15.8000 ;
	    RECT 81.4000 15.4000 81.8000 16.2000 ;
	    RECT 83.8000 15.8000 84.2000 16.2000 ;
	    RECT 87.0000 15.8000 87.4000 16.2000 ;
	    RECT 87.8000 15.9000 88.5000 16.2000 ;
	    RECT 87.8000 15.8000 88.2000 15.9000 ;
	    RECT 75.4000 13.8000 77.0000 14.1000 ;
	    RECT 73.5000 13.1000 73.8000 13.8000 ;
	    RECT 75.4000 13.6000 75.8000 13.8000 ;
	    RECT 74.3000 13.1000 76.1000 13.3000 ;
	    RECT 71.0000 11.1000 71.4000 12.1000 ;
	    RECT 72.6000 11.1000 73.0000 13.1000 ;
	    RECT 73.4000 11.1000 73.8000 13.1000 ;
	    RECT 74.2000 13.0000 76.2000 13.1000 ;
	    RECT 74.2000 11.1000 74.6000 13.0000 ;
	    RECT 75.8000 11.1000 76.2000 13.0000 ;
	    RECT 76.6000 11.1000 77.0000 13.8000 ;
	    RECT 80.0000 13.5000 80.3000 15.0000 ;
	    RECT 80.6000 14.8000 81.0000 15.2000 ;
	    RECT 82.2000 14.8000 83.0000 15.2000 ;
	    RECT 79.1000 13.2000 80.3000 13.5000 ;
	    RECT 78.2000 12.4000 78.6000 13.2000 ;
	    RECT 79.1000 12.1000 79.4000 13.2000 ;
	    RECT 80.7000 13.1000 81.0000 14.8000 ;
	    RECT 83.8000 14.2000 84.1000 15.8000 ;
	    RECT 85.4000 14.8000 86.2000 15.2000 ;
	    RECT 87.0000 14.2000 87.3000 15.8000 ;
	    RECT 83.3000 14.1000 84.1000 14.2000 ;
	    RECT 86.5000 14.1000 87.3000 14.2000 ;
	    RECT 79.0000 11.1000 79.4000 12.1000 ;
	    RECT 80.6000 11.1000 81.0000 13.1000 ;
	    RECT 83.2000 13.9000 84.1000 14.1000 ;
	    RECT 86.4000 13.9000 87.3000 14.1000 ;
	    RECT 87.8000 15.2000 88.1000 15.8000 ;
	    RECT 90.2000 15.6000 90.6000 19.9000 ;
	    RECT 91.8000 17.9000 92.2000 19.9000 ;
	    RECT 91.9000 17.8000 92.2000 17.9000 ;
	    RECT 93.4000 17.9000 93.8000 19.9000 ;
	    RECT 93.4000 17.8000 93.7000 17.9000 ;
	    RECT 91.9000 17.5000 93.7000 17.8000 ;
	    RECT 92.6000 16.4000 93.0000 17.2000 ;
	    RECT 93.4000 16.2000 93.7000 17.5000 ;
	    RECT 94.5000 16.2000 94.9000 19.9000 ;
	    RECT 88.6000 15.4000 90.6000 15.6000 ;
	    RECT 91.0000 15.4000 91.4000 16.2000 ;
	    RECT 93.4000 15.8000 93.8000 16.2000 ;
	    RECT 94.2000 15.9000 94.9000 16.2000 ;
	    RECT 88.5000 15.3000 90.6000 15.4000 ;
	    RECT 87.8000 14.8000 88.2000 15.2000 ;
	    RECT 88.5000 15.0000 88.9000 15.3000 ;
	    RECT 83.2000 11.1000 83.6000 13.9000 ;
	    RECT 86.4000 11.1000 86.8000 13.9000 ;
	    RECT 87.8000 13.1000 88.1000 14.8000 ;
	    RECT 88.5000 13.5000 88.8000 15.0000 ;
	    RECT 91.8000 14.8000 92.6000 15.2000 ;
	    RECT 93.4000 14.2000 93.7000 15.8000 ;
	    RECT 92.9000 14.1000 93.7000 14.2000 ;
	    RECT 92.8000 13.9000 93.7000 14.1000 ;
	    RECT 94.2000 15.2000 94.5000 15.9000 ;
	    RECT 96.6000 15.6000 97.0000 19.9000 ;
	    RECT 98.2000 17.1000 98.6000 19.9000 ;
	    RECT 97.4000 16.8000 98.6000 17.1000 ;
	    RECT 97.4000 16.2000 97.7000 16.8000 ;
	    RECT 97.4000 15.8000 97.8000 16.2000 ;
	    RECT 95.0000 15.4000 97.0000 15.6000 ;
	    RECT 94.9000 15.3000 97.0000 15.4000 ;
	    RECT 94.2000 14.8000 94.6000 15.2000 ;
	    RECT 94.9000 15.0000 95.3000 15.3000 ;
	    RECT 88.5000 13.2000 89.7000 13.5000 ;
	    RECT 87.8000 11.1000 88.2000 13.1000 ;
	    RECT 89.4000 12.1000 89.7000 13.2000 ;
	    RECT 90.2000 12.4000 90.6000 13.2000 ;
	    RECT 89.4000 11.1000 89.8000 12.1000 ;
	    RECT 92.8000 11.1000 93.2000 13.9000 ;
	    RECT 94.2000 13.1000 94.5000 14.8000 ;
	    RECT 94.9000 13.5000 95.2000 15.0000 ;
	    RECT 97.4000 14.1000 97.8000 14.2000 ;
	    RECT 96.6000 13.8000 97.8000 14.1000 ;
	    RECT 94.9000 13.2000 96.1000 13.5000 ;
	    RECT 94.2000 11.1000 94.6000 13.1000 ;
	    RECT 95.8000 12.1000 96.1000 13.2000 ;
	    RECT 96.6000 13.2000 96.9000 13.8000 ;
	    RECT 97.4000 13.4000 97.8000 13.8000 ;
	    RECT 96.6000 12.4000 97.0000 13.2000 ;
	    RECT 98.2000 13.1000 98.6000 16.8000 ;
	    RECT 99.0000 16.1000 99.4000 16.6000 ;
	    RECT 99.8000 16.1000 100.2000 19.9000 ;
	    RECT 101.4000 17.9000 101.8000 19.9000 ;
	    RECT 101.5000 17.8000 101.8000 17.9000 ;
	    RECT 103.0000 17.9000 103.4000 19.9000 ;
	    RECT 103.0000 17.8000 103.3000 17.9000 ;
	    RECT 101.5000 17.5000 103.3000 17.8000 ;
	    RECT 101.5000 16.2000 101.8000 17.5000 ;
	    RECT 102.2000 16.4000 102.6000 17.2000 ;
	    RECT 99.0000 15.8000 100.2000 16.1000 ;
	    RECT 101.4000 15.8000 101.8000 16.2000 ;
	    RECT 98.2000 12.8000 99.1000 13.1000 ;
	    RECT 95.8000 11.1000 96.2000 12.1000 ;
	    RECT 98.7000 11.1000 99.1000 12.8000 ;
	    RECT 99.8000 11.1000 100.2000 15.8000 ;
	    RECT 101.5000 14.2000 101.8000 15.8000 ;
	    RECT 104.6000 15.6000 105.0000 19.9000 ;
	    RECT 106.7000 16.2000 107.1000 19.9000 ;
	    RECT 107.8000 17.9000 108.2000 19.9000 ;
	    RECT 107.9000 17.8000 108.2000 17.9000 ;
	    RECT 109.4000 17.9000 109.8000 19.9000 ;
	    RECT 111.8000 19.1000 112.2000 19.2000 ;
	    RECT 112.6000 19.1000 113.0000 19.9000 ;
	    RECT 111.8000 18.8000 113.0000 19.1000 ;
	    RECT 112.6000 17.9000 113.0000 18.8000 ;
	    RECT 109.4000 17.8000 109.7000 17.9000 ;
	    RECT 107.9000 17.5000 109.7000 17.8000 ;
	    RECT 112.7000 17.8000 113.0000 17.9000 ;
	    RECT 114.2000 17.9000 114.6000 19.9000 ;
	    RECT 114.2000 17.8000 114.5000 17.9000 ;
	    RECT 112.7000 17.5000 114.5000 17.8000 ;
	    RECT 107.9000 16.2000 108.2000 17.5000 ;
	    RECT 108.6000 16.4000 109.0000 17.2000 ;
	    RECT 112.7000 16.2000 113.0000 17.5000 ;
	    RECT 113.4000 16.4000 113.8000 17.2000 ;
	    RECT 116.1000 16.2000 116.5000 19.9000 ;
	    RECT 106.7000 15.9000 107.4000 16.2000 ;
	    RECT 104.6000 15.4000 106.6000 15.6000 ;
	    RECT 104.6000 15.3000 106.7000 15.4000 ;
	    RECT 102.6000 14.8000 103.4000 15.2000 ;
	    RECT 106.3000 15.0000 106.7000 15.3000 ;
	    RECT 107.1000 15.2000 107.4000 15.9000 ;
	    RECT 107.8000 15.8000 108.2000 16.2000 ;
	    RECT 101.5000 14.1000 102.3000 14.2000 ;
	    RECT 101.5000 13.9000 102.4000 14.1000 ;
	    RECT 102.0000 11.1000 102.4000 13.9000 ;
	    RECT 106.4000 13.5000 106.7000 15.0000 ;
	    RECT 107.0000 14.8000 107.4000 15.2000 ;
	    RECT 105.5000 13.2000 106.7000 13.5000 ;
	    RECT 104.6000 12.4000 105.0000 13.2000 ;
	    RECT 105.5000 12.1000 105.8000 13.2000 ;
	    RECT 107.1000 13.1000 107.4000 14.8000 ;
	    RECT 107.9000 14.2000 108.2000 15.8000 ;
	    RECT 110.2000 16.1000 110.6000 16.2000 ;
	    RECT 111.0000 16.1000 111.4000 16.2000 ;
	    RECT 110.2000 15.8000 111.4000 16.1000 ;
	    RECT 112.6000 15.8000 113.0000 16.2000 ;
	    RECT 110.2000 15.4000 110.6000 15.8000 ;
	    RECT 109.0000 14.8000 109.8000 15.2000 ;
	    RECT 112.7000 14.2000 113.0000 15.8000 ;
	    RECT 115.8000 15.9000 116.5000 16.2000 ;
	    RECT 115.8000 15.2000 116.1000 15.9000 ;
	    RECT 118.2000 15.6000 118.6000 19.9000 ;
	    RECT 119.3000 16.2000 119.7000 19.9000 ;
	    RECT 116.6000 15.4000 118.6000 15.6000 ;
	    RECT 116.5000 15.3000 118.6000 15.4000 ;
	    RECT 119.0000 15.9000 119.7000 16.2000 ;
	    RECT 119.0000 15.8000 119.4000 15.9000 ;
	    RECT 113.8000 14.8000 114.6000 15.2000 ;
	    RECT 115.8000 14.8000 116.2000 15.2000 ;
	    RECT 116.5000 15.0000 116.9000 15.3000 ;
	    RECT 119.0000 15.2000 119.3000 15.8000 ;
	    RECT 121.4000 15.6000 121.8000 19.9000 ;
	    RECT 122.2000 17.9000 122.6000 19.9000 ;
	    RECT 122.3000 17.8000 122.6000 17.9000 ;
	    RECT 123.8000 17.9000 124.2000 19.9000 ;
	    RECT 125.4000 17.9000 125.8000 19.9000 ;
	    RECT 123.8000 17.8000 124.1000 17.9000 ;
	    RECT 122.3000 17.5000 124.1000 17.8000 ;
	    RECT 125.5000 17.8000 125.8000 17.9000 ;
	    RECT 127.0000 17.9000 127.4000 19.9000 ;
	    RECT 127.0000 17.8000 127.3000 17.9000 ;
	    RECT 125.5000 17.5000 127.3000 17.8000 ;
	    RECT 122.3000 16.2000 122.6000 17.5000 ;
	    RECT 123.0000 16.4000 123.4000 17.2000 ;
	    RECT 125.5000 16.2000 125.8000 17.5000 ;
	    RECT 126.2000 16.4000 126.6000 17.2000 ;
	    RECT 128.6000 16.2000 129.0000 19.9000 ;
	    RECT 122.2000 15.8000 122.6000 16.2000 ;
	    RECT 119.8000 15.4000 121.8000 15.6000 ;
	    RECT 119.7000 15.3000 121.8000 15.4000 ;
	    RECT 107.9000 14.1000 108.7000 14.2000 ;
	    RECT 112.7000 14.1000 113.5000 14.2000 ;
	    RECT 107.9000 13.9000 108.8000 14.1000 ;
	    RECT 112.7000 13.9000 113.6000 14.1000 ;
	    RECT 105.4000 11.1000 105.8000 12.1000 ;
	    RECT 107.0000 11.1000 107.4000 13.1000 ;
	    RECT 108.4000 11.1000 108.8000 13.9000 ;
	    RECT 113.2000 11.1000 113.6000 13.9000 ;
	    RECT 115.8000 13.1000 116.1000 14.8000 ;
	    RECT 116.5000 13.5000 116.8000 15.0000 ;
	    RECT 119.0000 14.8000 119.4000 15.2000 ;
	    RECT 119.7000 15.0000 120.1000 15.3000 ;
	    RECT 116.5000 13.2000 117.7000 13.5000 ;
	    RECT 115.8000 11.1000 116.2000 13.1000 ;
	    RECT 117.4000 12.1000 117.7000 13.2000 ;
	    RECT 118.2000 12.4000 118.6000 13.2000 ;
	    RECT 119.0000 13.1000 119.3000 14.8000 ;
	    RECT 119.7000 13.5000 120.0000 15.0000 ;
	    RECT 122.3000 14.2000 122.6000 15.8000 ;
	    RECT 124.6000 15.4000 125.0000 16.2000 ;
	    RECT 125.4000 15.8000 125.8000 16.2000 ;
	    RECT 123.4000 14.8000 124.2000 15.2000 ;
	    RECT 125.5000 14.2000 125.8000 15.8000 ;
	    RECT 127.8000 15.4000 128.2000 16.2000 ;
	    RECT 128.6000 15.9000 129.7000 16.2000 ;
	    RECT 130.2000 15.9000 130.6000 19.9000 ;
	    RECT 131.3000 18.2000 131.7000 19.9000 ;
	    RECT 131.0000 17.8000 131.7000 18.2000 ;
	    RECT 131.3000 16.2000 131.7000 17.8000 ;
	    RECT 129.4000 15.6000 129.7000 15.9000 ;
	    RECT 129.4000 15.2000 130.0000 15.6000 ;
	    RECT 126.6000 14.8000 127.4000 15.2000 ;
	    RECT 122.3000 14.1000 123.1000 14.2000 ;
	    RECT 125.5000 14.1000 126.3000 14.2000 ;
	    RECT 122.3000 13.9000 123.2000 14.1000 ;
	    RECT 125.5000 13.9000 126.4000 14.1000 ;
	    RECT 119.7000 13.2000 120.9000 13.5000 ;
	    RECT 117.4000 11.1000 117.8000 12.1000 ;
	    RECT 119.0000 11.1000 119.4000 13.1000 ;
	    RECT 120.6000 12.1000 120.9000 13.2000 ;
	    RECT 121.4000 12.4000 121.8000 13.2000 ;
	    RECT 120.6000 11.1000 121.0000 12.1000 ;
	    RECT 122.8000 11.1000 123.2000 13.9000 ;
	    RECT 126.0000 11.1000 126.4000 13.9000 ;
	    RECT 129.4000 13.7000 129.7000 15.2000 ;
	    RECT 130.3000 14.8000 130.6000 15.9000 ;
	    RECT 128.6000 13.4000 129.7000 13.7000 ;
	    RECT 128.6000 11.1000 129.0000 13.4000 ;
	    RECT 130.2000 11.1000 130.6000 14.8000 ;
	    RECT 131.0000 15.9000 131.7000 16.2000 ;
	    RECT 131.0000 15.2000 131.3000 15.9000 ;
	    RECT 133.4000 15.6000 133.8000 19.9000 ;
	    RECT 134.5000 16.2000 134.9000 19.9000 ;
	    RECT 131.8000 15.4000 133.8000 15.6000 ;
	    RECT 131.7000 15.3000 133.8000 15.4000 ;
	    RECT 134.2000 15.9000 134.9000 16.2000 ;
	    RECT 131.0000 14.8000 131.4000 15.2000 ;
	    RECT 131.7000 15.0000 132.1000 15.3000 ;
	    RECT 134.2000 15.2000 134.5000 15.9000 ;
	    RECT 136.6000 15.6000 137.0000 19.9000 ;
	    RECT 135.0000 15.4000 137.0000 15.6000 ;
	    RECT 134.9000 15.3000 137.0000 15.4000 ;
	    RECT 131.0000 13.1000 131.3000 14.8000 ;
	    RECT 131.7000 13.5000 132.0000 15.0000 ;
	    RECT 134.2000 14.8000 134.6000 15.2000 ;
	    RECT 134.9000 15.0000 135.3000 15.3000 ;
	    RECT 131.7000 13.2000 132.9000 13.5000 ;
	    RECT 131.0000 11.1000 131.4000 13.1000 ;
	    RECT 132.6000 12.1000 132.9000 13.2000 ;
	    RECT 133.4000 12.4000 133.8000 13.2000 ;
	    RECT 134.2000 13.1000 134.5000 14.8000 ;
	    RECT 134.9000 13.5000 135.2000 15.0000 ;
	    RECT 137.4000 14.1000 137.8000 14.2000 ;
	    RECT 138.2000 14.1000 138.6000 19.9000 ;
	    RECT 140.1000 19.2000 140.5000 19.9000 ;
	    RECT 140.1000 18.8000 141.0000 19.2000 ;
	    RECT 139.4000 16.8000 139.8000 17.2000 ;
	    RECT 139.4000 16.2000 139.7000 16.8000 ;
	    RECT 140.1000 16.2000 140.5000 18.8000 ;
	    RECT 143.3000 17.2000 143.7000 19.9000 ;
	    RECT 142.6000 16.8000 143.0000 17.2000 ;
	    RECT 143.3000 16.8000 144.2000 17.2000 ;
	    RECT 142.6000 16.2000 142.9000 16.8000 ;
	    RECT 143.3000 16.2000 143.7000 16.8000 ;
	    RECT 139.0000 15.9000 139.7000 16.2000 ;
	    RECT 140.0000 15.9000 140.5000 16.2000 ;
	    RECT 142.2000 15.9000 142.9000 16.2000 ;
	    RECT 143.2000 15.9000 143.7000 16.2000 ;
	    RECT 139.0000 15.8000 139.4000 15.9000 ;
	    RECT 140.0000 14.2000 140.3000 15.9000 ;
	    RECT 142.2000 15.8000 142.6000 15.9000 ;
	    RECT 140.6000 15.1000 141.0000 15.2000 ;
	    RECT 142.2000 15.1000 142.6000 15.2000 ;
	    RECT 140.6000 14.8000 142.6000 15.1000 ;
	    RECT 140.6000 14.4000 141.0000 14.8000 ;
	    RECT 143.2000 14.2000 143.5000 15.9000 ;
	    RECT 143.8000 14.4000 144.2000 15.2000 ;
	    RECT 137.4000 13.8000 138.6000 14.1000 ;
	    RECT 139.0000 13.8000 140.3000 14.2000 ;
	    RECT 141.4000 14.1000 141.8000 14.2000 ;
	    RECT 141.0000 13.8000 141.8000 14.1000 ;
	    RECT 142.2000 13.8000 143.5000 14.2000 ;
	    RECT 144.6000 14.1000 145.0000 14.2000 ;
	    RECT 145.4000 14.1000 145.8000 19.9000 ;
	    RECT 147.0000 17.9000 147.4000 19.9000 ;
	    RECT 147.1000 17.8000 147.4000 17.9000 ;
	    RECT 148.6000 17.9000 149.0000 19.9000 ;
	    RECT 148.6000 17.8000 148.9000 17.9000 ;
	    RECT 147.1000 17.5000 148.9000 17.8000 ;
	    RECT 147.1000 16.2000 147.4000 17.5000 ;
	    RECT 147.8000 16.4000 148.2000 17.2000 ;
	    RECT 150.5000 16.2000 150.9000 19.9000 ;
	    RECT 147.0000 15.8000 147.4000 16.2000 ;
	    RECT 144.2000 13.8000 145.8000 14.1000 ;
	    RECT 147.1000 14.2000 147.4000 15.8000 ;
	    RECT 149.4000 15.4000 149.8000 16.2000 ;
	    RECT 150.2000 15.9000 150.9000 16.2000 ;
	    RECT 150.2000 15.2000 150.5000 15.9000 ;
	    RECT 152.6000 15.6000 153.0000 19.9000 ;
	    RECT 153.8000 16.8000 154.2000 17.2000 ;
	    RECT 153.8000 16.2000 154.1000 16.8000 ;
	    RECT 154.5000 16.2000 154.9000 19.9000 ;
	    RECT 153.4000 15.9000 154.1000 16.2000 ;
	    RECT 154.4000 15.9000 154.9000 16.2000 ;
	    RECT 153.4000 15.8000 153.8000 15.9000 ;
	    RECT 151.0000 15.4000 153.0000 15.6000 ;
	    RECT 150.9000 15.3000 153.0000 15.4000 ;
	    RECT 148.2000 14.8000 149.0000 15.2000 ;
	    RECT 150.2000 14.8000 150.6000 15.2000 ;
	    RECT 150.9000 15.0000 151.3000 15.3000 ;
	    RECT 153.4000 15.1000 153.8000 15.2000 ;
	    RECT 154.4000 15.1000 154.7000 15.9000 ;
	    RECT 147.1000 14.1000 147.9000 14.2000 ;
	    RECT 147.1000 13.9000 148.0000 14.1000 ;
	    RECT 134.9000 13.2000 136.1000 13.5000 ;
	    RECT 132.6000 11.1000 133.0000 12.1000 ;
	    RECT 134.2000 11.1000 134.6000 13.1000 ;
	    RECT 135.8000 12.1000 136.1000 13.2000 ;
	    RECT 136.6000 12.4000 137.0000 13.2000 ;
	    RECT 135.8000 11.1000 136.2000 12.1000 ;
	    RECT 138.2000 11.1000 138.6000 13.8000 ;
	    RECT 139.1000 13.1000 139.4000 13.8000 ;
	    RECT 141.0000 13.6000 141.4000 13.8000 ;
	    RECT 139.9000 13.1000 141.7000 13.3000 ;
	    RECT 142.3000 13.1000 142.6000 13.8000 ;
	    RECT 144.2000 13.6000 144.6000 13.8000 ;
	    RECT 143.1000 13.1000 144.9000 13.3000 ;
	    RECT 139.0000 11.1000 139.4000 13.1000 ;
	    RECT 139.8000 13.0000 141.8000 13.1000 ;
	    RECT 139.8000 11.1000 140.2000 13.0000 ;
	    RECT 141.4000 11.1000 141.8000 13.0000 ;
	    RECT 142.2000 11.1000 142.6000 13.1000 ;
	    RECT 143.0000 13.0000 145.0000 13.1000 ;
	    RECT 143.0000 11.1000 143.4000 13.0000 ;
	    RECT 144.6000 11.1000 145.0000 13.0000 ;
	    RECT 145.4000 11.1000 145.8000 13.8000 ;
	    RECT 147.6000 11.1000 148.0000 13.9000 ;
	    RECT 150.2000 13.1000 150.5000 14.8000 ;
	    RECT 150.9000 13.5000 151.2000 15.0000 ;
	    RECT 153.4000 14.8000 154.7000 15.1000 ;
	    RECT 154.4000 14.2000 154.7000 14.8000 ;
	    RECT 155.0000 14.4000 155.4000 15.2000 ;
	    RECT 153.4000 13.8000 154.7000 14.2000 ;
	    RECT 155.8000 14.1000 156.2000 14.2000 ;
	    RECT 157.4000 14.1000 157.8000 19.9000 ;
	    RECT 159.0000 17.9000 159.4000 19.9000 ;
	    RECT 159.1000 17.8000 159.4000 17.9000 ;
	    RECT 160.6000 17.9000 161.0000 19.9000 ;
	    RECT 162.2000 17.9000 162.6000 19.9000 ;
	    RECT 160.6000 17.8000 160.9000 17.9000 ;
	    RECT 159.1000 17.5000 160.9000 17.8000 ;
	    RECT 162.3000 17.8000 162.6000 17.9000 ;
	    RECT 163.8000 17.9000 164.2000 19.9000 ;
	    RECT 163.8000 17.8000 164.1000 17.9000 ;
	    RECT 162.3000 17.5000 164.1000 17.8000 ;
	    RECT 159.8000 16.4000 160.2000 17.2000 ;
	    RECT 160.6000 16.2000 160.9000 17.5000 ;
	    RECT 163.0000 16.4000 163.4000 17.2000 ;
	    RECT 163.8000 16.2000 164.1000 17.5000 ;
	    RECT 165.0000 16.8000 165.4000 17.2000 ;
	    RECT 165.0000 16.2000 165.3000 16.8000 ;
	    RECT 165.7000 16.2000 166.1000 19.9000 ;
	    RECT 160.6000 15.8000 161.0000 16.2000 ;
	    RECT 159.0000 14.8000 159.8000 15.2000 ;
	    RECT 160.6000 14.2000 160.9000 15.8000 ;
	    RECT 161.4000 15.4000 161.8000 16.2000 ;
	    RECT 163.8000 15.8000 164.2000 16.2000 ;
	    RECT 164.6000 15.9000 165.3000 16.2000 ;
	    RECT 165.6000 15.9000 166.1000 16.2000 ;
	    RECT 164.6000 15.8000 165.0000 15.9000 ;
	    RECT 162.2000 14.8000 163.0000 15.2000 ;
	    RECT 163.8000 14.2000 164.1000 15.8000 ;
	    RECT 165.6000 15.2000 165.9000 15.9000 ;
	    RECT 165.4000 14.8000 165.9000 15.2000 ;
	    RECT 165.6000 14.2000 165.9000 14.8000 ;
	    RECT 166.2000 14.4000 166.6000 15.2000 ;
	    RECT 160.1000 14.1000 160.9000 14.2000 ;
	    RECT 163.3000 14.1000 164.1000 14.2000 ;
	    RECT 155.4000 13.8000 157.8000 14.1000 ;
	    RECT 150.9000 13.2000 152.1000 13.5000 ;
	    RECT 150.2000 11.1000 150.6000 13.1000 ;
	    RECT 151.8000 12.1000 152.1000 13.2000 ;
	    RECT 152.6000 12.4000 153.0000 13.2000 ;
	    RECT 153.5000 13.1000 153.8000 13.8000 ;
	    RECT 155.4000 13.6000 155.8000 13.8000 ;
	    RECT 154.3000 13.1000 156.1000 13.3000 ;
	    RECT 151.8000 11.1000 152.2000 12.1000 ;
	    RECT 153.4000 11.1000 153.8000 13.1000 ;
	    RECT 154.2000 13.0000 156.2000 13.1000 ;
	    RECT 154.2000 11.1000 154.6000 13.0000 ;
	    RECT 155.8000 11.1000 156.2000 13.0000 ;
	    RECT 157.4000 11.1000 157.8000 13.8000 ;
	    RECT 160.0000 13.9000 160.9000 14.1000 ;
	    RECT 163.2000 13.9000 164.1000 14.1000 ;
	    RECT 160.0000 11.1000 160.4000 13.9000 ;
	    RECT 163.2000 11.1000 163.6000 13.9000 ;
	    RECT 164.6000 13.8000 165.9000 14.2000 ;
	    RECT 167.0000 14.1000 167.4000 14.2000 ;
	    RECT 167.8000 14.1000 168.2000 19.9000 ;
	    RECT 166.6000 13.8000 168.2000 14.1000 ;
	    RECT 164.7000 13.1000 165.0000 13.8000 ;
	    RECT 166.6000 13.6000 167.0000 13.8000 ;
	    RECT 165.5000 13.1000 167.3000 13.3000 ;
	    RECT 164.6000 11.1000 165.0000 13.1000 ;
	    RECT 165.4000 13.0000 167.4000 13.1000 ;
	    RECT 165.4000 11.1000 165.8000 13.0000 ;
	    RECT 167.0000 11.1000 167.4000 13.0000 ;
	    RECT 167.8000 11.1000 168.2000 13.8000 ;
	    RECT 169.4000 15.9000 169.8000 19.9000 ;
	    RECT 171.0000 16.2000 171.4000 19.9000 ;
	    RECT 170.3000 15.9000 171.4000 16.2000 ;
	    RECT 169.4000 14.8000 169.7000 15.9000 ;
	    RECT 170.3000 15.6000 170.6000 15.9000 ;
	    RECT 170.0000 15.2000 170.6000 15.6000 ;
	    RECT 169.4000 11.1000 169.8000 14.8000 ;
	    RECT 170.3000 13.7000 170.6000 15.2000 ;
	    RECT 170.3000 13.4000 171.4000 13.7000 ;
	    RECT 171.0000 11.1000 171.4000 13.4000 ;
	    RECT 1.9000 9.2000 2.3000 9.9000 ;
	    RECT 1.4000 8.8000 2.3000 9.2000 ;
	    RECT 1.9000 8.2000 2.3000 8.8000 ;
	    RECT 4.3000 8.2000 4.7000 9.9000 ;
	    RECT 6.7000 9.2000 7.1000 9.9000 ;
	    RECT 6.7000 8.8000 7.4000 9.2000 ;
	    RECT 6.7000 8.2000 7.1000 8.8000 ;
	    RECT 1.4000 7.9000 2.3000 8.2000 ;
	    RECT 3.8000 7.9000 4.7000 8.2000 ;
	    RECT 6.2000 7.9000 7.1000 8.2000 ;
	    RECT 7.8000 7.9000 8.2000 9.9000 ;
	    RECT 8.6000 8.0000 9.0000 9.9000 ;
	    RECT 10.2000 8.0000 10.6000 9.9000 ;
	    RECT 8.6000 7.9000 10.6000 8.0000 ;
	    RECT 0.6000 6.8000 1.0000 7.6000 ;
	    RECT 1.4000 1.1000 1.8000 7.9000 ;
	    RECT 3.0000 6.8000 3.4000 7.6000 ;
	    RECT 2.2000 4.4000 2.6000 5.2000 ;
	    RECT 3.0000 5.1000 3.4000 5.2000 ;
	    RECT 3.8000 5.1000 4.2000 7.9000 ;
	    RECT 3.0000 4.8000 4.2000 5.1000 ;
	    RECT 3.8000 1.1000 4.2000 4.8000 ;
	    RECT 6.2000 1.1000 6.6000 7.9000 ;
	    RECT 7.9000 7.2000 8.2000 7.9000 ;
	    RECT 8.7000 7.7000 10.5000 7.9000 ;
	    RECT 9.8000 7.2000 10.2000 7.4000 ;
	    RECT 7.8000 6.8000 9.1000 7.2000 ;
	    RECT 9.8000 7.1000 10.6000 7.2000 ;
	    RECT 11.0000 7.1000 11.4000 9.9000 ;
	    RECT 13.4000 8.9000 13.8000 9.9000 ;
	    RECT 12.6000 7.8000 13.0000 8.6000 ;
	    RECT 13.5000 7.8000 13.8000 8.9000 ;
	    RECT 15.0000 7.9000 15.4000 9.9000 ;
	    RECT 13.5000 7.5000 14.7000 7.8000 ;
	    RECT 9.8000 6.9000 11.4000 7.1000 ;
	    RECT 10.2000 6.8000 11.4000 6.9000 ;
	    RECT 8.8000 6.1000 9.1000 6.8000 ;
	    RECT 7.0000 5.8000 9.1000 6.1000 ;
	    RECT 9.4000 5.8000 9.8000 6.6000 ;
	    RECT 7.0000 5.2000 7.3000 5.8000 ;
	    RECT 7.0000 4.4000 7.4000 5.2000 ;
	    RECT 7.8000 5.1000 8.2000 5.2000 ;
	    RECT 8.8000 5.1000 9.1000 5.8000 ;
	    RECT 7.8000 4.8000 8.5000 5.1000 ;
	    RECT 8.8000 4.8000 9.3000 5.1000 ;
	    RECT 8.2000 4.2000 8.5000 4.8000 ;
	    RECT 8.2000 3.8000 8.6000 4.2000 ;
	    RECT 8.9000 1.1000 9.3000 4.8000 ;
	    RECT 11.0000 1.1000 11.4000 6.8000 ;
	    RECT 14.4000 6.0000 14.7000 7.5000 ;
	    RECT 15.1000 6.2000 15.4000 7.9000 ;
	    RECT 14.3000 5.7000 14.7000 6.0000 ;
	    RECT 15.0000 5.8000 15.4000 6.2000 ;
	    RECT 12.6000 5.6000 14.7000 5.7000 ;
	    RECT 12.6000 5.4000 14.6000 5.6000 ;
	    RECT 12.6000 1.1000 13.0000 5.4000 ;
	    RECT 15.1000 5.1000 15.4000 5.8000 ;
	    RECT 14.7000 4.8000 15.4000 5.1000 ;
	    RECT 15.8000 6.1000 16.2000 9.9000 ;
	    RECT 17.7000 9.2000 18.1000 9.9000 ;
	    RECT 17.4000 8.8000 18.1000 9.2000 ;
	    RECT 17.7000 8.2000 18.1000 8.8000 ;
	    RECT 17.7000 7.9000 18.6000 8.2000 ;
	    RECT 16.6000 6.1000 17.0000 6.2000 ;
	    RECT 15.8000 5.8000 17.0000 6.1000 ;
	    RECT 14.7000 1.1000 15.1000 4.8000 ;
	    RECT 15.8000 1.1000 16.2000 5.8000 ;
	    RECT 17.4000 4.4000 17.8000 5.2000 ;
	    RECT 18.2000 1.1000 18.6000 7.9000 ;
	    RECT 19.8000 7.6000 20.2000 9.9000 ;
	    RECT 19.8000 7.3000 20.9000 7.6000 ;
	    RECT 20.6000 5.8000 20.9000 7.3000 ;
	    RECT 21.4000 7.1000 21.8000 9.9000 ;
	    RECT 23.5000 9.2000 23.9000 9.9000 ;
	    RECT 23.0000 8.8000 23.9000 9.2000 ;
	    RECT 23.5000 8.2000 23.9000 8.8000 ;
	    RECT 23.0000 7.9000 23.9000 8.2000 ;
	    RECT 22.2000 7.1000 22.6000 7.6000 ;
	    RECT 21.4000 6.8000 22.6000 7.1000 ;
	    RECT 21.4000 6.2000 21.8000 6.8000 ;
	    RECT 20.6000 5.4000 21.2000 5.8000 ;
	    RECT 20.6000 5.1000 20.9000 5.4000 ;
	    RECT 21.5000 5.1000 21.8000 6.2000 ;
	    RECT 22.2000 6.2000 22.5000 6.8000 ;
	    RECT 22.2000 5.8000 22.6000 6.2000 ;
	    RECT 19.8000 4.8000 20.9000 5.1000 ;
	    RECT 19.8000 1.1000 20.2000 4.8000 ;
	    RECT 21.4000 1.1000 21.8000 5.1000 ;
	    RECT 23.0000 1.1000 23.4000 7.9000 ;
	    RECT 23.8000 5.1000 24.2000 5.2000 ;
	    RECT 24.6000 5.1000 25.0000 9.9000 ;
	    RECT 27.5000 9.2000 27.9000 9.9000 ;
	    RECT 27.0000 8.8000 27.9000 9.2000 ;
	    RECT 27.5000 8.2000 27.9000 8.8000 ;
	    RECT 29.9000 9.2000 30.3000 9.9000 ;
	    RECT 29.9000 8.8000 30.6000 9.2000 ;
	    RECT 29.9000 8.2000 30.3000 8.8000 ;
	    RECT 27.0000 7.9000 27.9000 8.2000 ;
	    RECT 29.4000 7.9000 30.3000 8.2000 ;
	    RECT 26.2000 6.8000 26.6000 7.6000 ;
	    RECT 23.8000 4.8000 25.0000 5.1000 ;
	    RECT 23.8000 4.4000 24.2000 4.8000 ;
	    RECT 24.6000 1.1000 25.0000 4.8000 ;
	    RECT 27.0000 1.1000 27.4000 7.9000 ;
	    RECT 28.6000 6.8000 29.0000 7.6000 ;
	    RECT 27.8000 4.4000 28.2000 5.2000 ;
	    RECT 29.4000 1.1000 29.8000 7.9000 ;
	    RECT 30.2000 5.1000 30.6000 5.2000 ;
	    RECT 31.0000 5.1000 31.4000 9.9000 ;
	    RECT 33.9000 9.2000 34.3000 9.9000 ;
	    RECT 36.3000 9.2000 36.7000 9.9000 ;
	    RECT 33.9000 8.8000 34.6000 9.2000 ;
	    RECT 35.8000 8.8000 36.7000 9.2000 ;
	    RECT 33.9000 8.2000 34.3000 8.8000 ;
	    RECT 36.3000 8.2000 36.7000 8.8000 ;
	    RECT 38.7000 8.2000 39.1000 9.9000 ;
	    RECT 33.4000 7.9000 34.3000 8.2000 ;
	    RECT 35.8000 7.9000 36.7000 8.2000 ;
	    RECT 38.2000 7.9000 39.1000 8.2000 ;
	    RECT 39.8000 7.9000 40.2000 9.9000 ;
	    RECT 40.6000 8.0000 41.0000 9.9000 ;
	    RECT 42.2000 8.0000 42.6000 9.9000 ;
	    RECT 40.6000 7.9000 42.6000 8.0000 ;
	    RECT 32.6000 6.8000 33.0000 7.6000 ;
	    RECT 30.2000 4.8000 31.4000 5.1000 ;
	    RECT 30.2000 4.4000 30.6000 4.8000 ;
	    RECT 31.0000 1.1000 31.4000 4.8000 ;
	    RECT 33.4000 1.1000 33.8000 7.9000 ;
	    RECT 35.0000 6.8000 35.4000 7.6000 ;
	    RECT 34.2000 4.4000 34.6000 5.2000 ;
	    RECT 35.8000 1.1000 36.2000 7.9000 ;
	    RECT 36.6000 7.1000 37.0000 7.2000 ;
	    RECT 37.4000 7.1000 37.8000 7.6000 ;
	    RECT 36.6000 6.8000 37.8000 7.1000 ;
	    RECT 38.2000 6.1000 38.6000 7.9000 ;
	    RECT 39.9000 7.2000 40.2000 7.9000 ;
	    RECT 40.7000 7.7000 42.5000 7.9000 ;
	    RECT 41.8000 7.2000 42.2000 7.4000 ;
	    RECT 39.8000 6.8000 41.1000 7.2000 ;
	    RECT 41.8000 6.9000 42.6000 7.2000 ;
	    RECT 38.2000 5.8000 40.1000 6.1000 ;
	    RECT 36.6000 5.1000 37.0000 5.2000 ;
	    RECT 37.4000 5.1000 37.8000 5.2000 ;
	    RECT 36.6000 4.8000 37.8000 5.1000 ;
	    RECT 36.6000 4.4000 37.0000 4.8000 ;
	    RECT 38.2000 1.1000 38.6000 5.8000 ;
	    RECT 39.8000 5.2000 40.1000 5.8000 ;
	    RECT 39.8000 5.1000 40.2000 5.2000 ;
	    RECT 40.8000 5.1000 41.1000 6.8000 ;
	    RECT 42.2000 6.8000 42.6000 6.9000 ;
	    RECT 41.4000 5.8000 41.8000 6.6000 ;
	    RECT 42.2000 6.2000 42.5000 6.8000 ;
	    RECT 42.2000 5.8000 42.6000 6.2000 ;
	    RECT 39.8000 4.8000 40.5000 5.1000 ;
	    RECT 40.8000 4.8000 41.3000 5.1000 ;
	    RECT 40.2000 4.2000 40.5000 4.8000 ;
	    RECT 40.9000 4.2000 41.3000 4.8000 ;
	    RECT 40.2000 3.8000 40.6000 4.2000 ;
	    RECT 40.9000 3.8000 41.8000 4.2000 ;
	    RECT 40.9000 1.1000 41.3000 3.8000 ;
	    RECT 43.0000 1.1000 43.4000 9.9000 ;
	    RECT 44.6000 1.1000 45.0000 9.9000 ;
	    RECT 47.5000 9.2000 47.9000 9.9000 ;
	    RECT 47.0000 8.8000 47.9000 9.2000 ;
	    RECT 47.5000 8.2000 47.9000 8.8000 ;
	    RECT 47.0000 7.9000 47.9000 8.2000 ;
	    RECT 46.2000 6.8000 46.6000 7.6000 ;
	    RECT 47.0000 1.1000 47.4000 7.9000 ;
	    RECT 48.6000 7.1000 49.0000 9.9000 ;
	    RECT 47.8000 6.8000 49.0000 7.1000 ;
	    RECT 47.8000 6.2000 48.1000 6.8000 ;
	    RECT 47.8000 5.8000 48.2000 6.2000 ;
	    RECT 48.6000 1.1000 49.0000 6.8000 ;
	    RECT 50.2000 5.1000 50.6000 9.9000 ;
	    RECT 52.1000 9.2000 52.5000 9.9000 ;
	    RECT 51.8000 8.8000 52.5000 9.2000 ;
	    RECT 52.1000 8.2000 52.5000 8.8000 ;
	    RECT 55.5000 9.2000 55.9000 9.9000 ;
	    RECT 56.9000 9.2000 57.3000 9.9000 ;
	    RECT 55.5000 8.8000 56.2000 9.2000 ;
	    RECT 56.9000 8.8000 57.8000 9.2000 ;
	    RECT 55.5000 8.2000 55.9000 8.8000 ;
	    RECT 52.1000 7.9000 53.0000 8.2000 ;
	    RECT 51.8000 5.1000 52.2000 5.2000 ;
	    RECT 50.2000 4.8000 52.2000 5.1000 ;
	    RECT 50.2000 1.1000 50.6000 4.8000 ;
	    RECT 51.8000 4.4000 52.2000 4.8000 ;
	    RECT 52.6000 1.1000 53.0000 7.9000 ;
	    RECT 55.0000 7.9000 55.9000 8.2000 ;
	    RECT 56.9000 8.2000 57.3000 8.8000 ;
	    RECT 56.9000 7.9000 57.8000 8.2000 ;
	    RECT 53.4000 7.1000 53.8000 7.6000 ;
	    RECT 54.2000 7.1000 54.6000 7.6000 ;
	    RECT 53.4000 6.8000 54.6000 7.1000 ;
	    RECT 55.0000 1.1000 55.4000 7.9000 ;
	    RECT 57.4000 1.1000 57.8000 7.9000 ;
	    RECT 59.0000 7.6000 59.4000 9.9000 ;
	    RECT 60.6000 8.1000 61.0000 9.9000 ;
	    RECT 64.3000 9.2000 64.7000 9.9000 ;
	    RECT 64.3000 8.8000 65.0000 9.2000 ;
	    RECT 64.3000 8.2000 64.7000 8.8000 ;
	    RECT 61.4000 8.1000 61.8000 8.2000 ;
	    RECT 60.6000 7.8000 61.8000 8.1000 ;
	    RECT 63.8000 7.9000 64.7000 8.2000 ;
	    RECT 58.2000 6.8000 58.6000 7.6000 ;
	    RECT 59.0000 7.3000 60.1000 7.6000 ;
	    RECT 59.8000 5.8000 60.1000 7.3000 ;
	    RECT 60.6000 7.1000 61.0000 7.8000 ;
	    RECT 63.0000 7.1000 63.4000 7.6000 ;
	    RECT 60.6000 6.8000 63.4000 7.1000 ;
	    RECT 60.6000 6.2000 61.0000 6.8000 ;
	    RECT 59.8000 5.4000 60.4000 5.8000 ;
	    RECT 59.8000 5.1000 60.1000 5.4000 ;
	    RECT 60.7000 5.1000 61.0000 6.2000 ;
	    RECT 59.0000 4.8000 60.1000 5.1000 ;
	    RECT 59.0000 1.1000 59.4000 4.8000 ;
	    RECT 60.6000 1.1000 61.0000 5.1000 ;
	    RECT 63.8000 1.1000 64.2000 7.9000 ;
	    RECT 64.6000 5.1000 65.0000 5.2000 ;
	    RECT 66.2000 5.1000 66.6000 9.9000 ;
	    RECT 64.6000 4.8000 66.6000 5.1000 ;
	    RECT 64.6000 4.4000 65.0000 4.8000 ;
	    RECT 66.2000 1.1000 66.6000 4.8000 ;
	    RECT 67.0000 1.1000 67.4000 9.9000 ;
	    RECT 68.9000 9.2000 69.3000 9.9000 ;
	    RECT 72.3000 9.2000 72.7000 9.9000 ;
	    RECT 68.9000 8.8000 69.8000 9.2000 ;
	    RECT 72.3000 8.8000 73.0000 9.2000 ;
	    RECT 68.9000 8.2000 69.3000 8.8000 ;
	    RECT 72.3000 8.2000 72.7000 8.8000 ;
	    RECT 68.9000 7.9000 69.8000 8.2000 ;
	    RECT 69.4000 1.1000 69.8000 7.9000 ;
	    RECT 71.8000 7.9000 72.7000 8.2000 ;
	    RECT 70.2000 7.1000 70.6000 7.6000 ;
	    RECT 71.0000 7.1000 71.4000 7.6000 ;
	    RECT 70.2000 6.8000 71.4000 7.1000 ;
	    RECT 71.8000 1.1000 72.2000 7.9000 ;
	    RECT 72.6000 5.1000 73.0000 5.2000 ;
	    RECT 73.4000 5.1000 73.8000 9.9000 ;
	    RECT 76.3000 9.2000 76.7000 9.9000 ;
	    RECT 75.8000 8.8000 76.7000 9.2000 ;
	    RECT 76.3000 8.2000 76.7000 8.8000 ;
	    RECT 75.8000 7.9000 76.7000 8.2000 ;
	    RECT 75.0000 6.8000 75.4000 7.6000 ;
	    RECT 72.6000 4.8000 73.8000 5.1000 ;
	    RECT 72.6000 4.4000 73.0000 4.8000 ;
	    RECT 73.4000 1.1000 73.8000 4.8000 ;
	    RECT 75.8000 1.1000 76.2000 7.9000 ;
	    RECT 76.6000 5.1000 77.0000 5.2000 ;
	    RECT 77.4000 5.1000 77.8000 9.9000 ;
	    RECT 79.0000 7.6000 79.4000 9.9000 ;
	    RECT 79.0000 7.3000 80.1000 7.6000 ;
	    RECT 79.8000 5.8000 80.1000 7.3000 ;
	    RECT 80.6000 6.2000 81.0000 9.9000 ;
	    RECT 79.8000 5.4000 80.4000 5.8000 ;
	    RECT 79.8000 5.1000 80.1000 5.4000 ;
	    RECT 80.7000 5.1000 81.0000 6.2000 ;
	    RECT 76.6000 4.8000 77.8000 5.1000 ;
	    RECT 76.6000 4.4000 77.0000 4.8000 ;
	    RECT 77.4000 1.1000 77.8000 4.8000 ;
	    RECT 79.0000 4.8000 80.1000 5.1000 ;
	    RECT 79.0000 1.1000 79.4000 4.8000 ;
	    RECT 80.6000 1.1000 81.0000 5.1000 ;
	    RECT 82.2000 5.1000 82.6000 9.9000 ;
	    RECT 83.3000 9.2000 83.7000 9.9000 ;
	    RECT 83.3000 8.8000 84.2000 9.2000 ;
	    RECT 83.3000 8.2000 83.7000 8.8000 ;
	    RECT 83.3000 7.9000 84.2000 8.2000 ;
	    RECT 83.0000 5.1000 83.4000 5.2000 ;
	    RECT 82.2000 4.8000 83.4000 5.1000 ;
	    RECT 82.2000 1.1000 82.6000 4.8000 ;
	    RECT 83.0000 4.4000 83.4000 4.8000 ;
	    RECT 83.8000 1.1000 84.2000 7.9000 ;
	    RECT 84.6000 6.8000 85.0000 7.6000 ;
	    RECT 86.2000 5.1000 86.6000 9.9000 ;
	    RECT 87.3000 9.2000 87.7000 9.9000 ;
	    RECT 90.7000 9.2000 91.1000 9.9000 ;
	    RECT 87.3000 8.8000 88.2000 9.2000 ;
	    RECT 90.7000 8.8000 91.4000 9.2000 ;
	    RECT 87.3000 8.2000 87.7000 8.8000 ;
	    RECT 90.7000 8.2000 91.1000 8.8000 ;
	    RECT 87.3000 7.9000 88.2000 8.2000 ;
	    RECT 87.0000 5.1000 87.4000 5.2000 ;
	    RECT 86.2000 4.8000 87.4000 5.1000 ;
	    RECT 86.2000 1.1000 86.6000 4.8000 ;
	    RECT 87.0000 4.4000 87.4000 4.8000 ;
	    RECT 87.8000 1.1000 88.2000 7.9000 ;
	    RECT 90.2000 7.9000 91.1000 8.2000 ;
	    RECT 88.6000 7.1000 89.0000 7.6000 ;
	    RECT 89.4000 7.1000 89.8000 7.6000 ;
	    RECT 88.6000 6.8000 89.8000 7.1000 ;
	    RECT 90.2000 1.1000 90.6000 7.9000 ;
	    RECT 91.0000 5.1000 91.4000 5.2000 ;
	    RECT 91.8000 5.1000 92.2000 9.9000 ;
	    RECT 94.7000 8.2000 95.1000 9.9000 ;
	    RECT 94.2000 7.9000 95.1000 8.2000 ;
	    RECT 93.4000 6.8000 93.8000 7.6000 ;
	    RECT 91.0000 4.8000 92.2000 5.1000 ;
	    RECT 91.0000 4.4000 91.4000 4.8000 ;
	    RECT 91.8000 1.1000 92.2000 4.8000 ;
	    RECT 94.2000 6.1000 94.6000 7.9000 ;
	    RECT 95.8000 7.1000 96.2000 7.2000 ;
	    RECT 96.6000 7.1000 97.0000 9.9000 ;
	    RECT 97.4000 7.9000 97.8000 9.9000 ;
	    RECT 98.2000 8.0000 98.6000 9.9000 ;
	    RECT 99.8000 8.0000 100.2000 9.9000 ;
	    RECT 100.9000 9.2000 101.3000 9.9000 ;
	    RECT 104.3000 9.2000 104.7000 9.9000 ;
	    RECT 100.6000 8.8000 101.3000 9.2000 ;
	    RECT 103.8000 8.8000 104.7000 9.2000 ;
	    RECT 98.2000 7.9000 100.2000 8.0000 ;
	    RECT 100.9000 8.2000 101.3000 8.8000 ;
	    RECT 104.3000 8.2000 104.7000 8.8000 ;
	    RECT 100.9000 7.9000 101.8000 8.2000 ;
	    RECT 97.5000 7.2000 97.8000 7.9000 ;
	    RECT 98.3000 7.7000 100.1000 7.9000 ;
	    RECT 99.4000 7.2000 99.8000 7.4000 ;
	    RECT 95.8000 6.8000 97.0000 7.1000 ;
	    RECT 97.4000 6.8000 98.7000 7.2000 ;
	    RECT 99.4000 6.9000 100.2000 7.2000 ;
	    RECT 99.8000 6.8000 100.2000 6.9000 ;
	    RECT 95.8000 6.1000 96.2000 6.2000 ;
	    RECT 94.2000 5.8000 96.2000 6.1000 ;
	    RECT 94.2000 1.1000 94.6000 5.8000 ;
	    RECT 96.6000 1.1000 97.0000 6.8000 ;
	    RECT 97.4000 6.1000 97.8000 6.2000 ;
	    RECT 98.4000 6.1000 98.7000 6.8000 ;
	    RECT 97.4000 5.8000 98.7000 6.1000 ;
	    RECT 99.0000 5.8000 99.4000 6.6000 ;
	    RECT 97.4000 5.1000 97.8000 5.2000 ;
	    RECT 98.4000 5.1000 98.7000 5.8000 ;
	    RECT 97.4000 4.8000 98.1000 5.1000 ;
	    RECT 98.4000 4.8000 98.9000 5.1000 ;
	    RECT 97.8000 4.2000 98.1000 4.8000 ;
	    RECT 97.8000 3.8000 98.2000 4.2000 ;
	    RECT 98.5000 1.1000 98.9000 4.8000 ;
	    RECT 100.6000 4.4000 101.0000 5.2000 ;
	    RECT 101.4000 1.1000 101.8000 7.9000 ;
	    RECT 103.8000 7.9000 104.7000 8.2000 ;
	    RECT 103.0000 6.8000 103.4000 7.6000 ;
	    RECT 103.8000 1.1000 104.2000 7.9000 ;
	    RECT 104.6000 5.1000 105.0000 5.2000 ;
	    RECT 105.4000 5.1000 105.8000 9.9000 ;
	    RECT 104.6000 4.8000 105.8000 5.1000 ;
	    RECT 104.6000 4.4000 105.0000 4.8000 ;
	    RECT 105.4000 1.1000 105.8000 4.8000 ;
	    RECT 107.8000 5.1000 108.2000 9.9000 ;
	    RECT 108.9000 9.2000 109.3000 9.9000 ;
	    RECT 108.9000 8.8000 109.8000 9.2000 ;
	    RECT 108.9000 8.2000 109.3000 8.8000 ;
	    RECT 113.9000 8.2000 114.3000 9.9000 ;
	    RECT 108.9000 7.9000 109.8000 8.2000 ;
	    RECT 108.6000 5.1000 109.0000 5.2000 ;
	    RECT 107.8000 4.8000 109.0000 5.1000 ;
	    RECT 107.8000 1.1000 108.2000 4.8000 ;
	    RECT 108.6000 4.4000 109.0000 4.8000 ;
	    RECT 109.4000 1.1000 109.8000 7.9000 ;
	    RECT 113.4000 7.9000 114.3000 8.2000 ;
	    RECT 115.0000 7.9000 115.4000 9.9000 ;
	    RECT 115.8000 8.0000 116.2000 9.9000 ;
	    RECT 117.4000 8.0000 117.8000 9.9000 ;
	    RECT 115.8000 7.9000 117.8000 8.0000 ;
	    RECT 110.2000 6.8000 110.6000 7.6000 ;
	    RECT 112.6000 6.8000 113.0000 7.6000 ;
	    RECT 113.4000 6.1000 113.8000 7.9000 ;
	    RECT 115.1000 7.2000 115.4000 7.9000 ;
	    RECT 115.9000 7.7000 117.7000 7.9000 ;
	    RECT 117.0000 7.2000 117.4000 7.4000 ;
	    RECT 115.0000 6.8000 116.3000 7.2000 ;
	    RECT 117.0000 7.1000 117.8000 7.2000 ;
	    RECT 118.2000 7.1000 118.6000 9.9000 ;
	    RECT 117.0000 6.9000 118.6000 7.1000 ;
	    RECT 117.4000 6.8000 118.6000 6.9000 ;
	    RECT 113.4000 5.8000 115.3000 6.1000 ;
	    RECT 113.4000 1.1000 113.8000 5.8000 ;
	    RECT 115.0000 5.2000 115.3000 5.8000 ;
	    RECT 115.0000 5.1000 115.4000 5.2000 ;
	    RECT 116.0000 5.1000 116.3000 6.8000 ;
	    RECT 116.6000 5.8000 117.0000 6.6000 ;
	    RECT 115.0000 4.8000 115.7000 5.1000 ;
	    RECT 116.0000 4.8000 116.5000 5.1000 ;
	    RECT 115.4000 4.2000 115.7000 4.8000 ;
	    RECT 115.4000 3.8000 115.8000 4.2000 ;
	    RECT 116.1000 1.1000 116.5000 4.8000 ;
	    RECT 118.2000 1.1000 118.6000 6.8000 ;
	    RECT 119.8000 6.2000 120.2000 9.9000 ;
	    RECT 121.4000 7.6000 121.8000 9.9000 ;
	    RECT 123.5000 9.2000 123.9000 9.9000 ;
	    RECT 125.9000 9.2000 126.3000 9.9000 ;
	    RECT 123.5000 8.8000 124.2000 9.2000 ;
	    RECT 125.9000 8.8000 126.6000 9.2000 ;
	    RECT 123.5000 8.2000 123.9000 8.8000 ;
	    RECT 125.9000 8.2000 126.3000 8.8000 ;
	    RECT 123.0000 7.9000 123.9000 8.2000 ;
	    RECT 125.4000 7.9000 126.3000 8.2000 ;
	    RECT 120.7000 7.3000 121.8000 7.6000 ;
	    RECT 119.8000 5.1000 120.1000 6.2000 ;
	    RECT 120.7000 5.8000 121.0000 7.3000 ;
	    RECT 122.2000 6.8000 122.6000 7.6000 ;
	    RECT 120.4000 5.4000 121.0000 5.8000 ;
	    RECT 120.7000 5.1000 121.0000 5.4000 ;
	    RECT 119.8000 1.1000 120.2000 5.1000 ;
	    RECT 120.7000 4.8000 121.8000 5.1000 ;
	    RECT 121.4000 1.1000 121.8000 4.8000 ;
	    RECT 123.0000 1.1000 123.4000 7.9000 ;
	    RECT 124.6000 6.8000 125.0000 7.6000 ;
	    RECT 125.4000 1.1000 125.8000 7.9000 ;
	    RECT 126.2000 5.1000 126.6000 5.2000 ;
	    RECT 127.0000 5.1000 127.4000 9.9000 ;
	    RECT 128.6000 6.1000 129.0000 6.2000 ;
	    RECT 129.4000 6.1000 129.8000 9.9000 ;
	    RECT 128.6000 5.8000 129.8000 6.1000 ;
	    RECT 126.2000 4.8000 127.4000 5.1000 ;
	    RECT 126.2000 4.4000 126.6000 4.8000 ;
	    RECT 127.0000 1.1000 127.4000 4.8000 ;
	    RECT 129.4000 1.1000 129.8000 5.8000 ;
	    RECT 131.0000 5.1000 131.4000 9.9000 ;
	    RECT 132.1000 9.2000 132.5000 9.9000 ;
	    RECT 131.8000 8.8000 132.5000 9.2000 ;
	    RECT 132.1000 8.2000 132.5000 8.8000 ;
	    RECT 132.1000 7.9000 133.0000 8.2000 ;
	    RECT 131.8000 5.1000 132.2000 5.2000 ;
	    RECT 131.0000 4.8000 132.2000 5.1000 ;
	    RECT 131.0000 1.1000 131.4000 4.8000 ;
	    RECT 131.8000 4.4000 132.2000 4.8000 ;
	    RECT 132.6000 1.1000 133.0000 7.9000 ;
	    RECT 133.4000 6.8000 133.8000 7.6000 ;
	    RECT 135.0000 7.1000 135.4000 9.9000 ;
	    RECT 136.1000 9.2000 136.5000 9.9000 ;
	    RECT 138.5000 9.2000 138.9000 9.9000 ;
	    RECT 140.9000 9.2000 141.3000 9.9000 ;
	    RECT 136.1000 8.8000 137.0000 9.2000 ;
	    RECT 138.5000 8.8000 139.4000 9.2000 ;
	    RECT 140.9000 8.8000 141.8000 9.2000 ;
	    RECT 136.1000 8.2000 136.5000 8.8000 ;
	    RECT 138.5000 8.2000 138.9000 8.8000 ;
	    RECT 140.9000 8.2000 141.3000 8.8000 ;
	    RECT 136.1000 7.9000 137.0000 8.2000 ;
	    RECT 138.5000 7.9000 139.4000 8.2000 ;
	    RECT 140.9000 7.9000 141.8000 8.2000 ;
	    RECT 135.8000 7.1000 136.2000 7.2000 ;
	    RECT 135.0000 6.8000 136.2000 7.1000 ;
	    RECT 135.0000 1.1000 135.4000 6.8000 ;
	    RECT 135.8000 4.4000 136.2000 5.2000 ;
	    RECT 136.6000 1.1000 137.0000 7.9000 ;
	    RECT 137.4000 7.1000 137.8000 7.6000 ;
	    RECT 138.2000 7.1000 138.6000 7.2000 ;
	    RECT 137.4000 6.8000 138.6000 7.1000 ;
	    RECT 139.0000 1.1000 139.4000 7.9000 ;
	    RECT 139.8000 6.8000 140.2000 7.6000 ;
	    RECT 141.4000 1.1000 141.8000 7.9000 ;
	    RECT 142.2000 6.8000 142.6000 7.6000 ;
	    RECT 143.8000 5.1000 144.2000 9.9000 ;
	    RECT 144.9000 9.2000 145.3000 9.9000 ;
	    RECT 144.6000 8.8000 145.3000 9.2000 ;
	    RECT 144.9000 8.2000 145.3000 8.8000 ;
	    RECT 147.3000 9.2000 147.7000 9.9000 ;
	    RECT 149.7000 9.2000 150.1000 9.9000 ;
	    RECT 147.3000 8.8000 148.2000 9.2000 ;
	    RECT 149.7000 8.8000 150.6000 9.2000 ;
	    RECT 152.6000 8.9000 153.0000 9.9000 ;
	    RECT 147.3000 8.2000 147.7000 8.8000 ;
	    RECT 149.7000 8.2000 150.1000 8.8000 ;
	    RECT 144.9000 7.9000 145.8000 8.2000 ;
	    RECT 147.3000 7.9000 148.2000 8.2000 ;
	    RECT 149.7000 7.9000 150.6000 8.2000 ;
	    RECT 144.6000 5.1000 145.0000 5.2000 ;
	    RECT 143.8000 4.8000 145.0000 5.1000 ;
	    RECT 143.8000 1.1000 144.2000 4.8000 ;
	    RECT 144.6000 4.4000 145.0000 4.8000 ;
	    RECT 145.4000 1.1000 145.8000 7.9000 ;
	    RECT 146.2000 6.8000 146.6000 7.6000 ;
	    RECT 147.8000 1.1000 148.2000 7.9000 ;
	    RECT 148.6000 6.8000 149.0000 7.6000 ;
	    RECT 149.4000 4.4000 149.8000 5.2000 ;
	    RECT 150.2000 1.1000 150.6000 7.9000 ;
	    RECT 151.8000 7.8000 152.2000 8.6000 ;
	    RECT 152.7000 7.8000 153.0000 8.9000 ;
	    RECT 154.2000 7.9000 154.6000 9.9000 ;
	    RECT 155.8000 8.9000 156.2000 9.9000 ;
	    RECT 151.0000 7.1000 151.4000 7.6000 ;
	    RECT 151.8000 7.1000 152.1000 7.8000 ;
	    RECT 152.7000 7.5000 153.9000 7.8000 ;
	    RECT 151.0000 6.8000 152.1000 7.1000 ;
	    RECT 153.6000 6.0000 153.9000 7.5000 ;
	    RECT 154.3000 6.2000 154.6000 7.9000 ;
	    RECT 155.0000 7.8000 155.4000 8.6000 ;
	    RECT 155.9000 7.8000 156.2000 8.9000 ;
	    RECT 157.4000 7.9000 157.8000 9.9000 ;
	    RECT 155.9000 7.5000 157.1000 7.8000 ;
	    RECT 153.5000 5.7000 153.9000 6.0000 ;
	    RECT 154.2000 5.8000 154.6000 6.2000 ;
	    RECT 156.8000 6.0000 157.1000 7.5000 ;
	    RECT 157.5000 6.2000 157.8000 7.9000 ;
	    RECT 151.8000 5.6000 153.9000 5.7000 ;
	    RECT 151.8000 5.4000 153.8000 5.6000 ;
	    RECT 151.8000 1.1000 152.2000 5.4000 ;
	    RECT 154.3000 5.1000 154.6000 5.8000 ;
	    RECT 156.7000 5.7000 157.1000 6.0000 ;
	    RECT 157.4000 5.8000 157.8000 6.2000 ;
	    RECT 153.9000 4.8000 154.6000 5.1000 ;
	    RECT 155.0000 5.6000 157.1000 5.7000 ;
	    RECT 155.0000 5.4000 157.0000 5.6000 ;
	    RECT 153.9000 1.1000 154.3000 4.8000 ;
	    RECT 155.0000 1.1000 155.4000 5.4000 ;
	    RECT 157.5000 5.1000 157.8000 5.8000 ;
	    RECT 157.1000 4.8000 157.8000 5.1000 ;
	    RECT 157.1000 1.1000 157.5000 4.8000 ;
	    RECT 158.2000 1.1000 158.6000 9.9000 ;
	    RECT 160.6000 7.6000 161.0000 9.9000 ;
	    RECT 162.2000 7.6000 162.6000 9.9000 ;
	    RECT 163.8000 7.6000 164.2000 9.9000 ;
	    RECT 165.4000 7.6000 165.8000 9.9000 ;
	    RECT 159.0000 6.8000 159.4000 7.6000 ;
	    RECT 159.8000 7.2000 161.0000 7.6000 ;
	    RECT 161.5000 7.2000 162.6000 7.6000 ;
	    RECT 163.1000 7.2000 164.2000 7.6000 ;
	    RECT 164.9000 7.2000 165.8000 7.6000 ;
	    RECT 159.8000 5.8000 160.2000 7.2000 ;
	    RECT 161.5000 6.9000 161.9000 7.2000 ;
	    RECT 163.1000 6.9000 163.5000 7.2000 ;
	    RECT 164.9000 6.9000 165.3000 7.2000 ;
	    RECT 160.6000 6.5000 161.9000 6.9000 ;
	    RECT 162.3000 6.5000 163.5000 6.9000 ;
	    RECT 164.0000 6.5000 165.3000 6.9000 ;
	    RECT 161.5000 5.8000 161.9000 6.5000 ;
	    RECT 163.1000 5.8000 163.5000 6.5000 ;
	    RECT 164.9000 5.8000 165.3000 6.5000 ;
	    RECT 167.0000 6.2000 167.4000 9.9000 ;
	    RECT 168.6000 7.6000 169.0000 9.9000 ;
	    RECT 169.4000 7.9000 169.8000 9.9000 ;
	    RECT 171.5000 9.2000 171.9000 9.9000 ;
	    RECT 171.5000 8.8000 172.2000 9.2000 ;
	    RECT 171.5000 8.4000 171.9000 8.8000 ;
	    RECT 171.5000 7.9000 172.2000 8.4000 ;
	    RECT 167.9000 7.3000 169.0000 7.6000 ;
	    RECT 169.5000 7.8000 169.8000 7.9000 ;
	    RECT 169.5000 7.6000 170.4000 7.8000 ;
	    RECT 169.5000 7.5000 171.6000 7.6000 ;
	    RECT 170.1000 7.3000 171.6000 7.5000 ;
	    RECT 159.8000 5.4000 161.0000 5.8000 ;
	    RECT 161.5000 5.4000 162.6000 5.8000 ;
	    RECT 163.1000 5.4000 164.2000 5.8000 ;
	    RECT 164.9000 5.4000 165.8000 5.8000 ;
	    RECT 160.6000 1.1000 161.0000 5.4000 ;
	    RECT 162.2000 1.1000 162.6000 5.4000 ;
	    RECT 163.8000 1.1000 164.2000 5.4000 ;
	    RECT 165.4000 1.1000 165.8000 5.4000 ;
	    RECT 167.0000 5.1000 167.3000 6.2000 ;
	    RECT 167.9000 5.8000 168.2000 7.3000 ;
	    RECT 171.2000 7.2000 171.6000 7.3000 ;
	    RECT 169.4000 6.4000 169.8000 7.2000 ;
	    RECT 170.2000 6.6000 170.8000 7.0000 ;
	    RECT 170.3000 6.2000 170.6000 6.6000 ;
	    RECT 170.2000 5.8000 170.6000 6.2000 ;
	    RECT 167.6000 5.4000 168.2000 5.8000 ;
	    RECT 171.2000 5.5000 171.5000 7.2000 ;
	    RECT 171.9000 6.2000 172.2000 7.9000 ;
	    RECT 171.8000 5.8000 172.2000 6.2000 ;
	    RECT 167.9000 5.1000 168.2000 5.4000 ;
	    RECT 170.3000 5.2000 171.5000 5.5000 ;
	    RECT 167.0000 1.1000 167.4000 5.1000 ;
	    RECT 167.9000 4.8000 169.0000 5.1000 ;
	    RECT 168.6000 1.1000 169.0000 4.8000 ;
	    RECT 170.3000 3.1000 170.6000 5.2000 ;
	    RECT 171.9000 5.1000 172.2000 5.8000 ;
	    RECT 170.2000 1.1000 170.6000 3.1000 ;
	    RECT 171.8000 1.1000 172.2000 5.1000 ;
         LAYER metal2 ;
	    RECT 80.6000 156.8000 81.0000 157.2000 ;
	    RECT 49.4000 155.8000 49.8000 156.2000 ;
	    RECT 61.4000 155.8000 61.8000 156.2000 ;
	    RECT 62.2000 155.8000 62.6000 156.2000 ;
	    RECT 69.4000 156.1000 69.8000 156.2000 ;
	    RECT 70.2000 156.1000 70.6000 156.2000 ;
	    RECT 69.4000 155.8000 70.6000 156.1000 ;
	    RECT 75.8000 155.8000 76.2000 156.2000 ;
	    RECT 78.2000 156.1000 78.6000 156.2000 ;
	    RECT 79.0000 156.1000 79.4000 156.2000 ;
	    RECT 78.2000 155.8000 79.4000 156.1000 ;
	    RECT 9.4000 154.8000 9.8000 155.2000 ;
	    RECT 33.4000 154.8000 33.8000 155.2000 ;
	    RECT 39.8000 154.8000 40.2000 155.2000 ;
	    RECT 9.4000 154.2000 9.7000 154.8000 ;
	    RECT 4.6000 153.8000 5.0000 154.2000 ;
	    RECT 9.4000 153.8000 9.8000 154.2000 ;
	    RECT 11.8000 153.8000 12.2000 154.2000 ;
	    RECT 12.6000 154.1000 13.0000 154.2000 ;
	    RECT 13.4000 154.1000 13.8000 154.2000 ;
	    RECT 12.6000 153.8000 13.8000 154.1000 ;
	    RECT 14.2000 153.8000 14.6000 154.2000 ;
	    RECT 15.8000 154.1000 16.2000 154.2000 ;
	    RECT 16.6000 154.1000 17.0000 154.2000 ;
	    RECT 15.8000 153.8000 17.0000 154.1000 ;
	    RECT 18.2000 154.1000 18.6000 154.2000 ;
	    RECT 19.0000 154.1000 19.4000 154.2000 ;
	    RECT 18.2000 153.8000 19.4000 154.1000 ;
	    RECT 21.4000 154.1000 21.8000 154.2000 ;
	    RECT 22.2000 154.1000 22.6000 154.2000 ;
	    RECT 21.4000 153.8000 22.6000 154.1000 ;
	    RECT 25.4000 154.1000 25.8000 154.2000 ;
	    RECT 27.8000 154.1000 28.2000 154.2000 ;
	    RECT 28.6000 154.1000 29.0000 154.2000 ;
	    RECT 25.4000 153.8000 26.5000 154.1000 ;
	    RECT 27.8000 153.8000 29.0000 154.1000 ;
	    RECT 31.8000 154.1000 32.2000 154.2000 ;
	    RECT 32.6000 154.1000 33.0000 154.2000 ;
	    RECT 31.8000 153.8000 33.0000 154.1000 ;
	    RECT 2.2000 151.8000 2.6000 152.2000 ;
	    RECT 2.2000 147.1000 2.5000 151.8000 ;
	    RECT 1.4000 146.8000 2.5000 147.1000 ;
	    RECT 3.8000 146.8000 4.2000 147.2000 ;
	    RECT 1.4000 144.2000 1.7000 146.8000 ;
	    RECT 3.8000 146.2000 4.1000 146.8000 ;
	    RECT 4.6000 146.2000 4.9000 153.8000 ;
	    RECT 6.2000 151.8000 6.6000 152.2000 ;
	    RECT 6.2000 149.2000 6.5000 151.8000 ;
	    RECT 6.2000 148.8000 6.6000 149.2000 ;
	    RECT 11.8000 148.2000 12.1000 153.8000 ;
	    RECT 6.2000 147.8000 6.6000 148.2000 ;
	    RECT 11.8000 147.8000 12.2000 148.2000 ;
	    RECT 6.2000 146.2000 6.5000 147.8000 ;
	    RECT 7.0000 146.8000 7.4000 147.2000 ;
	    RECT 13.4000 146.8000 13.8000 147.2000 ;
	    RECT 7.0000 146.2000 7.3000 146.8000 ;
	    RECT 13.4000 146.2000 13.7000 146.8000 ;
	    RECT 14.2000 146.2000 14.5000 153.8000 ;
	    RECT 15.0000 151.8000 15.4000 152.2000 ;
	    RECT 20.6000 151.8000 21.0000 152.2000 ;
	    RECT 22.2000 151.8000 22.6000 152.2000 ;
	    RECT 2.2000 146.1000 2.6000 146.2000 ;
	    RECT 3.0000 146.1000 3.4000 146.2000 ;
	    RECT 2.2000 145.8000 3.4000 146.1000 ;
	    RECT 3.8000 145.8000 4.2000 146.2000 ;
	    RECT 4.6000 145.8000 5.0000 146.2000 ;
	    RECT 6.2000 145.8000 6.6000 146.2000 ;
	    RECT 7.0000 145.8000 7.4000 146.2000 ;
	    RECT 7.8000 146.1000 8.2000 146.2000 ;
	    RECT 8.6000 146.1000 9.0000 146.2000 ;
	    RECT 7.8000 145.8000 9.0000 146.1000 ;
	    RECT 13.4000 145.8000 13.8000 146.2000 ;
	    RECT 14.2000 145.8000 14.6000 146.2000 ;
	    RECT 3.0000 144.8000 3.4000 145.2000 ;
	    RECT 1.4000 143.8000 1.8000 144.2000 ;
	    RECT 2.2000 141.8000 2.6000 142.2000 ;
	    RECT 2.2000 140.2000 2.5000 141.8000 ;
	    RECT 3.0000 141.2000 3.3000 144.8000 ;
	    RECT 3.0000 140.8000 3.4000 141.2000 ;
	    RECT 2.2000 139.8000 2.6000 140.2000 ;
	    RECT 3.8000 139.8000 4.2000 140.2000 ;
	    RECT 2.2000 138.8000 2.6000 139.2000 ;
	    RECT 2.2000 138.2000 2.5000 138.8000 ;
	    RECT 2.2000 137.8000 2.6000 138.2000 ;
	    RECT 3.8000 133.1000 4.1000 139.8000 ;
	    RECT 5.4000 138.1000 5.8000 138.2000 ;
	    RECT 6.2000 138.1000 6.5000 145.8000 ;
	    RECT 7.0000 144.8000 7.4000 145.2000 ;
	    RECT 14.2000 145.1000 14.6000 145.2000 ;
	    RECT 15.0000 145.1000 15.3000 151.8000 ;
	    RECT 19.0000 147.8000 19.4000 148.2000 ;
	    RECT 15.8000 146.8000 16.2000 147.2000 ;
	    RECT 16.6000 147.1000 17.0000 147.2000 ;
	    RECT 17.4000 147.1000 17.8000 147.2000 ;
	    RECT 16.6000 146.8000 17.8000 147.1000 ;
	    RECT 18.2000 146.8000 18.6000 147.2000 ;
	    RECT 15.8000 146.2000 16.1000 146.8000 ;
	    RECT 18.2000 146.2000 18.5000 146.8000 ;
	    RECT 15.8000 145.8000 16.2000 146.2000 ;
	    RECT 18.2000 145.8000 18.6000 146.2000 ;
	    RECT 14.2000 144.8000 15.3000 145.1000 ;
	    RECT 7.0000 144.2000 7.3000 144.8000 ;
	    RECT 7.0000 143.8000 7.4000 144.2000 ;
	    RECT 15.8000 141.8000 16.2000 142.2000 ;
	    RECT 17.4000 141.8000 17.8000 142.2000 ;
	    RECT 5.4000 137.8000 6.5000 138.1000 ;
	    RECT 8.6000 140.8000 9.0000 141.2000 ;
	    RECT 4.6000 136.8000 5.0000 137.2000 ;
	    RECT 4.6000 136.2000 4.9000 136.8000 ;
	    RECT 4.6000 135.8000 5.0000 136.2000 ;
	    RECT 5.4000 135.2000 5.7000 137.8000 ;
	    RECT 8.6000 136.2000 8.9000 140.8000 ;
	    RECT 13.4000 137.8000 13.8000 138.2000 ;
	    RECT 10.2000 137.1000 10.6000 137.2000 ;
	    RECT 11.0000 137.1000 11.4000 137.2000 ;
	    RECT 10.2000 136.8000 11.4000 137.1000 ;
	    RECT 11.8000 136.8000 12.2000 137.2000 ;
	    RECT 12.6000 136.8000 13.0000 137.2000 ;
	    RECT 11.8000 136.2000 12.1000 136.8000 ;
	    RECT 8.6000 135.8000 9.0000 136.2000 ;
	    RECT 11.8000 135.8000 12.2000 136.2000 ;
	    RECT 5.4000 134.8000 5.8000 135.2000 ;
	    RECT 5.4000 133.2000 5.7000 134.8000 ;
	    RECT 7.8000 133.8000 8.2000 134.2000 ;
	    RECT 7.8000 133.2000 8.1000 133.8000 ;
	    RECT 3.8000 132.8000 4.9000 133.1000 ;
	    RECT 5.4000 132.8000 5.8000 133.2000 ;
	    RECT 7.8000 132.8000 8.2000 133.2000 ;
	    RECT 3.8000 131.8000 4.2000 132.2000 ;
	    RECT 1.4000 129.8000 1.8000 130.2000 ;
	    RECT 1.4000 129.2000 1.7000 129.8000 ;
	    RECT 1.4000 128.8000 1.8000 129.2000 ;
	    RECT 3.8000 124.2000 4.1000 131.8000 ;
	    RECT 4.6000 126.2000 4.9000 132.8000 ;
	    RECT 8.6000 130.2000 8.9000 135.8000 ;
	    RECT 9.4000 134.8000 9.8000 135.2000 ;
	    RECT 11.8000 134.8000 12.2000 135.2000 ;
	    RECT 9.4000 134.2000 9.7000 134.8000 ;
	    RECT 11.8000 134.2000 12.1000 134.8000 ;
	    RECT 9.4000 133.8000 9.8000 134.2000 ;
	    RECT 11.8000 133.8000 12.2000 134.2000 ;
	    RECT 9.4000 131.8000 9.8000 132.2000 ;
	    RECT 8.6000 129.8000 9.0000 130.2000 ;
	    RECT 9.4000 126.2000 9.7000 131.8000 ;
	    RECT 10.2000 127.8000 10.6000 128.2000 ;
	    RECT 4.6000 125.8000 5.0000 126.2000 ;
	    RECT 9.4000 125.8000 9.8000 126.2000 ;
	    RECT 10.2000 124.2000 10.5000 127.8000 ;
	    RECT 12.6000 126.2000 12.9000 136.8000 ;
	    RECT 13.4000 136.2000 13.7000 137.8000 ;
	    RECT 15.8000 136.2000 16.1000 141.8000 ;
	    RECT 13.4000 135.8000 13.8000 136.2000 ;
	    RECT 14.2000 136.1000 14.6000 136.2000 ;
	    RECT 15.0000 136.1000 15.4000 136.2000 ;
	    RECT 14.2000 135.8000 15.4000 136.1000 ;
	    RECT 15.8000 135.8000 16.2000 136.2000 ;
	    RECT 16.6000 136.1000 17.0000 136.2000 ;
	    RECT 17.4000 136.1000 17.7000 141.8000 ;
	    RECT 16.6000 135.8000 17.7000 136.1000 ;
	    RECT 19.0000 136.2000 19.3000 147.8000 ;
	    RECT 20.6000 145.2000 20.9000 151.8000 ;
	    RECT 21.4000 146.8000 21.8000 147.2000 ;
	    RECT 21.4000 146.2000 21.7000 146.8000 ;
	    RECT 21.4000 145.8000 21.8000 146.2000 ;
	    RECT 19.8000 144.8000 20.2000 145.2000 ;
	    RECT 20.6000 144.8000 21.0000 145.2000 ;
	    RECT 19.8000 141.2000 20.1000 144.8000 ;
	    RECT 22.2000 144.2000 22.5000 151.8000 ;
	    RECT 26.2000 148.2000 26.5000 153.8000 ;
	    RECT 33.4000 153.2000 33.7000 154.8000 ;
	    RECT 39.8000 154.2000 40.1000 154.8000 ;
	    RECT 49.4000 154.2000 49.7000 155.8000 ;
	    RECT 51.8000 154.8000 52.2000 155.2000 ;
	    RECT 55.8000 154.8000 56.2000 155.2000 ;
	    RECT 58.2000 155.1000 58.6000 155.2000 ;
	    RECT 59.0000 155.1000 59.4000 155.2000 ;
	    RECT 58.2000 154.8000 59.4000 155.1000 ;
	    RECT 60.6000 154.8000 61.0000 155.2000 ;
	    RECT 51.8000 154.2000 52.1000 154.8000 ;
	    RECT 55.8000 154.2000 56.1000 154.8000 ;
	    RECT 35.0000 154.1000 35.4000 154.2000 ;
	    RECT 35.8000 154.1000 36.2000 154.2000 ;
	    RECT 35.0000 153.8000 36.2000 154.1000 ;
	    RECT 37.4000 154.1000 37.8000 154.2000 ;
	    RECT 38.2000 154.1000 38.6000 154.2000 ;
	    RECT 37.4000 153.8000 38.6000 154.1000 ;
	    RECT 39.8000 153.8000 40.2000 154.2000 ;
	    RECT 40.6000 153.8000 41.0000 154.2000 ;
	    RECT 42.2000 154.1000 42.6000 154.2000 ;
	    RECT 43.0000 154.1000 43.4000 154.2000 ;
	    RECT 42.2000 153.8000 43.4000 154.1000 ;
	    RECT 44.6000 154.1000 45.0000 154.2000 ;
	    RECT 45.4000 154.1000 45.8000 154.2000 ;
	    RECT 44.6000 153.8000 45.8000 154.1000 ;
	    RECT 49.4000 153.8000 49.8000 154.2000 ;
	    RECT 51.8000 153.8000 52.2000 154.2000 ;
	    RECT 55.8000 153.8000 56.2000 154.2000 ;
	    RECT 33.4000 152.8000 33.8000 153.2000 ;
	    RECT 27.0000 151.8000 27.4000 152.2000 ;
	    RECT 29.4000 151.8000 29.8000 152.2000 ;
	    RECT 31.8000 151.8000 32.2000 152.2000 ;
	    RECT 39.0000 151.8000 39.4000 152.2000 ;
	    RECT 26.2000 147.8000 26.6000 148.2000 ;
	    RECT 23.8000 147.1000 24.2000 147.2000 ;
	    RECT 24.6000 147.1000 25.0000 147.2000 ;
	    RECT 23.8000 146.8000 25.0000 147.1000 ;
	    RECT 26.2000 146.2000 26.5000 147.8000 ;
	    RECT 26.2000 145.8000 26.6000 146.2000 ;
	    RECT 27.0000 145.2000 27.3000 151.8000 ;
	    RECT 29.4000 147.2000 29.7000 151.8000 ;
	    RECT 31.8000 147.2000 32.1000 151.8000 ;
	    RECT 29.4000 146.8000 29.8000 147.2000 ;
	    RECT 31.8000 146.8000 32.2000 147.2000 ;
	    RECT 35.0000 147.1000 35.4000 147.2000 ;
	    RECT 35.8000 147.1000 36.2000 147.2000 ;
	    RECT 35.0000 146.8000 36.2000 147.1000 ;
	    RECT 27.8000 146.1000 28.2000 146.2000 ;
	    RECT 28.6000 146.1000 29.0000 146.2000 ;
	    RECT 27.8000 145.8000 29.0000 146.1000 ;
	    RECT 33.4000 145.8000 33.8000 146.2000 ;
	    RECT 37.4000 146.1000 37.8000 146.2000 ;
	    RECT 38.2000 146.1000 38.6000 146.2000 ;
	    RECT 37.4000 145.8000 38.6000 146.1000 ;
	    RECT 27.0000 144.8000 27.4000 145.2000 ;
	    RECT 31.0000 145.1000 31.4000 145.2000 ;
	    RECT 31.8000 145.1000 32.2000 145.2000 ;
	    RECT 31.0000 144.8000 32.2000 145.1000 ;
	    RECT 22.2000 143.8000 22.6000 144.2000 ;
	    RECT 33.4000 143.2000 33.7000 145.8000 ;
	    RECT 39.0000 145.2000 39.3000 151.8000 ;
	    RECT 39.8000 149.2000 40.1000 153.8000 ;
	    RECT 40.6000 153.2000 40.9000 153.8000 ;
	    RECT 40.6000 152.8000 41.0000 153.2000 ;
	    RECT 43.8000 151.8000 44.2000 152.2000 ;
	    RECT 39.8000 148.8000 40.2000 149.2000 ;
	    RECT 39.8000 146.2000 40.1000 148.8000 ;
	    RECT 39.8000 145.8000 40.2000 146.2000 ;
	    RECT 39.0000 144.8000 39.4000 145.2000 ;
	    RECT 29.4000 142.8000 29.8000 143.2000 ;
	    RECT 33.4000 142.8000 33.8000 143.2000 ;
	    RECT 21.4000 141.8000 21.8000 142.2000 ;
	    RECT 28.6000 141.8000 29.0000 142.2000 ;
	    RECT 19.8000 140.8000 20.2000 141.2000 ;
	    RECT 21.4000 137.2000 21.7000 141.8000 ;
	    RECT 28.6000 139.2000 28.9000 141.8000 ;
	    RECT 23.0000 138.8000 23.4000 139.2000 ;
	    RECT 28.6000 138.8000 29.0000 139.2000 ;
	    RECT 21.4000 136.8000 21.8000 137.2000 ;
	    RECT 23.0000 136.2000 23.3000 138.8000 ;
	    RECT 26.2000 137.8000 26.6000 138.2000 ;
	    RECT 26.2000 137.2000 26.5000 137.8000 ;
	    RECT 26.2000 136.8000 26.6000 137.2000 ;
	    RECT 19.0000 135.8000 19.4000 136.2000 ;
	    RECT 23.0000 135.8000 23.4000 136.2000 ;
	    RECT 27.8000 136.1000 28.2000 136.2000 ;
	    RECT 28.6000 136.1000 29.0000 136.2000 ;
	    RECT 27.8000 135.8000 29.0000 136.1000 ;
	    RECT 29.4000 135.2000 29.7000 142.8000 ;
	    RECT 30.2000 141.8000 30.6000 142.2000 ;
	    RECT 33.4000 141.8000 33.8000 142.2000 ;
	    RECT 37.4000 141.8000 37.8000 142.2000 ;
	    RECT 30.2000 136.2000 30.5000 141.8000 ;
	    RECT 33.4000 136.2000 33.7000 141.8000 ;
	    RECT 37.4000 140.2000 37.7000 141.8000 ;
	    RECT 37.4000 139.8000 37.8000 140.2000 ;
	    RECT 30.2000 135.8000 30.6000 136.2000 ;
	    RECT 31.8000 136.1000 32.2000 136.2000 ;
	    RECT 32.6000 136.1000 33.0000 136.2000 ;
	    RECT 31.8000 135.8000 33.0000 136.1000 ;
	    RECT 33.4000 135.8000 33.8000 136.2000 ;
	    RECT 37.4000 136.1000 37.8000 136.2000 ;
	    RECT 38.2000 136.1000 38.6000 136.2000 ;
	    RECT 37.4000 135.8000 38.6000 136.1000 ;
	    RECT 39.8000 135.2000 40.1000 145.8000 ;
	    RECT 43.8000 145.2000 44.1000 151.8000 ;
	    RECT 44.6000 148.2000 44.9000 153.8000 ;
	    RECT 46.2000 152.1000 46.6000 152.2000 ;
	    RECT 47.0000 152.1000 47.4000 152.2000 ;
	    RECT 46.2000 151.8000 47.4000 152.1000 ;
	    RECT 50.2000 151.8000 50.6000 152.2000 ;
	    RECT 51.8000 151.8000 52.2000 152.2000 ;
	    RECT 52.6000 152.1000 53.0000 152.2000 ;
	    RECT 53.4000 152.1000 53.8000 152.2000 ;
	    RECT 52.6000 151.8000 53.8000 152.1000 ;
	    RECT 50.2000 151.2000 50.5000 151.8000 ;
	    RECT 50.2000 150.8000 50.6000 151.2000 ;
	    RECT 44.6000 147.8000 45.0000 148.2000 ;
	    RECT 46.2000 148.1000 46.6000 148.2000 ;
	    RECT 47.0000 148.1000 47.4000 148.2000 ;
	    RECT 46.2000 147.8000 47.4000 148.1000 ;
	    RECT 44.6000 146.2000 44.9000 147.8000 ;
	    RECT 50.2000 146.8000 50.6000 147.2000 ;
	    RECT 50.2000 146.2000 50.5000 146.8000 ;
	    RECT 44.6000 145.8000 45.0000 146.2000 ;
	    RECT 46.2000 145.8000 46.6000 146.2000 ;
	    RECT 50.2000 145.8000 50.6000 146.2000 ;
	    RECT 46.2000 145.2000 46.5000 145.8000 ;
	    RECT 43.8000 144.8000 44.2000 145.2000 ;
	    RECT 46.2000 144.8000 46.6000 145.2000 ;
	    RECT 51.8000 144.1000 52.1000 151.8000 ;
	    RECT 57.4000 150.8000 57.8000 151.2000 ;
	    RECT 53.4000 147.8000 53.8000 148.2000 ;
	    RECT 53.4000 147.2000 53.7000 147.8000 ;
	    RECT 53.4000 146.8000 53.8000 147.2000 ;
	    RECT 52.6000 146.1000 53.0000 146.2000 ;
	    RECT 53.4000 146.1000 53.8000 146.2000 ;
	    RECT 52.6000 145.8000 53.8000 146.1000 ;
	    RECT 55.0000 145.1000 55.4000 145.2000 ;
	    RECT 55.8000 145.1000 56.2000 145.2000 ;
	    RECT 55.0000 144.8000 56.2000 145.1000 ;
	    RECT 57.4000 144.2000 57.7000 150.8000 ;
	    RECT 60.6000 148.2000 60.9000 154.8000 ;
	    RECT 61.4000 154.2000 61.7000 155.8000 ;
	    RECT 62.2000 155.2000 62.5000 155.8000 ;
	    RECT 75.8000 155.2000 76.1000 155.8000 ;
	    RECT 80.6000 155.2000 80.9000 156.8000 ;
	    RECT 62.2000 154.8000 62.6000 155.2000 ;
	    RECT 64.6000 154.8000 65.0000 155.2000 ;
	    RECT 71.8000 154.8000 72.2000 155.2000 ;
	    RECT 75.8000 154.8000 76.2000 155.2000 ;
	    RECT 77.4000 154.8000 77.8000 155.2000 ;
	    RECT 80.6000 154.8000 81.0000 155.2000 ;
	    RECT 64.6000 154.2000 64.9000 154.8000 ;
	    RECT 71.8000 154.2000 72.1000 154.8000 ;
	    RECT 61.4000 153.8000 61.8000 154.2000 ;
	    RECT 64.6000 153.8000 65.0000 154.2000 ;
	    RECT 71.8000 153.8000 72.2000 154.2000 ;
	    RECT 66.2000 151.8000 66.6000 152.2000 ;
	    RECT 69.4000 151.8000 69.8000 152.2000 ;
	    RECT 60.6000 147.8000 61.0000 148.2000 ;
	    RECT 58.2000 146.8000 58.6000 147.2000 ;
	    RECT 63.8000 147.1000 64.2000 147.2000 ;
	    RECT 64.6000 147.1000 65.0000 147.2000 ;
	    RECT 63.8000 146.8000 65.0000 147.1000 ;
	    RECT 65.4000 146.8000 65.8000 147.2000 ;
	    RECT 58.2000 146.2000 58.5000 146.8000 ;
	    RECT 65.4000 146.2000 65.7000 146.8000 ;
	    RECT 58.2000 145.8000 58.6000 146.2000 ;
	    RECT 65.4000 145.8000 65.8000 146.2000 ;
	    RECT 64.6000 144.8000 65.0000 145.2000 ;
	    RECT 64.6000 144.2000 64.9000 144.8000 ;
	    RECT 66.2000 144.2000 66.5000 151.8000 ;
	    RECT 67.0000 147.8000 67.4000 148.2000 ;
	    RECT 67.0000 147.2000 67.3000 147.8000 ;
	    RECT 67.0000 146.8000 67.4000 147.2000 ;
	    RECT 68.6000 146.8000 69.0000 147.2000 ;
	    RECT 68.6000 146.2000 68.9000 146.8000 ;
	    RECT 68.6000 145.8000 69.0000 146.2000 ;
	    RECT 69.4000 144.2000 69.7000 151.8000 ;
	    RECT 52.6000 144.1000 53.0000 144.2000 ;
	    RECT 51.8000 143.8000 53.0000 144.1000 ;
	    RECT 57.4000 143.8000 57.8000 144.2000 ;
	    RECT 64.6000 143.8000 65.0000 144.2000 ;
	    RECT 66.2000 143.8000 66.6000 144.2000 ;
	    RECT 69.4000 143.8000 69.8000 144.2000 ;
	    RECT 44.6000 142.8000 45.0000 143.2000 ;
	    RECT 71.8000 143.1000 72.1000 153.8000 ;
	    RECT 77.4000 153.2000 77.7000 154.8000 ;
	    RECT 75.8000 152.8000 76.2000 153.2000 ;
	    RECT 77.4000 152.8000 77.8000 153.2000 ;
	    RECT 73.4000 151.8000 73.8000 152.2000 ;
	    RECT 73.4000 149.2000 73.7000 151.8000 ;
	    RECT 73.4000 148.8000 73.8000 149.2000 ;
	    RECT 75.8000 149.1000 76.1000 152.8000 ;
	    RECT 79.0000 151.8000 79.4000 152.2000 ;
	    RECT 83.0000 152.1000 83.4000 157.9000 ;
	    RECT 87.0000 154.7000 87.4000 155.1000 ;
	    RECT 85.4000 153.8000 85.8000 154.2000 ;
	    RECT 83.8000 152.8000 84.2000 153.2000 ;
	    RECT 75.0000 148.8000 76.1000 149.1000 ;
	    RECT 76.6000 148.8000 77.0000 149.2000 ;
	    RECT 77.4000 148.8000 77.8000 149.2000 ;
	    RECT 75.0000 148.2000 75.3000 148.8000 ;
	    RECT 72.6000 147.8000 73.0000 148.2000 ;
	    RECT 75.0000 147.8000 75.4000 148.2000 ;
	    RECT 75.8000 147.8000 76.2000 148.2000 ;
	    RECT 72.6000 146.2000 72.9000 147.8000 ;
	    RECT 75.8000 147.2000 76.1000 147.8000 ;
	    RECT 73.4000 147.1000 73.8000 147.2000 ;
	    RECT 74.2000 147.1000 74.6000 147.2000 ;
	    RECT 73.4000 146.8000 74.6000 147.1000 ;
	    RECT 75.0000 146.8000 75.4000 147.2000 ;
	    RECT 75.8000 146.8000 76.2000 147.2000 ;
	    RECT 75.0000 146.2000 75.3000 146.8000 ;
	    RECT 72.6000 145.8000 73.0000 146.2000 ;
	    RECT 75.0000 145.8000 75.4000 146.2000 ;
	    RECT 71.8000 142.8000 72.9000 143.1000 ;
	    RECT 44.6000 142.2000 44.9000 142.8000 ;
	    RECT 44.6000 141.8000 45.0000 142.2000 ;
	    RECT 51.0000 141.8000 51.4000 142.2000 ;
	    RECT 55.8000 141.8000 56.2000 142.2000 ;
	    RECT 58.2000 141.8000 58.6000 142.2000 ;
	    RECT 70.2000 141.8000 70.6000 142.2000 ;
	    RECT 71.8000 141.8000 72.2000 142.2000 ;
	    RECT 51.0000 140.1000 51.3000 141.8000 ;
	    RECT 51.0000 139.8000 52.1000 140.1000 ;
	    RECT 40.6000 136.8000 41.0000 137.2000 ;
	    RECT 40.6000 136.2000 40.9000 136.8000 ;
	    RECT 51.8000 136.2000 52.1000 139.8000 ;
	    RECT 55.0000 136.8000 55.4000 137.2000 ;
	    RECT 55.0000 136.2000 55.3000 136.8000 ;
	    RECT 40.6000 135.8000 41.0000 136.2000 ;
	    RECT 49.4000 135.8000 49.8000 136.2000 ;
	    RECT 51.8000 135.8000 52.2000 136.2000 ;
	    RECT 55.0000 135.8000 55.4000 136.2000 ;
	    RECT 18.2000 134.8000 18.6000 135.2000 ;
	    RECT 29.4000 134.8000 29.8000 135.2000 ;
	    RECT 39.8000 134.8000 40.2000 135.2000 ;
	    RECT 40.6000 134.8000 41.0000 135.2000 ;
	    RECT 43.8000 134.8000 44.2000 135.2000 ;
	    RECT 47.0000 135.1000 47.4000 135.2000 ;
	    RECT 47.8000 135.1000 48.2000 135.2000 ;
	    RECT 47.0000 134.8000 48.2000 135.1000 ;
	    RECT 18.2000 134.2000 18.5000 134.8000 ;
	    RECT 29.4000 134.2000 29.7000 134.8000 ;
	    RECT 18.2000 133.8000 18.6000 134.2000 ;
	    RECT 29.4000 133.8000 29.8000 134.2000 ;
	    RECT 32.6000 132.8000 33.0000 133.2000 ;
	    RECT 32.6000 132.2000 32.9000 132.8000 ;
	    RECT 40.6000 132.2000 40.9000 134.8000 ;
	    RECT 43.0000 133.8000 43.4000 134.2000 ;
	    RECT 43.0000 132.2000 43.3000 133.8000 ;
	    RECT 14.2000 131.8000 14.6000 132.2000 ;
	    RECT 16.6000 131.8000 17.0000 132.2000 ;
	    RECT 19.0000 131.8000 19.4000 132.2000 ;
	    RECT 22.2000 131.8000 22.6000 132.2000 ;
	    RECT 25.4000 131.8000 25.8000 132.2000 ;
	    RECT 28.6000 131.8000 29.0000 132.2000 ;
	    RECT 31.8000 131.8000 32.2000 132.2000 ;
	    RECT 32.6000 131.8000 33.0000 132.2000 ;
	    RECT 35.0000 131.8000 35.4000 132.2000 ;
	    RECT 36.6000 131.8000 37.0000 132.2000 ;
	    RECT 39.0000 131.8000 39.4000 132.2000 ;
	    RECT 40.6000 131.8000 41.0000 132.2000 ;
	    RECT 43.0000 131.8000 43.4000 132.2000 ;
	    RECT 12.6000 125.8000 13.0000 126.2000 ;
	    RECT 3.8000 123.8000 4.2000 124.2000 ;
	    RECT 10.2000 123.8000 10.6000 124.2000 ;
	    RECT 13.4000 124.1000 13.8000 124.2000 ;
	    RECT 14.2000 124.1000 14.5000 131.8000 ;
	    RECT 16.6000 127.1000 16.9000 131.8000 ;
	    RECT 13.4000 123.8000 14.5000 124.1000 ;
	    RECT 15.8000 126.8000 16.9000 127.1000 ;
	    RECT 15.8000 124.2000 16.1000 126.8000 ;
	    RECT 16.6000 126.1000 17.0000 126.2000 ;
	    RECT 17.4000 126.1000 17.8000 126.2000 ;
	    RECT 16.6000 125.8000 17.8000 126.1000 ;
	    RECT 17.4000 124.8000 17.8000 125.2000 ;
	    RECT 15.8000 123.8000 16.2000 124.2000 ;
	    RECT 16.6000 123.8000 17.0000 124.2000 ;
	    RECT 16.6000 123.2000 16.9000 123.8000 ;
	    RECT 16.6000 122.8000 17.0000 123.2000 ;
	    RECT 17.4000 122.2000 17.7000 124.8000 ;
	    RECT 19.0000 124.2000 19.3000 131.8000 ;
	    RECT 22.2000 128.2000 22.5000 131.8000 ;
	    RECT 22.2000 127.8000 22.6000 128.2000 ;
	    RECT 24.6000 128.1000 25.0000 128.2000 ;
	    RECT 25.4000 128.1000 25.7000 131.8000 ;
	    RECT 24.6000 127.8000 25.7000 128.1000 ;
	    RECT 21.4000 126.8000 21.8000 127.2000 ;
	    RECT 21.4000 126.2000 21.7000 126.8000 ;
	    RECT 19.8000 125.8000 20.2000 126.2000 ;
	    RECT 21.4000 125.8000 21.8000 126.2000 ;
	    RECT 19.8000 124.2000 20.1000 125.8000 ;
	    RECT 19.0000 123.8000 19.4000 124.2000 ;
	    RECT 19.8000 123.8000 20.2000 124.2000 ;
	    RECT 1.4000 121.8000 1.8000 122.2000 ;
	    RECT 4.6000 121.8000 5.0000 122.2000 ;
	    RECT 7.0000 121.8000 7.4000 122.2000 ;
	    RECT 11.0000 121.8000 11.4000 122.2000 ;
	    RECT 13.4000 121.8000 13.8000 122.2000 ;
	    RECT 14.2000 121.8000 14.6000 122.2000 ;
	    RECT 17.4000 121.8000 17.8000 122.2000 ;
	    RECT 19.8000 121.8000 20.2000 122.2000 ;
	    RECT 1.4000 121.2000 1.7000 121.8000 ;
	    RECT 1.4000 120.8000 1.8000 121.2000 ;
	    RECT 3.8000 113.8000 4.2000 114.2000 ;
	    RECT 3.8000 113.2000 4.1000 113.8000 ;
	    RECT 0.6000 113.1000 1.0000 113.2000 ;
	    RECT 1.4000 113.1000 1.8000 113.2000 ;
	    RECT 0.6000 112.8000 1.8000 113.1000 ;
	    RECT 2.2000 112.8000 2.6000 113.2000 ;
	    RECT 3.8000 112.8000 4.2000 113.2000 ;
	    RECT 0.6000 105.1000 1.0000 105.2000 ;
	    RECT 1.4000 105.1000 1.8000 105.2000 ;
	    RECT 0.6000 104.8000 1.8000 105.1000 ;
	    RECT 2.2000 99.2000 2.5000 112.8000 ;
	    RECT 3.0000 111.8000 3.4000 112.2000 ;
	    RECT 3.0000 106.2000 3.3000 111.8000 ;
	    RECT 3.0000 105.8000 3.4000 106.2000 ;
	    RECT 3.8000 105.8000 4.2000 106.2000 ;
	    RECT 3.0000 104.8000 3.4000 105.2000 ;
	    RECT 3.0000 103.2000 3.3000 104.8000 ;
	    RECT 3.8000 104.2000 4.1000 105.8000 ;
	    RECT 3.8000 103.8000 4.2000 104.2000 ;
	    RECT 3.0000 102.8000 3.4000 103.2000 ;
	    RECT 3.0000 101.8000 3.4000 102.2000 ;
	    RECT 2.2000 98.8000 2.6000 99.2000 ;
	    RECT 3.0000 94.1000 3.3000 101.8000 ;
	    RECT 3.0000 93.8000 4.1000 94.1000 ;
	    RECT 2.2000 91.8000 2.6000 92.2000 ;
	    RECT 2.2000 88.2000 2.5000 91.8000 ;
	    RECT 2.2000 87.8000 2.6000 88.2000 ;
	    RECT 2.2000 87.2000 2.5000 87.8000 ;
	    RECT 2.2000 86.8000 2.6000 87.2000 ;
	    RECT 0.6000 83.8000 1.0000 84.2000 ;
	    RECT 0.6000 76.2000 0.9000 83.8000 ;
	    RECT 0.6000 75.8000 1.0000 76.2000 ;
	    RECT 2.2000 74.2000 2.5000 86.8000 ;
	    RECT 3.8000 86.2000 4.1000 93.8000 ;
	    RECT 3.8000 85.8000 4.2000 86.2000 ;
	    RECT 3.0000 84.8000 3.4000 85.2000 ;
	    RECT 3.0000 84.2000 3.3000 84.8000 ;
	    RECT 3.0000 83.8000 3.4000 84.2000 ;
	    RECT 4.6000 77.2000 4.9000 121.8000 ;
	    RECT 7.0000 116.2000 7.3000 121.8000 ;
	    RECT 11.0000 118.2000 11.3000 121.8000 ;
	    RECT 11.0000 117.8000 11.4000 118.2000 ;
	    RECT 11.0000 116.8000 11.4000 117.2000 ;
	    RECT 11.8000 117.1000 12.2000 117.2000 ;
	    RECT 12.6000 117.1000 13.0000 117.2000 ;
	    RECT 11.8000 116.8000 13.0000 117.1000 ;
	    RECT 11.0000 116.2000 11.3000 116.8000 ;
	    RECT 13.4000 116.2000 13.7000 121.8000 ;
	    RECT 14.2000 116.2000 14.5000 121.8000 ;
	    RECT 19.8000 119.2000 20.1000 121.8000 ;
	    RECT 19.8000 118.8000 20.2000 119.2000 ;
	    RECT 7.0000 115.8000 7.4000 116.2000 ;
	    RECT 11.0000 115.8000 11.4000 116.2000 ;
	    RECT 12.6000 116.1000 13.0000 116.2000 ;
	    RECT 13.4000 116.1000 13.8000 116.2000 ;
	    RECT 12.6000 115.8000 13.8000 116.1000 ;
	    RECT 14.2000 115.8000 14.6000 116.2000 ;
	    RECT 13.4000 115.1000 13.8000 115.2000 ;
	    RECT 15.0000 115.1000 15.4000 115.2000 ;
	    RECT 13.4000 114.8000 15.4000 115.1000 ;
	    RECT 11.0000 113.8000 11.4000 114.2000 ;
	    RECT 23.8000 113.8000 24.2000 114.2000 ;
	    RECT 11.0000 112.2000 11.3000 113.8000 ;
	    RECT 17.4000 112.8000 17.8000 113.2000 ;
	    RECT 17.4000 112.2000 17.7000 112.8000 ;
	    RECT 23.8000 112.2000 24.1000 113.8000 ;
	    RECT 24.6000 113.2000 24.9000 127.8000 ;
	    RECT 28.6000 127.2000 28.9000 131.8000 ;
	    RECT 29.4000 127.8000 29.8000 128.2000 ;
	    RECT 29.4000 127.2000 29.7000 127.8000 ;
	    RECT 27.0000 126.8000 27.4000 127.2000 ;
	    RECT 28.6000 126.8000 29.0000 127.2000 ;
	    RECT 29.4000 126.8000 29.8000 127.2000 ;
	    RECT 27.0000 126.2000 27.3000 126.8000 ;
	    RECT 27.0000 125.8000 27.4000 126.2000 ;
	    RECT 28.6000 126.1000 29.0000 126.2000 ;
	    RECT 29.4000 126.1000 29.8000 126.2000 ;
	    RECT 28.6000 125.8000 29.8000 126.1000 ;
	    RECT 30.2000 124.8000 30.6000 125.2000 ;
	    RECT 28.6000 124.1000 29.0000 124.2000 ;
	    RECT 29.4000 124.1000 29.8000 124.2000 ;
	    RECT 28.6000 123.8000 29.8000 124.1000 ;
	    RECT 30.2000 122.2000 30.5000 124.8000 ;
	    RECT 31.8000 124.2000 32.1000 131.8000 ;
	    RECT 32.6000 126.8000 33.0000 127.2000 ;
	    RECT 32.6000 126.2000 32.9000 126.8000 ;
	    RECT 35.0000 126.2000 35.3000 131.8000 ;
	    RECT 32.6000 125.8000 33.0000 126.2000 ;
	    RECT 35.0000 125.8000 35.4000 126.2000 ;
	    RECT 34.2000 124.8000 34.6000 125.2000 ;
	    RECT 31.8000 123.8000 32.2000 124.2000 ;
	    RECT 34.2000 122.2000 34.5000 124.8000 ;
	    RECT 35.8000 123.8000 36.2000 124.2000 ;
	    RECT 35.8000 123.2000 36.1000 123.8000 ;
	    RECT 35.8000 122.8000 36.2000 123.2000 ;
	    RECT 26.2000 121.8000 26.6000 122.2000 ;
	    RECT 30.2000 121.8000 30.6000 122.2000 ;
	    RECT 32.6000 121.8000 33.0000 122.2000 ;
	    RECT 34.2000 121.8000 34.6000 122.2000 ;
	    RECT 35.0000 121.8000 35.4000 122.2000 ;
	    RECT 24.6000 112.8000 25.0000 113.2000 ;
	    RECT 5.4000 111.8000 5.8000 112.2000 ;
	    RECT 11.0000 111.8000 11.4000 112.2000 ;
	    RECT 11.8000 111.8000 12.2000 112.2000 ;
	    RECT 13.4000 111.8000 13.8000 112.2000 ;
	    RECT 17.4000 111.8000 17.8000 112.2000 ;
	    RECT 19.8000 111.8000 20.2000 112.2000 ;
	    RECT 23.0000 111.8000 23.4000 112.2000 ;
	    RECT 23.8000 111.8000 24.2000 112.2000 ;
	    RECT 5.4000 106.2000 5.7000 111.8000 ;
	    RECT 7.0000 107.1000 7.4000 107.2000 ;
	    RECT 7.0000 106.8000 8.1000 107.1000 ;
	    RECT 5.4000 105.8000 5.8000 106.2000 ;
	    RECT 5.4000 104.8000 5.8000 105.2000 ;
	    RECT 7.0000 104.8000 7.4000 105.2000 ;
	    RECT 5.4000 104.2000 5.7000 104.8000 ;
	    RECT 7.0000 104.2000 7.3000 104.8000 ;
	    RECT 5.4000 103.8000 5.8000 104.2000 ;
	    RECT 7.0000 103.8000 7.4000 104.2000 ;
	    RECT 5.4000 96.8000 5.8000 97.2000 ;
	    RECT 5.4000 96.2000 5.7000 96.8000 ;
	    RECT 5.4000 95.8000 5.8000 96.2000 ;
	    RECT 7.8000 95.2000 8.1000 106.8000 ;
	    RECT 9.4000 106.8000 9.8000 107.2000 ;
	    RECT 11.0000 106.8000 11.4000 107.2000 ;
	    RECT 9.4000 106.2000 9.7000 106.8000 ;
	    RECT 11.0000 106.2000 11.3000 106.8000 ;
	    RECT 11.8000 106.2000 12.1000 111.8000 ;
	    RECT 13.4000 108.2000 13.7000 111.8000 ;
	    RECT 19.8000 108.2000 20.1000 111.8000 ;
	    RECT 13.4000 107.8000 13.8000 108.2000 ;
	    RECT 15.8000 107.8000 16.2000 108.2000 ;
	    RECT 19.8000 107.8000 20.2000 108.2000 ;
	    RECT 22.2000 107.8000 22.6000 108.2000 ;
	    RECT 15.8000 107.2000 16.1000 107.8000 ;
	    RECT 22.2000 107.2000 22.5000 107.8000 ;
	    RECT 15.8000 106.8000 16.2000 107.2000 ;
	    RECT 22.2000 106.8000 22.6000 107.2000 ;
	    RECT 9.4000 105.8000 9.8000 106.2000 ;
	    RECT 11.0000 105.8000 11.4000 106.2000 ;
	    RECT 11.8000 105.8000 12.2000 106.2000 ;
	    RECT 15.0000 106.1000 15.4000 106.2000 ;
	    RECT 15.8000 106.1000 16.2000 106.2000 ;
	    RECT 15.0000 105.8000 16.2000 106.1000 ;
	    RECT 22.2000 105.8000 22.6000 106.2000 ;
	    RECT 8.6000 104.8000 9.0000 105.2000 ;
	    RECT 16.6000 104.8000 17.0000 105.2000 ;
	    RECT 8.6000 104.2000 8.9000 104.8000 ;
	    RECT 16.6000 104.2000 16.9000 104.8000 ;
	    RECT 8.6000 103.8000 9.0000 104.2000 ;
	    RECT 9.4000 103.8000 9.8000 104.2000 ;
	    RECT 14.2000 104.1000 14.6000 104.2000 ;
	    RECT 15.0000 104.1000 15.4000 104.2000 ;
	    RECT 14.2000 103.8000 15.4000 104.1000 ;
	    RECT 15.8000 103.8000 16.2000 104.2000 ;
	    RECT 16.6000 103.8000 17.0000 104.2000 ;
	    RECT 9.4000 103.2000 9.7000 103.8000 ;
	    RECT 9.4000 102.8000 9.8000 103.2000 ;
	    RECT 10.2000 97.1000 10.6000 97.2000 ;
	    RECT 11.0000 97.1000 11.4000 97.2000 ;
	    RECT 10.2000 96.8000 11.4000 97.1000 ;
	    RECT 12.6000 96.1000 13.0000 96.2000 ;
	    RECT 13.4000 96.1000 13.8000 96.2000 ;
	    RECT 12.6000 95.8000 13.8000 96.1000 ;
	    RECT 15.8000 95.2000 16.1000 103.8000 ;
	    RECT 22.2000 99.2000 22.5000 105.8000 ;
	    RECT 23.0000 104.1000 23.3000 111.8000 ;
	    RECT 24.6000 106.8000 25.0000 107.2000 ;
	    RECT 24.6000 106.2000 24.9000 106.8000 ;
	    RECT 24.6000 105.8000 25.0000 106.2000 ;
	    RECT 25.4000 105.1000 25.8000 105.2000 ;
	    RECT 26.2000 105.1000 26.5000 121.8000 ;
	    RECT 31.8000 120.8000 32.2000 121.2000 ;
	    RECT 31.8000 119.2000 32.1000 120.8000 ;
	    RECT 31.8000 118.8000 32.2000 119.2000 ;
	    RECT 28.6000 116.8000 29.0000 117.2000 ;
	    RECT 29.4000 117.1000 29.8000 117.2000 ;
	    RECT 30.2000 117.1000 30.6000 117.2000 ;
	    RECT 29.4000 116.8000 30.6000 117.1000 ;
	    RECT 31.8000 116.8000 32.2000 117.2000 ;
	    RECT 28.6000 115.2000 28.9000 116.8000 ;
	    RECT 28.6000 114.8000 29.0000 115.2000 ;
	    RECT 29.4000 111.8000 29.8000 112.2000 ;
	    RECT 31.0000 111.8000 31.4000 112.2000 ;
	    RECT 27.8000 106.1000 28.2000 106.2000 ;
	    RECT 28.6000 106.1000 29.0000 106.2000 ;
	    RECT 27.8000 105.8000 29.0000 106.1000 ;
	    RECT 25.4000 104.8000 26.5000 105.1000 ;
	    RECT 27.8000 104.8000 28.2000 105.2000 ;
	    RECT 23.8000 104.1000 24.2000 104.2000 ;
	    RECT 23.0000 103.8000 24.2000 104.1000 ;
	    RECT 24.6000 101.8000 25.0000 102.2000 ;
	    RECT 22.2000 98.8000 22.6000 99.2000 ;
	    RECT 16.6000 97.1000 17.0000 97.2000 ;
	    RECT 17.4000 97.1000 17.8000 97.2000 ;
	    RECT 16.6000 96.8000 17.8000 97.1000 ;
	    RECT 20.6000 97.1000 21.0000 97.2000 ;
	    RECT 21.4000 97.1000 21.8000 97.2000 ;
	    RECT 20.6000 96.8000 21.8000 97.1000 ;
	    RECT 23.0000 96.8000 23.4000 97.2000 ;
	    RECT 23.0000 96.2000 23.3000 96.8000 ;
	    RECT 23.0000 95.8000 23.4000 96.2000 ;
	    RECT 24.6000 95.2000 24.9000 101.8000 ;
	    RECT 25.4000 96.2000 25.7000 104.8000 ;
	    RECT 27.8000 104.2000 28.1000 104.8000 ;
	    RECT 29.4000 104.2000 29.7000 111.8000 ;
	    RECT 31.0000 107.2000 31.3000 111.8000 ;
	    RECT 31.8000 109.2000 32.1000 116.8000 ;
	    RECT 32.6000 115.2000 32.9000 121.8000 ;
	    RECT 33.4000 117.1000 33.8000 117.2000 ;
	    RECT 34.2000 117.1000 34.6000 117.2000 ;
	    RECT 33.4000 116.8000 34.6000 117.1000 ;
	    RECT 35.0000 115.2000 35.3000 121.8000 ;
	    RECT 35.8000 117.1000 36.2000 117.2000 ;
	    RECT 36.6000 117.1000 36.9000 131.8000 ;
	    RECT 39.0000 127.2000 39.3000 131.8000 ;
	    RECT 43.8000 128.2000 44.1000 134.8000 ;
	    RECT 49.4000 134.2000 49.7000 135.8000 ;
	    RECT 55.8000 135.2000 56.1000 141.8000 ;
	    RECT 57.4000 139.8000 57.8000 140.2000 ;
	    RECT 56.6000 137.8000 57.0000 138.2000 ;
	    RECT 56.6000 137.2000 56.9000 137.8000 ;
	    RECT 56.6000 136.8000 57.0000 137.2000 ;
	    RECT 57.4000 136.1000 57.7000 139.8000 ;
	    RECT 58.2000 138.2000 58.5000 141.8000 ;
	    RECT 58.2000 137.8000 58.6000 138.2000 ;
	    RECT 67.8000 136.8000 68.2000 137.2000 ;
	    RECT 67.8000 136.2000 68.1000 136.8000 ;
	    RECT 58.2000 136.1000 58.6000 136.2000 ;
	    RECT 57.4000 135.8000 58.6000 136.1000 ;
	    RECT 61.4000 136.1000 61.8000 136.2000 ;
	    RECT 62.2000 136.1000 62.6000 136.2000 ;
	    RECT 61.4000 135.8000 62.6000 136.1000 ;
	    RECT 67.8000 135.8000 68.2000 136.2000 ;
	    RECT 70.2000 135.2000 70.5000 141.8000 ;
	    RECT 71.8000 136.2000 72.1000 141.8000 ;
	    RECT 71.8000 135.8000 72.2000 136.2000 ;
	    RECT 50.2000 134.8000 50.6000 135.2000 ;
	    RECT 55.8000 134.8000 56.2000 135.2000 ;
	    RECT 56.6000 134.8000 57.0000 135.2000 ;
	    RECT 57.4000 134.8000 57.8000 135.2000 ;
	    RECT 70.2000 134.8000 70.6000 135.2000 ;
	    RECT 49.4000 133.8000 49.8000 134.2000 ;
	    RECT 50.2000 128.2000 50.5000 134.8000 ;
	    RECT 56.6000 134.2000 56.9000 134.8000 ;
	    RECT 57.4000 134.2000 57.7000 134.8000 ;
	    RECT 51.8000 134.1000 52.2000 134.2000 ;
	    RECT 52.6000 134.1000 53.0000 134.2000 ;
	    RECT 51.8000 133.8000 53.0000 134.1000 ;
	    RECT 54.2000 134.1000 54.6000 134.2000 ;
	    RECT 55.0000 134.1000 55.4000 134.2000 ;
	    RECT 54.2000 133.8000 55.4000 134.1000 ;
	    RECT 56.6000 133.8000 57.0000 134.2000 ;
	    RECT 57.4000 133.8000 57.8000 134.2000 ;
	    RECT 67.8000 133.8000 68.2000 134.2000 ;
	    RECT 70.2000 133.8000 70.6000 134.2000 ;
	    RECT 56.6000 133.2000 56.9000 133.8000 ;
	    RECT 56.6000 132.8000 57.0000 133.2000 ;
	    RECT 63.8000 133.1000 64.2000 133.2000 ;
	    RECT 64.6000 133.1000 65.0000 133.2000 ;
	    RECT 63.8000 132.8000 65.0000 133.1000 ;
	    RECT 53.4000 131.8000 53.8000 132.2000 ;
	    RECT 43.8000 127.8000 44.2000 128.2000 ;
	    RECT 50.2000 127.8000 50.6000 128.2000 ;
	    RECT 39.0000 126.8000 39.4000 127.2000 ;
	    RECT 46.2000 126.8000 46.6000 127.2000 ;
	    RECT 52.6000 126.8000 53.0000 127.2000 ;
	    RECT 46.2000 126.2000 46.5000 126.8000 ;
	    RECT 52.6000 126.2000 52.9000 126.8000 ;
	    RECT 39.0000 125.8000 39.4000 126.2000 ;
	    RECT 46.2000 125.8000 46.6000 126.2000 ;
	    RECT 47.8000 126.1000 48.2000 126.2000 ;
	    RECT 48.6000 126.1000 49.0000 126.2000 ;
	    RECT 47.8000 125.8000 49.0000 126.1000 ;
	    RECT 52.6000 125.8000 53.0000 126.2000 ;
	    RECT 39.0000 125.2000 39.3000 125.8000 ;
	    RECT 37.4000 125.1000 37.8000 125.2000 ;
	    RECT 38.2000 125.1000 38.6000 125.2000 ;
	    RECT 37.4000 124.8000 38.6000 125.1000 ;
	    RECT 39.0000 124.8000 39.4000 125.2000 ;
	    RECT 41.4000 124.8000 41.8000 125.2000 ;
	    RECT 43.0000 124.8000 43.4000 125.2000 ;
	    RECT 49.4000 125.1000 49.8000 125.2000 ;
	    RECT 50.2000 125.1000 50.6000 125.2000 ;
	    RECT 49.4000 124.8000 50.6000 125.1000 ;
	    RECT 38.2000 124.1000 38.6000 124.2000 ;
	    RECT 39.0000 124.1000 39.4000 124.2000 ;
	    RECT 38.2000 123.8000 39.4000 124.1000 ;
	    RECT 41.4000 121.2000 41.7000 124.8000 ;
	    RECT 43.0000 124.2000 43.3000 124.8000 ;
	    RECT 43.0000 123.8000 43.4000 124.2000 ;
	    RECT 47.0000 124.1000 47.4000 124.2000 ;
	    RECT 47.8000 124.1000 48.2000 124.2000 ;
	    RECT 47.0000 123.8000 48.2000 124.1000 ;
	    RECT 53.4000 124.1000 53.7000 131.8000 ;
	    RECT 56.6000 129.2000 56.9000 132.8000 ;
	    RECT 59.0000 131.8000 59.4000 132.2000 ;
	    RECT 63.0000 131.8000 63.4000 132.2000 ;
	    RECT 56.6000 128.8000 57.0000 129.2000 ;
	    RECT 54.2000 126.1000 54.6000 126.2000 ;
	    RECT 55.0000 126.1000 55.4000 126.2000 ;
	    RECT 54.2000 125.8000 55.4000 126.1000 ;
	    RECT 55.8000 125.1000 56.2000 125.2000 ;
	    RECT 56.6000 125.1000 57.0000 125.2000 ;
	    RECT 55.8000 124.8000 57.0000 125.1000 ;
	    RECT 59.0000 124.2000 59.3000 131.8000 ;
	    RECT 63.0000 126.2000 63.3000 131.8000 ;
	    RECT 63.8000 128.2000 64.1000 132.8000 ;
	    RECT 63.8000 127.8000 64.2000 128.2000 ;
	    RECT 66.2000 127.8000 66.6000 128.2000 ;
	    RECT 66.2000 127.2000 66.5000 127.8000 ;
	    RECT 66.2000 126.8000 66.6000 127.2000 ;
	    RECT 67.8000 126.2000 68.1000 133.8000 ;
	    RECT 70.2000 133.2000 70.5000 133.8000 ;
	    RECT 72.6000 133.2000 72.9000 142.8000 ;
	    RECT 75.0000 141.8000 75.4000 142.2000 ;
	    RECT 75.0000 136.2000 75.3000 141.8000 ;
	    RECT 76.6000 137.2000 76.9000 148.8000 ;
	    RECT 77.4000 146.2000 77.7000 148.8000 ;
	    RECT 79.0000 148.2000 79.3000 151.8000 ;
	    RECT 79.8000 148.8000 80.2000 149.2000 ;
	    RECT 79.0000 147.8000 79.4000 148.2000 ;
	    RECT 78.2000 147.1000 78.6000 147.2000 ;
	    RECT 79.0000 147.1000 79.4000 147.2000 ;
	    RECT 78.2000 146.8000 79.4000 147.1000 ;
	    RECT 77.4000 145.8000 77.8000 146.2000 ;
	    RECT 79.8000 145.2000 80.1000 148.8000 ;
	    RECT 83.8000 148.2000 84.1000 152.8000 ;
	    RECT 82.2000 147.8000 82.6000 148.2000 ;
	    RECT 83.8000 147.8000 84.2000 148.2000 ;
	    RECT 81.4000 145.8000 81.8000 146.2000 ;
	    RECT 79.8000 144.8000 80.2000 145.2000 ;
	    RECT 78.2000 143.8000 78.6000 144.2000 ;
	    RECT 76.6000 136.8000 77.0000 137.2000 ;
	    RECT 78.2000 136.2000 78.5000 143.8000 ;
	    RECT 81.4000 143.1000 81.7000 145.8000 ;
	    RECT 82.2000 144.2000 82.5000 147.8000 ;
	    RECT 85.4000 147.2000 85.7000 153.8000 ;
	    RECT 87.0000 153.2000 87.3000 154.7000 ;
	    RECT 87.0000 152.8000 87.4000 153.2000 ;
	    RECT 87.8000 152.1000 88.2000 157.9000 ;
	    RECT 90.2000 156.8000 90.6000 157.2000 ;
	    RECT 115.8000 156.8000 116.2000 157.2000 ;
	    RECT 139.8000 157.1000 140.2000 157.2000 ;
	    RECT 140.6000 157.1000 141.0000 157.2000 ;
	    RECT 147.0000 157.1000 147.4000 157.2000 ;
	    RECT 139.8000 156.8000 141.0000 157.1000 ;
	    RECT 146.2000 156.8000 147.4000 157.1000 ;
	    RECT 147.8000 156.8000 148.2000 157.2000 ;
	    RECT 150.2000 157.1000 150.6000 157.2000 ;
	    RECT 151.0000 157.1000 151.4000 157.2000 ;
	    RECT 150.2000 156.8000 151.4000 157.1000 ;
	    RECT 151.8000 156.8000 152.2000 157.2000 ;
	    RECT 159.0000 156.8000 159.4000 157.2000 ;
	    RECT 90.2000 156.2000 90.5000 156.8000 ;
	    RECT 115.8000 156.2000 116.1000 156.8000 ;
	    RECT 88.6000 153.8000 89.0000 154.2000 ;
	    RECT 87.0000 150.8000 87.4000 151.2000 ;
	    RECT 86.2000 147.8000 86.6000 148.2000 ;
	    RECT 86.2000 147.2000 86.5000 147.8000 ;
	    RECT 85.4000 146.8000 85.8000 147.2000 ;
	    RECT 86.2000 146.8000 86.6000 147.2000 ;
	    RECT 83.8000 146.1000 84.2000 146.2000 ;
	    RECT 84.6000 146.1000 85.0000 146.2000 ;
	    RECT 83.8000 145.8000 85.0000 146.1000 ;
	    RECT 82.2000 143.8000 82.6000 144.2000 ;
	    RECT 81.4000 142.8000 82.5000 143.1000 ;
	    RECT 79.0000 141.8000 79.4000 142.2000 ;
	    RECT 79.0000 136.2000 79.3000 141.8000 ;
	    RECT 81.4000 136.8000 81.8000 137.2000 ;
	    RECT 81.4000 136.2000 81.7000 136.8000 ;
	    RECT 75.0000 135.8000 75.4000 136.2000 ;
	    RECT 78.2000 135.8000 78.6000 136.2000 ;
	    RECT 79.0000 135.8000 79.4000 136.2000 ;
	    RECT 81.4000 135.8000 81.8000 136.2000 ;
	    RECT 77.4000 134.8000 77.8000 135.2000 ;
	    RECT 77.4000 134.2000 77.7000 134.8000 ;
	    RECT 75.0000 133.8000 75.4000 134.2000 ;
	    RECT 77.4000 133.8000 77.8000 134.2000 ;
	    RECT 75.0000 133.2000 75.3000 133.8000 ;
	    RECT 70.2000 132.8000 70.6000 133.2000 ;
	    RECT 72.6000 132.8000 73.0000 133.2000 ;
	    RECT 75.0000 132.8000 75.4000 133.2000 ;
	    RECT 68.6000 131.8000 69.0000 132.2000 ;
	    RECT 68.6000 128.2000 68.9000 131.8000 ;
	    RECT 70.2000 128.2000 70.5000 132.8000 ;
	    RECT 71.8000 131.8000 72.2000 132.2000 ;
	    RECT 77.4000 131.8000 77.8000 132.2000 ;
	    RECT 68.6000 127.8000 69.0000 128.2000 ;
	    RECT 70.2000 127.8000 70.6000 128.2000 ;
	    RECT 71.0000 126.8000 71.4000 127.2000 ;
	    RECT 71.0000 126.2000 71.3000 126.8000 ;
	    RECT 62.2000 125.8000 62.6000 126.2000 ;
	    RECT 63.0000 125.8000 63.4000 126.2000 ;
	    RECT 66.2000 125.8000 66.6000 126.2000 ;
	    RECT 67.8000 125.8000 68.2000 126.2000 ;
	    RECT 68.6000 125.8000 69.0000 126.2000 ;
	    RECT 71.0000 125.8000 71.4000 126.2000 ;
	    RECT 54.2000 124.1000 54.6000 124.2000 ;
	    RECT 53.4000 123.8000 54.6000 124.1000 ;
	    RECT 55.0000 123.8000 55.4000 124.2000 ;
	    RECT 59.0000 123.8000 59.4000 124.2000 ;
	    RECT 60.6000 124.1000 61.0000 124.2000 ;
	    RECT 61.4000 124.1000 61.8000 124.2000 ;
	    RECT 60.6000 123.8000 61.8000 124.1000 ;
	    RECT 55.0000 123.2000 55.3000 123.8000 ;
	    RECT 62.2000 123.2000 62.5000 125.8000 ;
	    RECT 55.0000 122.8000 55.4000 123.2000 ;
	    RECT 62.2000 122.8000 62.6000 123.2000 ;
	    RECT 48.6000 121.8000 49.0000 122.2000 ;
	    RECT 62.2000 121.8000 62.6000 122.2000 ;
	    RECT 41.4000 120.8000 41.8000 121.2000 ;
	    RECT 48.6000 117.2000 48.9000 121.8000 ;
	    RECT 52.6000 118.8000 53.0000 119.2000 ;
	    RECT 52.6000 118.2000 52.9000 118.8000 ;
	    RECT 52.6000 117.8000 53.0000 118.2000 ;
	    RECT 57.4000 117.8000 57.8000 118.2000 ;
	    RECT 57.4000 117.2000 57.7000 117.8000 ;
	    RECT 35.8000 116.8000 36.9000 117.1000 ;
	    RECT 37.4000 116.8000 37.8000 117.2000 ;
	    RECT 39.0000 116.8000 39.4000 117.2000 ;
	    RECT 45.4000 117.1000 45.8000 117.2000 ;
	    RECT 46.2000 117.1000 46.6000 117.2000 ;
	    RECT 45.4000 116.8000 46.6000 117.1000 ;
	    RECT 48.6000 116.8000 49.0000 117.2000 ;
	    RECT 57.4000 116.8000 57.8000 117.2000 ;
	    RECT 37.4000 116.2000 37.7000 116.8000 ;
	    RECT 39.0000 116.2000 39.3000 116.8000 ;
	    RECT 37.4000 115.8000 37.8000 116.2000 ;
	    RECT 39.0000 115.8000 39.4000 116.2000 ;
	    RECT 47.8000 116.1000 48.2000 116.2000 ;
	    RECT 48.6000 116.1000 49.0000 116.2000 ;
	    RECT 47.8000 115.8000 49.0000 116.1000 ;
	    RECT 32.6000 114.8000 33.0000 115.2000 ;
	    RECT 35.0000 114.8000 35.4000 115.2000 ;
	    RECT 38.2000 114.8000 38.6000 115.2000 ;
	    RECT 47.0000 114.8000 47.4000 115.2000 ;
	    RECT 56.6000 114.8000 57.0000 115.2000 ;
	    RECT 35.0000 111.8000 35.4000 112.2000 ;
	    RECT 31.8000 108.8000 32.2000 109.2000 ;
	    RECT 31.0000 106.8000 31.4000 107.2000 ;
	    RECT 31.0000 105.8000 31.4000 106.2000 ;
	    RECT 31.0000 105.2000 31.3000 105.8000 ;
	    RECT 31.0000 104.8000 31.4000 105.2000 ;
	    RECT 26.2000 103.8000 26.6000 104.2000 ;
	    RECT 27.8000 103.8000 28.2000 104.2000 ;
	    RECT 29.4000 103.8000 29.8000 104.2000 ;
	    RECT 26.2000 102.2000 26.5000 103.8000 ;
	    RECT 26.2000 101.8000 26.6000 102.2000 ;
	    RECT 26.2000 96.2000 26.5000 101.8000 ;
	    RECT 30.2000 97.8000 30.6000 98.2000 ;
	    RECT 30.2000 97.2000 30.5000 97.8000 ;
	    RECT 35.0000 97.2000 35.3000 111.8000 ;
	    RECT 35.8000 106.1000 36.2000 106.2000 ;
	    RECT 36.6000 106.1000 37.0000 106.2000 ;
	    RECT 35.8000 105.8000 37.0000 106.1000 ;
	    RECT 35.8000 104.8000 36.2000 105.2000 ;
	    RECT 37.4000 104.8000 37.8000 105.2000 ;
	    RECT 35.8000 104.2000 36.1000 104.8000 ;
	    RECT 35.8000 103.8000 36.2000 104.2000 ;
	    RECT 36.6000 101.8000 37.0000 102.2000 ;
	    RECT 36.6000 99.2000 36.9000 101.8000 ;
	    RECT 36.6000 98.8000 37.0000 99.2000 ;
	    RECT 27.8000 97.1000 28.2000 97.2000 ;
	    RECT 28.6000 97.1000 29.0000 97.2000 ;
	    RECT 27.8000 96.8000 29.0000 97.1000 ;
	    RECT 30.2000 96.8000 30.6000 97.2000 ;
	    RECT 31.0000 97.1000 31.4000 97.2000 ;
	    RECT 31.0000 96.8000 32.1000 97.1000 ;
	    RECT 35.0000 96.8000 35.4000 97.2000 ;
	    RECT 35.8000 97.1000 36.2000 97.2000 ;
	    RECT 36.6000 97.1000 37.0000 97.2000 ;
	    RECT 35.8000 96.8000 37.0000 97.1000 ;
	    RECT 25.4000 95.8000 25.8000 96.2000 ;
	    RECT 26.2000 95.8000 26.6000 96.2000 ;
	    RECT 27.0000 95.8000 27.4000 96.2000 ;
	    RECT 7.8000 94.8000 8.2000 95.2000 ;
	    RECT 11.8000 94.8000 12.2000 95.2000 ;
	    RECT 13.4000 94.8000 13.8000 95.2000 ;
	    RECT 15.8000 95.1000 16.2000 95.2000 ;
	    RECT 15.8000 94.8000 16.9000 95.1000 ;
	    RECT 7.8000 94.2000 8.1000 94.8000 ;
	    RECT 11.8000 94.2000 12.1000 94.8000 ;
	    RECT 7.8000 93.8000 8.2000 94.2000 ;
	    RECT 9.4000 93.8000 9.8000 94.2000 ;
	    RECT 11.8000 93.8000 12.2000 94.2000 ;
	    RECT 9.4000 93.2000 9.7000 93.8000 ;
	    RECT 13.4000 93.2000 13.7000 94.8000 ;
	    RECT 16.6000 94.2000 16.9000 94.8000 ;
	    RECT 17.4000 94.8000 17.8000 95.2000 ;
	    RECT 22.2000 94.8000 22.6000 95.2000 ;
	    RECT 24.6000 94.8000 25.0000 95.2000 ;
	    RECT 15.8000 93.8000 16.2000 94.2000 ;
	    RECT 16.6000 93.8000 17.0000 94.2000 ;
	    RECT 15.8000 93.2000 16.1000 93.8000 ;
	    RECT 9.4000 92.8000 9.8000 93.2000 ;
	    RECT 13.4000 92.8000 13.8000 93.2000 ;
	    RECT 15.8000 92.8000 16.2000 93.2000 ;
	    RECT 11.8000 91.8000 12.2000 92.2000 ;
	    RECT 11.8000 89.2000 12.1000 91.8000 ;
	    RECT 6.2000 88.8000 6.6000 89.2000 ;
	    RECT 11.8000 88.8000 12.2000 89.2000 ;
	    RECT 6.2000 88.2000 6.5000 88.8000 ;
	    RECT 17.4000 88.2000 17.7000 94.8000 ;
	    RECT 22.2000 94.2000 22.5000 94.8000 ;
	    RECT 22.2000 93.8000 22.6000 94.2000 ;
	    RECT 25.4000 93.8000 25.8000 94.2000 ;
	    RECT 25.4000 93.2000 25.7000 93.8000 ;
	    RECT 25.4000 92.8000 25.8000 93.2000 ;
	    RECT 23.8000 88.8000 24.2000 89.2000 ;
	    RECT 6.2000 87.8000 6.6000 88.2000 ;
	    RECT 8.6000 87.8000 9.0000 88.2000 ;
	    RECT 17.4000 87.8000 17.8000 88.2000 ;
	    RECT 19.0000 88.1000 19.4000 88.2000 ;
	    RECT 19.8000 88.1000 20.2000 88.2000 ;
	    RECT 19.0000 87.8000 20.2000 88.1000 ;
	    RECT 23.0000 87.8000 23.4000 88.2000 ;
	    RECT 8.6000 87.2000 8.9000 87.8000 ;
	    RECT 17.4000 87.2000 17.7000 87.8000 ;
	    RECT 8.6000 86.8000 9.0000 87.2000 ;
	    RECT 11.0000 86.8000 11.4000 87.2000 ;
	    RECT 17.4000 86.8000 17.8000 87.2000 ;
	    RECT 19.0000 87.1000 19.4000 87.2000 ;
	    RECT 19.8000 87.1000 20.2000 87.2000 ;
	    RECT 19.0000 86.8000 20.2000 87.1000 ;
	    RECT 22.2000 86.8000 22.6000 87.2000 ;
	    RECT 11.0000 86.2000 11.3000 86.8000 ;
	    RECT 22.2000 86.2000 22.5000 86.8000 ;
	    RECT 11.0000 85.8000 11.4000 86.2000 ;
	    RECT 13.4000 86.1000 13.8000 86.2000 ;
	    RECT 14.2000 86.1000 14.6000 86.2000 ;
	    RECT 13.4000 85.8000 14.6000 86.1000 ;
	    RECT 17.4000 85.8000 17.8000 86.2000 ;
	    RECT 22.2000 85.8000 22.6000 86.2000 ;
	    RECT 17.4000 85.2000 17.7000 85.8000 ;
	    RECT 23.0000 85.2000 23.3000 87.8000 ;
	    RECT 23.8000 86.2000 24.1000 88.8000 ;
	    RECT 26.2000 88.2000 26.5000 95.8000 ;
	    RECT 27.0000 95.2000 27.3000 95.8000 ;
	    RECT 27.0000 94.8000 27.4000 95.2000 ;
	    RECT 28.6000 94.8000 29.0000 95.2000 ;
	    RECT 30.2000 95.1000 30.6000 95.2000 ;
	    RECT 31.0000 95.1000 31.4000 95.2000 ;
	    RECT 30.2000 94.8000 31.4000 95.1000 ;
	    RECT 28.6000 94.2000 28.9000 94.8000 ;
	    RECT 28.6000 93.8000 29.0000 94.2000 ;
	    RECT 31.8000 94.1000 32.1000 96.8000 ;
	    RECT 32.6000 95.8000 33.0000 96.2000 ;
	    RECT 37.4000 96.1000 37.7000 104.8000 ;
	    RECT 38.2000 104.1000 38.5000 114.8000 ;
	    RECT 47.0000 114.2000 47.3000 114.8000 ;
	    RECT 56.6000 114.2000 56.9000 114.8000 ;
	    RECT 39.0000 113.8000 39.4000 114.2000 ;
	    RECT 44.6000 113.8000 45.0000 114.2000 ;
	    RECT 47.0000 113.8000 47.4000 114.2000 ;
	    RECT 51.0000 113.8000 51.4000 114.2000 ;
	    RECT 51.8000 113.8000 52.2000 114.2000 ;
	    RECT 56.6000 113.8000 57.0000 114.2000 ;
	    RECT 39.0000 112.2000 39.3000 113.8000 ;
	    RECT 44.6000 113.2000 44.9000 113.8000 ;
	    RECT 51.0000 113.2000 51.3000 113.8000 ;
	    RECT 51.8000 113.2000 52.1000 113.8000 ;
	    RECT 42.2000 112.8000 42.6000 113.2000 ;
	    RECT 44.6000 112.8000 45.0000 113.2000 ;
	    RECT 48.6000 112.8000 49.0000 113.2000 ;
	    RECT 51.0000 112.8000 51.4000 113.2000 ;
	    RECT 51.8000 112.8000 52.2000 113.2000 ;
	    RECT 59.0000 112.8000 59.4000 113.2000 ;
	    RECT 39.0000 111.8000 39.4000 112.2000 ;
	    RECT 41.4000 111.8000 41.8000 112.2000 ;
	    RECT 41.4000 108.2000 41.7000 111.8000 ;
	    RECT 41.4000 107.8000 41.8000 108.2000 ;
	    RECT 39.0000 106.1000 39.4000 106.2000 ;
	    RECT 39.8000 106.1000 40.2000 106.2000 ;
	    RECT 39.0000 105.8000 40.2000 106.1000 ;
	    RECT 39.8000 105.1000 40.2000 105.2000 ;
	    RECT 40.6000 105.1000 41.0000 105.2000 ;
	    RECT 39.8000 104.8000 41.0000 105.1000 ;
	    RECT 39.0000 104.1000 39.4000 104.2000 ;
	    RECT 38.2000 103.8000 39.4000 104.1000 ;
	    RECT 39.8000 101.8000 40.2000 102.2000 ;
	    RECT 39.8000 101.2000 40.1000 101.8000 ;
	    RECT 39.8000 100.8000 40.2000 101.2000 ;
	    RECT 42.2000 98.1000 42.5000 112.8000 ;
	    RECT 48.6000 112.2000 48.9000 112.8000 ;
	    RECT 51.8000 112.2000 52.1000 112.8000 ;
	    RECT 59.0000 112.2000 59.3000 112.8000 ;
	    RECT 47.0000 111.8000 47.4000 112.2000 ;
	    RECT 48.6000 112.1000 49.0000 112.2000 ;
	    RECT 47.8000 111.8000 49.0000 112.1000 ;
	    RECT 51.8000 111.8000 52.2000 112.2000 ;
	    RECT 57.4000 111.8000 57.8000 112.2000 ;
	    RECT 59.0000 111.8000 59.4000 112.2000 ;
	    RECT 47.0000 110.2000 47.3000 111.8000 ;
	    RECT 47.0000 109.8000 47.4000 110.2000 ;
	    RECT 47.8000 107.2000 48.1000 111.8000 ;
	    RECT 51.8000 108.2000 52.1000 111.8000 ;
	    RECT 51.8000 107.8000 52.2000 108.2000 ;
	    RECT 57.4000 107.2000 57.7000 111.8000 ;
	    RECT 43.8000 106.8000 44.2000 107.2000 ;
	    RECT 47.8000 106.8000 48.2000 107.2000 ;
	    RECT 54.2000 106.8000 54.6000 107.2000 ;
	    RECT 57.4000 106.8000 57.8000 107.2000 ;
	    RECT 58.2000 107.1000 58.6000 107.2000 ;
	    RECT 59.0000 107.1000 59.3000 111.8000 ;
	    RECT 62.2000 108.2000 62.5000 121.8000 ;
	    RECT 66.2000 117.2000 66.5000 125.8000 ;
	    RECT 67.0000 125.1000 67.4000 125.2000 ;
	    RECT 67.8000 125.1000 68.2000 125.2000 ;
	    RECT 67.0000 124.8000 68.2000 125.1000 ;
	    RECT 68.6000 124.2000 68.9000 125.8000 ;
	    RECT 71.0000 124.8000 71.4000 125.2000 ;
	    RECT 71.0000 124.2000 71.3000 124.8000 ;
	    RECT 71.8000 124.2000 72.1000 131.8000 ;
	    RECT 73.4000 127.8000 73.8000 128.2000 ;
	    RECT 73.4000 127.2000 73.7000 127.8000 ;
	    RECT 73.4000 126.8000 73.8000 127.2000 ;
	    RECT 73.4000 125.8000 73.8000 126.2000 ;
	    RECT 77.4000 126.1000 77.7000 131.8000 ;
	    RECT 78.2000 131.2000 78.5000 135.8000 ;
	    RECT 82.2000 134.1000 82.5000 142.8000 ;
	    RECT 83.0000 141.8000 83.4000 142.2000 ;
	    RECT 83.0000 135.2000 83.3000 141.8000 ;
	    RECT 85.4000 136.2000 85.7000 146.8000 ;
	    RECT 87.0000 146.2000 87.3000 150.8000 ;
	    RECT 87.8000 149.8000 88.2000 150.2000 ;
	    RECT 87.8000 147.2000 88.1000 149.8000 ;
	    RECT 87.8000 146.8000 88.2000 147.2000 ;
	    RECT 86.2000 146.1000 86.6000 146.2000 ;
	    RECT 87.0000 146.1000 87.4000 146.2000 ;
	    RECT 86.2000 145.8000 87.4000 146.1000 ;
	    RECT 88.6000 141.2000 88.9000 153.8000 ;
	    RECT 89.4000 153.1000 89.8000 155.9000 ;
	    RECT 90.2000 155.8000 90.6000 156.2000 ;
	    RECT 97.4000 156.1000 97.8000 156.2000 ;
	    RECT 98.2000 156.1000 98.6000 156.2000 ;
	    RECT 97.4000 155.8000 98.6000 156.1000 ;
	    RECT 99.8000 155.8000 100.2000 156.2000 ;
	    RECT 100.6000 155.8000 101.0000 156.2000 ;
	    RECT 107.0000 156.1000 107.4000 156.2000 ;
	    RECT 107.8000 156.1000 108.2000 156.2000 ;
	    RECT 107.0000 155.8000 108.2000 156.1000 ;
	    RECT 109.4000 155.8000 109.8000 156.2000 ;
	    RECT 115.8000 155.8000 116.2000 156.2000 ;
	    RECT 116.6000 156.1000 117.0000 156.2000 ;
	    RECT 117.4000 156.1000 117.8000 156.2000 ;
	    RECT 116.6000 155.8000 117.8000 156.1000 ;
	    RECT 129.4000 156.1000 129.8000 156.2000 ;
	    RECT 130.2000 156.1000 130.6000 156.2000 ;
	    RECT 129.4000 155.8000 130.6000 156.1000 ;
	    RECT 136.6000 155.8000 137.0000 156.2000 ;
	    RECT 143.0000 155.8000 143.4000 156.2000 ;
	    RECT 145.4000 155.8000 145.8000 156.2000 ;
	    RECT 99.8000 155.2000 100.1000 155.8000 ;
	    RECT 92.6000 155.1000 93.0000 155.2000 ;
	    RECT 93.4000 155.1000 93.8000 155.2000 ;
	    RECT 92.6000 154.8000 93.8000 155.1000 ;
	    RECT 94.2000 154.8000 94.6000 155.2000 ;
	    RECT 96.6000 154.8000 97.0000 155.2000 ;
	    RECT 98.2000 154.8000 98.6000 155.2000 ;
	    RECT 99.8000 154.8000 100.2000 155.2000 ;
	    RECT 94.2000 154.2000 94.5000 154.8000 ;
	    RECT 96.6000 154.2000 96.9000 154.8000 ;
	    RECT 91.0000 153.8000 91.4000 154.2000 ;
	    RECT 94.2000 153.8000 94.6000 154.2000 ;
	    RECT 95.0000 153.8000 95.4000 154.2000 ;
	    RECT 95.8000 153.8000 96.2000 154.2000 ;
	    RECT 96.6000 153.8000 97.0000 154.2000 ;
	    RECT 91.0000 153.2000 91.3000 153.8000 ;
	    RECT 91.0000 152.8000 91.4000 153.2000 ;
	    RECT 91.0000 150.2000 91.3000 152.8000 ;
	    RECT 93.4000 152.1000 93.8000 152.2000 ;
	    RECT 94.2000 152.1000 94.6000 152.2000 ;
	    RECT 93.4000 151.8000 94.6000 152.1000 ;
	    RECT 91.0000 149.8000 91.4000 150.2000 ;
	    RECT 91.0000 148.8000 91.4000 149.2000 ;
	    RECT 91.0000 148.2000 91.3000 148.8000 ;
	    RECT 95.0000 148.2000 95.3000 153.8000 ;
	    RECT 95.8000 151.2000 96.1000 153.8000 ;
	    RECT 98.2000 152.2000 98.5000 154.8000 ;
	    RECT 99.8000 153.8000 100.2000 154.2000 ;
	    RECT 99.8000 153.2000 100.1000 153.8000 ;
	    RECT 99.8000 152.8000 100.2000 153.2000 ;
	    RECT 100.6000 152.2000 100.9000 155.8000 ;
	    RECT 109.4000 155.2000 109.7000 155.8000 ;
	    RECT 109.4000 154.8000 109.8000 155.2000 ;
	    RECT 115.8000 155.1000 116.2000 155.2000 ;
	    RECT 116.6000 155.1000 117.0000 155.2000 ;
	    RECT 115.8000 154.8000 117.0000 155.1000 ;
	    RECT 117.4000 154.2000 117.7000 155.8000 ;
	    RECT 118.2000 154.8000 118.6000 155.2000 ;
	    RECT 122.2000 154.8000 122.6000 155.2000 ;
	    RECT 123.8000 155.1000 124.2000 155.2000 ;
	    RECT 124.6000 155.1000 125.0000 155.2000 ;
	    RECT 123.8000 154.8000 125.0000 155.1000 ;
	    RECT 129.4000 155.1000 129.8000 155.2000 ;
	    RECT 130.2000 155.1000 130.6000 155.2000 ;
	    RECT 129.4000 154.8000 130.6000 155.1000 ;
	    RECT 131.0000 155.1000 131.4000 155.2000 ;
	    RECT 131.8000 155.1000 132.2000 155.2000 ;
	    RECT 131.0000 154.8000 132.2000 155.1000 ;
	    RECT 132.6000 154.8000 133.0000 155.2000 ;
	    RECT 118.2000 154.2000 118.5000 154.8000 ;
	    RECT 106.2000 153.8000 106.6000 154.2000 ;
	    RECT 109.4000 153.8000 109.8000 154.2000 ;
	    RECT 111.8000 153.8000 112.2000 154.2000 ;
	    RECT 113.4000 154.1000 113.8000 154.2000 ;
	    RECT 114.2000 154.1000 114.6000 154.2000 ;
	    RECT 113.4000 153.8000 114.6000 154.1000 ;
	    RECT 115.0000 154.1000 115.4000 154.2000 ;
	    RECT 115.8000 154.1000 116.2000 154.2000 ;
	    RECT 115.0000 153.8000 116.2000 154.1000 ;
	    RECT 117.4000 153.8000 117.8000 154.2000 ;
	    RECT 118.2000 153.8000 118.6000 154.2000 ;
	    RECT 121.4000 153.8000 121.8000 154.2000 ;
	    RECT 101.4000 152.8000 101.8000 153.2000 ;
	    RECT 104.6000 152.8000 105.0000 153.2000 ;
	    RECT 98.2000 151.8000 98.6000 152.2000 ;
	    RECT 100.6000 151.8000 101.0000 152.2000 ;
	    RECT 95.8000 150.8000 96.2000 151.2000 ;
	    RECT 99.0000 150.8000 99.4000 151.2000 ;
	    RECT 99.0000 149.2000 99.3000 150.8000 ;
	    RECT 99.0000 148.8000 99.4000 149.2000 ;
	    RECT 89.4000 147.8000 89.8000 148.2000 ;
	    RECT 91.0000 147.8000 91.4000 148.2000 ;
	    RECT 95.0000 147.8000 95.4000 148.2000 ;
	    RECT 95.8000 147.8000 96.2000 148.2000 ;
	    RECT 96.6000 147.8000 97.0000 148.2000 ;
	    RECT 99.8000 147.8000 100.2000 148.2000 ;
	    RECT 89.4000 147.2000 89.7000 147.8000 ;
	    RECT 95.8000 147.2000 96.1000 147.8000 ;
	    RECT 89.4000 146.8000 89.8000 147.2000 ;
	    RECT 90.2000 146.8000 90.6000 147.2000 ;
	    RECT 91.8000 147.1000 92.2000 147.2000 ;
	    RECT 92.6000 147.1000 93.0000 147.2000 ;
	    RECT 91.8000 146.8000 93.0000 147.1000 ;
	    RECT 95.8000 146.8000 96.2000 147.2000 ;
	    RECT 89.4000 145.2000 89.7000 146.8000 ;
	    RECT 90.2000 146.2000 90.5000 146.8000 ;
	    RECT 90.2000 145.8000 90.6000 146.2000 ;
	    RECT 92.6000 145.8000 93.0000 146.2000 ;
	    RECT 93.4000 146.1000 93.8000 146.2000 ;
	    RECT 94.2000 146.1000 94.6000 146.2000 ;
	    RECT 93.4000 145.8000 94.6000 146.1000 ;
	    RECT 95.0000 145.8000 95.4000 146.2000 ;
	    RECT 89.4000 144.8000 89.8000 145.2000 ;
	    RECT 89.4000 141.8000 89.8000 142.2000 ;
	    RECT 91.0000 141.8000 91.4000 142.2000 ;
	    RECT 88.6000 140.8000 89.0000 141.2000 ;
	    RECT 89.4000 136.2000 89.7000 141.8000 ;
	    RECT 91.0000 139.2000 91.3000 141.8000 ;
	    RECT 91.0000 138.8000 91.4000 139.2000 ;
	    RECT 92.6000 137.2000 92.9000 145.8000 ;
	    RECT 95.0000 145.2000 95.3000 145.8000 ;
	    RECT 94.2000 145.1000 94.6000 145.2000 ;
	    RECT 95.0000 145.1000 95.4000 145.2000 ;
	    RECT 94.2000 144.8000 95.4000 145.1000 ;
	    RECT 93.4000 143.8000 93.8000 144.2000 ;
	    RECT 94.2000 143.8000 94.6000 144.2000 ;
	    RECT 93.4000 137.2000 93.7000 143.8000 ;
	    RECT 94.2000 143.2000 94.5000 143.8000 ;
	    RECT 94.2000 142.8000 94.6000 143.2000 ;
	    RECT 95.8000 137.8000 96.2000 138.2000 ;
	    RECT 92.6000 136.8000 93.0000 137.2000 ;
	    RECT 93.4000 137.1000 93.8000 137.2000 ;
	    RECT 94.2000 137.1000 94.6000 137.2000 ;
	    RECT 93.4000 136.8000 94.6000 137.1000 ;
	    RECT 85.4000 135.8000 85.8000 136.2000 ;
	    RECT 89.4000 135.8000 89.8000 136.2000 ;
	    RECT 91.8000 135.8000 92.2000 136.2000 ;
	    RECT 83.0000 134.8000 83.4000 135.2000 ;
	    RECT 83.8000 134.8000 84.2000 135.2000 ;
	    RECT 83.8000 134.2000 84.1000 134.8000 ;
	    RECT 82.2000 133.8000 83.3000 134.1000 ;
	    RECT 83.8000 133.8000 84.2000 134.2000 ;
	    RECT 84.6000 133.8000 85.0000 134.2000 ;
	    RECT 81.4000 132.8000 81.8000 133.2000 ;
	    RECT 81.4000 132.2000 81.7000 132.8000 ;
	    RECT 79.0000 131.8000 79.4000 132.2000 ;
	    RECT 81.4000 131.8000 81.8000 132.2000 ;
	    RECT 78.2000 130.8000 78.6000 131.2000 ;
	    RECT 78.2000 126.1000 78.6000 126.2000 ;
	    RECT 77.4000 125.8000 78.6000 126.1000 ;
	    RECT 73.4000 125.2000 73.7000 125.8000 ;
	    RECT 72.6000 124.8000 73.0000 125.2000 ;
	    RECT 73.4000 124.8000 73.8000 125.2000 ;
	    RECT 68.6000 123.8000 69.0000 124.2000 ;
	    RECT 71.0000 123.8000 71.4000 124.2000 ;
	    RECT 71.8000 123.8000 72.2000 124.2000 ;
	    RECT 71.8000 122.8000 72.2000 123.2000 ;
	    RECT 67.8000 121.8000 68.2000 122.2000 ;
	    RECT 71.0000 121.8000 71.4000 122.2000 ;
	    RECT 66.2000 116.8000 66.6000 117.2000 ;
	    RECT 67.8000 117.1000 68.1000 121.8000 ;
	    RECT 67.0000 116.8000 68.1000 117.1000 ;
	    RECT 69.4000 117.8000 69.8000 118.2000 ;
	    RECT 69.4000 117.2000 69.7000 117.8000 ;
	    RECT 69.4000 116.8000 69.8000 117.2000 ;
	    RECT 71.0000 117.1000 71.3000 121.8000 ;
	    RECT 71.8000 119.2000 72.1000 122.8000 ;
	    RECT 71.8000 118.8000 72.2000 119.2000 ;
	    RECT 70.2000 116.8000 71.3000 117.1000 ;
	    RECT 67.0000 115.2000 67.3000 116.8000 ;
	    RECT 70.2000 115.2000 70.5000 116.8000 ;
	    RECT 67.0000 114.8000 67.4000 115.2000 ;
	    RECT 70.2000 114.8000 70.6000 115.2000 ;
	    RECT 64.6000 111.8000 65.0000 112.2000 ;
	    RECT 67.0000 111.8000 67.4000 112.2000 ;
	    RECT 70.2000 111.8000 70.6000 112.2000 ;
	    RECT 64.6000 110.2000 64.9000 111.8000 ;
	    RECT 67.0000 111.2000 67.3000 111.8000 ;
	    RECT 67.0000 110.8000 67.4000 111.2000 ;
	    RECT 64.6000 109.8000 65.0000 110.2000 ;
	    RECT 70.2000 109.2000 70.5000 111.8000 ;
	    RECT 72.6000 109.2000 72.9000 124.8000 ;
	    RECT 79.0000 124.2000 79.3000 131.8000 ;
	    RECT 81.4000 130.8000 81.8000 131.2000 ;
	    RECT 81.4000 129.2000 81.7000 130.8000 ;
	    RECT 83.0000 129.2000 83.3000 133.8000 ;
	    RECT 84.6000 133.2000 84.9000 133.8000 ;
	    RECT 84.6000 132.8000 85.0000 133.2000 ;
	    RECT 81.4000 128.8000 81.8000 129.2000 ;
	    RECT 83.0000 128.8000 83.4000 129.2000 ;
	    RECT 84.6000 127.2000 84.9000 132.8000 ;
	    RECT 85.4000 129.2000 85.7000 135.8000 ;
	    RECT 86.2000 134.8000 86.6000 135.2000 ;
	    RECT 87.8000 134.8000 88.2000 135.2000 ;
	    RECT 88.6000 135.1000 89.0000 135.2000 ;
	    RECT 89.4000 135.1000 89.8000 135.2000 ;
	    RECT 88.6000 134.8000 89.8000 135.1000 ;
	    RECT 90.2000 134.8000 90.6000 135.2000 ;
	    RECT 85.4000 128.8000 85.8000 129.2000 ;
	    RECT 84.6000 126.8000 85.0000 127.2000 ;
	    RECT 86.2000 125.2000 86.5000 134.8000 ;
	    RECT 87.8000 133.2000 88.1000 134.8000 ;
	    RECT 90.2000 134.2000 90.5000 134.8000 ;
	    RECT 91.8000 134.2000 92.1000 135.8000 ;
	    RECT 92.6000 135.2000 92.9000 136.8000 ;
	    RECT 94.2000 136.1000 94.6000 136.2000 ;
	    RECT 95.0000 136.1000 95.4000 136.2000 ;
	    RECT 94.2000 135.8000 95.4000 136.1000 ;
	    RECT 95.8000 135.2000 96.1000 137.8000 ;
	    RECT 96.6000 137.2000 96.9000 147.8000 ;
	    RECT 99.8000 147.2000 100.1000 147.8000 ;
	    RECT 98.2000 147.1000 98.6000 147.2000 ;
	    RECT 98.2000 146.8000 99.3000 147.1000 ;
	    RECT 99.0000 146.2000 99.3000 146.8000 ;
	    RECT 99.8000 146.8000 100.2000 147.2000 ;
	    RECT 97.4000 146.1000 97.8000 146.2000 ;
	    RECT 98.2000 146.1000 98.6000 146.2000 ;
	    RECT 97.4000 145.8000 98.6000 146.1000 ;
	    RECT 99.0000 145.8000 99.4000 146.2000 ;
	    RECT 97.4000 145.1000 97.8000 145.2000 ;
	    RECT 97.4000 144.8000 98.5000 145.1000 ;
	    RECT 96.6000 136.8000 97.0000 137.2000 ;
	    RECT 97.4000 135.8000 97.8000 136.2000 ;
	    RECT 97.4000 135.2000 97.7000 135.8000 ;
	    RECT 92.6000 134.8000 93.0000 135.2000 ;
	    RECT 94.2000 134.8000 94.6000 135.2000 ;
	    RECT 95.8000 134.8000 96.2000 135.2000 ;
	    RECT 97.4000 134.8000 97.8000 135.2000 ;
	    RECT 94.2000 134.2000 94.5000 134.8000 ;
	    RECT 90.2000 133.8000 90.6000 134.2000 ;
	    RECT 91.8000 133.8000 92.2000 134.2000 ;
	    RECT 94.2000 133.8000 94.6000 134.2000 ;
	    RECT 97.4000 133.8000 97.8000 134.2000 ;
	    RECT 87.8000 132.8000 88.2000 133.2000 ;
	    RECT 83.0000 125.1000 83.4000 125.2000 ;
	    RECT 83.8000 125.1000 84.2000 125.2000 ;
	    RECT 83.0000 124.8000 84.2000 125.1000 ;
	    RECT 86.2000 124.8000 86.6000 125.2000 ;
	    RECT 79.0000 123.8000 79.4000 124.2000 ;
	    RECT 87.8000 123.1000 88.2000 128.9000 ;
	    RECT 88.6000 125.8000 89.0000 126.2000 ;
	    RECT 79.8000 121.8000 80.2000 122.2000 ;
	    RECT 74.2000 112.1000 74.6000 117.9000 ;
	    RECT 78.2000 114.7000 78.6000 115.1000 ;
	    RECT 78.2000 114.2000 78.5000 114.7000 ;
	    RECT 78.2000 113.8000 78.6000 114.2000 ;
	    RECT 79.0000 112.1000 79.4000 117.9000 ;
	    RECT 79.8000 112.2000 80.1000 121.8000 ;
	    RECT 80.6000 113.1000 81.0000 115.9000 ;
	    RECT 81.4000 113.1000 81.8000 115.9000 ;
	    RECT 79.8000 111.8000 80.2000 112.2000 ;
	    RECT 83.0000 112.1000 83.4000 117.9000 ;
	    RECT 87.0000 115.8000 87.4000 116.2000 ;
	    RECT 87.0000 115.2000 87.3000 115.8000 ;
	    RECT 83.8000 114.7000 84.2000 115.1000 ;
	    RECT 87.0000 114.8000 87.4000 115.2000 ;
	    RECT 83.8000 114.2000 84.1000 114.7000 ;
	    RECT 83.8000 113.8000 84.2000 114.2000 ;
	    RECT 87.8000 112.1000 88.2000 117.9000 ;
	    RECT 88.6000 117.2000 88.9000 125.8000 ;
	    RECT 90.2000 119.2000 90.5000 133.8000 ;
	    RECT 97.4000 129.2000 97.7000 133.8000 ;
	    RECT 98.2000 132.2000 98.5000 144.8000 ;
	    RECT 99.8000 140.2000 100.1000 146.8000 ;
	    RECT 100.6000 142.2000 100.9000 151.8000 ;
	    RECT 101.4000 151.2000 101.7000 152.8000 ;
	    RECT 104.6000 152.2000 104.9000 152.8000 ;
	    RECT 106.2000 152.2000 106.5000 153.8000 ;
	    RECT 109.4000 153.2000 109.7000 153.8000 ;
	    RECT 111.8000 153.2000 112.1000 153.8000 ;
	    RECT 109.4000 152.8000 109.8000 153.2000 ;
	    RECT 111.8000 152.8000 112.2000 153.2000 ;
	    RECT 113.4000 152.8000 113.8000 153.2000 ;
	    RECT 103.0000 151.8000 103.4000 152.2000 ;
	    RECT 104.6000 151.8000 105.0000 152.2000 ;
	    RECT 106.2000 151.8000 106.6000 152.2000 ;
	    RECT 101.4000 150.8000 101.8000 151.2000 ;
	    RECT 102.2000 148.8000 102.6000 149.2000 ;
	    RECT 102.2000 148.2000 102.5000 148.8000 ;
	    RECT 103.0000 148.2000 103.3000 151.8000 ;
	    RECT 102.2000 147.8000 102.6000 148.2000 ;
	    RECT 103.0000 147.8000 103.4000 148.2000 ;
	    RECT 110.2000 147.8000 110.6000 148.2000 ;
	    RECT 110.2000 147.2000 110.5000 147.8000 ;
	    RECT 103.8000 146.8000 104.2000 147.2000 ;
	    RECT 108.6000 147.1000 109.0000 147.2000 ;
	    RECT 109.4000 147.1000 109.8000 147.2000 ;
	    RECT 108.6000 146.8000 109.8000 147.1000 ;
	    RECT 110.2000 146.8000 110.6000 147.2000 ;
	    RECT 111.8000 147.1000 112.2000 147.2000 ;
	    RECT 112.6000 147.1000 113.0000 147.2000 ;
	    RECT 111.8000 146.8000 113.0000 147.1000 ;
	    RECT 101.4000 146.1000 101.8000 146.2000 ;
	    RECT 102.2000 146.1000 102.6000 146.2000 ;
	    RECT 101.4000 145.8000 102.6000 146.1000 ;
	    RECT 103.0000 145.1000 103.4000 145.2000 ;
	    RECT 103.8000 145.1000 104.1000 146.8000 ;
	    RECT 113.4000 146.2000 113.7000 152.8000 ;
	    RECT 114.2000 147.2000 114.5000 153.8000 ;
	    RECT 120.6000 151.8000 121.0000 152.2000 ;
	    RECT 117.4000 149.8000 117.8000 150.2000 ;
	    RECT 119.8000 149.8000 120.2000 150.2000 ;
	    RECT 116.6000 147.8000 117.0000 148.2000 ;
	    RECT 114.2000 146.8000 114.6000 147.2000 ;
	    RECT 115.8000 146.8000 116.2000 147.2000 ;
	    RECT 115.8000 146.2000 116.1000 146.8000 ;
	    RECT 105.4000 146.1000 105.8000 146.2000 ;
	    RECT 106.2000 146.1000 106.6000 146.2000 ;
	    RECT 105.4000 145.8000 106.6000 146.1000 ;
	    RECT 107.0000 146.1000 107.4000 146.2000 ;
	    RECT 107.8000 146.1000 108.2000 146.2000 ;
	    RECT 107.0000 145.8000 108.2000 146.1000 ;
	    RECT 111.0000 145.8000 111.4000 146.2000 ;
	    RECT 113.4000 145.8000 113.8000 146.2000 ;
	    RECT 115.0000 145.8000 115.4000 146.2000 ;
	    RECT 115.8000 145.8000 116.2000 146.2000 ;
	    RECT 103.0000 144.8000 104.1000 145.1000 ;
	    RECT 106.2000 145.1000 106.6000 145.2000 ;
	    RECT 107.0000 145.1000 107.4000 145.2000 ;
	    RECT 106.2000 144.8000 107.4000 145.1000 ;
	    RECT 109.4000 144.8000 109.8000 145.2000 ;
	    RECT 101.4000 143.8000 101.8000 144.2000 ;
	    RECT 101.4000 143.2000 101.7000 143.8000 ;
	    RECT 101.4000 142.8000 101.8000 143.2000 ;
	    RECT 100.6000 141.8000 101.0000 142.2000 ;
	    RECT 103.0000 141.8000 103.4000 142.2000 ;
	    RECT 99.8000 139.8000 100.2000 140.2000 ;
	    RECT 99.0000 139.1000 99.4000 139.2000 ;
	    RECT 99.8000 139.1000 100.2000 139.2000 ;
	    RECT 99.0000 138.8000 100.2000 139.1000 ;
	    RECT 99.8000 137.8000 100.2000 138.2000 ;
	    RECT 99.0000 136.8000 99.4000 137.2000 ;
	    RECT 99.0000 136.2000 99.3000 136.8000 ;
	    RECT 99.0000 135.8000 99.4000 136.2000 ;
	    RECT 99.8000 135.2000 100.1000 137.8000 ;
	    RECT 100.6000 136.2000 100.9000 141.8000 ;
	    RECT 101.4000 139.8000 101.8000 140.2000 ;
	    RECT 100.6000 135.8000 101.0000 136.2000 ;
	    RECT 99.8000 134.8000 100.2000 135.2000 ;
	    RECT 99.0000 132.8000 99.4000 133.2000 ;
	    RECT 98.2000 131.8000 98.6000 132.2000 ;
	    RECT 91.0000 126.2000 91.4000 126.3000 ;
	    RECT 91.8000 126.2000 92.2000 126.3000 ;
	    RECT 91.0000 125.9000 92.2000 126.2000 ;
	    RECT 92.6000 123.1000 93.0000 128.9000 ;
	    RECT 97.4000 128.8000 97.8000 129.2000 ;
	    RECT 95.0000 128.1000 95.4000 128.2000 ;
	    RECT 95.8000 128.1000 96.2000 128.2000 ;
	    RECT 94.2000 125.1000 94.6000 127.9000 ;
	    RECT 95.0000 127.8000 96.2000 128.1000 ;
	    RECT 95.0000 119.2000 95.3000 127.8000 ;
	    RECT 98.2000 125.2000 98.5000 131.8000 ;
	    RECT 99.0000 129.2000 99.3000 132.8000 ;
	    RECT 101.4000 129.2000 101.7000 139.8000 ;
	    RECT 103.0000 139.2000 103.3000 141.8000 ;
	    RECT 102.2000 138.8000 102.6000 139.2000 ;
	    RECT 103.0000 138.8000 103.4000 139.2000 ;
	    RECT 102.2000 137.2000 102.5000 138.8000 ;
	    RECT 102.2000 136.8000 102.6000 137.2000 ;
	    RECT 103.8000 136.2000 104.1000 144.8000 ;
	    RECT 109.4000 144.2000 109.7000 144.8000 ;
	    RECT 107.8000 143.8000 108.2000 144.2000 ;
	    RECT 109.4000 143.8000 109.8000 144.2000 ;
	    RECT 107.8000 143.2000 108.1000 143.8000 ;
	    RECT 106.2000 142.8000 106.6000 143.2000 ;
	    RECT 107.8000 143.1000 108.2000 143.2000 ;
	    RECT 107.0000 142.8000 108.2000 143.1000 ;
	    RECT 105.4000 140.8000 105.8000 141.2000 ;
	    RECT 103.8000 135.8000 104.2000 136.2000 ;
	    RECT 102.2000 134.8000 102.6000 135.2000 ;
	    RECT 102.2000 134.2000 102.5000 134.8000 ;
	    RECT 102.2000 133.8000 102.6000 134.2000 ;
	    RECT 103.0000 133.8000 103.4000 134.2000 ;
	    RECT 103.0000 129.2000 103.3000 133.8000 ;
	    RECT 103.8000 130.2000 104.1000 135.8000 ;
	    RECT 104.6000 132.8000 105.0000 133.2000 ;
	    RECT 103.8000 129.8000 104.2000 130.2000 ;
	    RECT 99.0000 128.8000 99.4000 129.2000 ;
	    RECT 101.4000 128.8000 101.8000 129.2000 ;
	    RECT 103.0000 128.8000 103.4000 129.2000 ;
	    RECT 103.8000 128.8000 104.2000 129.2000 ;
	    RECT 100.6000 127.8000 101.0000 128.2000 ;
	    RECT 100.6000 127.2000 100.9000 127.8000 ;
	    RECT 101.4000 127.2000 101.7000 128.8000 ;
	    RECT 103.8000 128.2000 104.1000 128.8000 ;
	    RECT 103.8000 127.8000 104.2000 128.2000 ;
	    RECT 104.6000 127.2000 104.9000 132.8000 ;
	    RECT 100.6000 126.8000 101.0000 127.2000 ;
	    RECT 101.4000 126.8000 101.8000 127.2000 ;
	    RECT 104.6000 126.8000 105.0000 127.2000 ;
	    RECT 99.0000 125.8000 99.4000 126.2000 ;
	    RECT 99.0000 125.2000 99.3000 125.8000 ;
	    RECT 95.8000 125.1000 96.2000 125.2000 ;
	    RECT 96.6000 125.1000 97.0000 125.2000 ;
	    RECT 95.8000 124.8000 97.0000 125.1000 ;
	    RECT 98.2000 124.8000 98.6000 125.2000 ;
	    RECT 99.0000 124.8000 99.4000 125.2000 ;
	    RECT 102.2000 125.1000 102.6000 125.2000 ;
	    RECT 103.0000 125.1000 103.4000 125.2000 ;
	    RECT 102.2000 124.8000 103.4000 125.1000 ;
	    RECT 104.6000 123.2000 104.9000 126.8000 ;
	    RECT 105.4000 124.2000 105.7000 140.8000 ;
	    RECT 106.2000 139.2000 106.5000 142.8000 ;
	    RECT 106.2000 138.8000 106.6000 139.2000 ;
	    RECT 105.4000 123.8000 105.8000 124.2000 ;
	    RECT 104.6000 122.8000 105.0000 123.2000 ;
	    RECT 106.2000 123.1000 106.6000 128.9000 ;
	    RECT 90.2000 118.8000 90.6000 119.2000 ;
	    RECT 91.0000 119.1000 91.4000 119.2000 ;
	    RECT 91.8000 119.1000 92.2000 119.2000 ;
	    RECT 91.0000 118.8000 92.2000 119.1000 ;
	    RECT 95.0000 118.8000 95.4000 119.2000 ;
	    RECT 88.6000 116.8000 89.0000 117.2000 ;
	    RECT 92.6000 116.8000 93.0000 117.2000 ;
	    RECT 92.6000 115.2000 92.9000 116.8000 ;
	    RECT 92.6000 114.8000 93.0000 115.2000 ;
	    RECT 93.4000 112.1000 93.8000 117.9000 ;
	    RECT 97.4000 114.7000 97.8000 115.1000 ;
	    RECT 97.4000 111.2000 97.7000 114.7000 ;
	    RECT 98.2000 112.1000 98.6000 117.9000 ;
	    RECT 99.0000 113.8000 99.4000 114.2000 ;
	    RECT 97.4000 110.8000 97.8000 111.2000 ;
	    RECT 81.4000 109.8000 81.8000 110.2000 ;
	    RECT 67.0000 108.8000 67.4000 109.2000 ;
	    RECT 70.2000 108.8000 70.6000 109.2000 ;
	    RECT 72.6000 108.8000 73.0000 109.2000 ;
	    RECT 62.2000 107.8000 62.6000 108.2000 ;
	    RECT 58.2000 106.8000 59.3000 107.1000 ;
	    RECT 62.2000 106.8000 62.6000 107.2000 ;
	    RECT 43.8000 106.2000 44.1000 106.8000 ;
	    RECT 54.2000 106.2000 54.5000 106.8000 ;
	    RECT 43.8000 105.8000 44.2000 106.2000 ;
	    RECT 49.4000 106.1000 49.8000 106.2000 ;
	    RECT 50.2000 106.1000 50.6000 106.2000 ;
	    RECT 49.4000 105.8000 50.6000 106.1000 ;
	    RECT 54.2000 105.8000 54.6000 106.2000 ;
	    RECT 55.0000 106.1000 55.4000 106.2000 ;
	    RECT 55.8000 106.1000 56.2000 106.2000 ;
	    RECT 55.0000 105.8000 56.2000 106.1000 ;
	    RECT 57.4000 106.1000 57.8000 106.2000 ;
	    RECT 58.2000 106.1000 58.6000 106.2000 ;
	    RECT 57.4000 105.8000 58.6000 106.1000 ;
	    RECT 47.8000 104.8000 48.2000 105.2000 ;
	    RECT 55.8000 104.8000 56.2000 105.2000 ;
	    RECT 58.2000 104.8000 58.6000 105.2000 ;
	    RECT 59.8000 105.1000 60.2000 105.2000 ;
	    RECT 59.0000 104.8000 60.2000 105.1000 ;
	    RECT 47.8000 104.2000 48.1000 104.8000 ;
	    RECT 47.8000 103.8000 48.2000 104.2000 ;
	    RECT 48.6000 104.1000 49.0000 104.2000 ;
	    RECT 49.4000 104.1000 49.8000 104.2000 ;
	    RECT 48.6000 103.8000 49.8000 104.1000 ;
	    RECT 50.2000 103.8000 50.6000 104.2000 ;
	    RECT 50.2000 103.2000 50.5000 103.8000 ;
	    RECT 50.2000 102.8000 50.6000 103.2000 ;
	    RECT 47.8000 99.8000 48.2000 100.2000 ;
	    RECT 47.8000 99.2000 48.1000 99.8000 ;
	    RECT 47.8000 98.8000 48.2000 99.2000 ;
	    RECT 42.2000 97.8000 43.3000 98.1000 ;
	    RECT 42.2000 96.8000 42.6000 97.2000 ;
	    RECT 42.2000 96.2000 42.5000 96.8000 ;
	    RECT 38.2000 96.1000 38.6000 96.2000 ;
	    RECT 37.4000 95.8000 38.6000 96.1000 ;
	    RECT 42.2000 95.8000 42.6000 96.2000 ;
	    RECT 32.6000 95.2000 32.9000 95.8000 ;
	    RECT 32.6000 94.8000 33.0000 95.2000 ;
	    RECT 36.6000 95.1000 37.0000 95.2000 ;
	    RECT 37.4000 95.1000 37.8000 95.2000 ;
	    RECT 36.6000 94.8000 37.8000 95.1000 ;
	    RECT 31.8000 93.8000 32.9000 94.1000 ;
	    RECT 32.6000 89.2000 32.9000 93.8000 ;
	    RECT 37.4000 93.8000 37.8000 94.2000 ;
	    RECT 37.4000 93.2000 37.7000 93.8000 ;
	    RECT 34.2000 93.1000 34.6000 93.2000 ;
	    RECT 35.0000 93.1000 35.4000 93.2000 ;
	    RECT 34.2000 92.8000 35.4000 93.1000 ;
	    RECT 37.4000 92.8000 37.8000 93.2000 ;
	    RECT 32.6000 88.8000 33.0000 89.2000 ;
	    RECT 34.2000 88.2000 34.5000 92.8000 ;
	    RECT 38.2000 88.2000 38.5000 95.8000 ;
	    RECT 43.0000 94.2000 43.3000 97.8000 ;
	    RECT 46.2000 97.1000 46.6000 97.2000 ;
	    RECT 47.0000 97.1000 47.4000 97.2000 ;
	    RECT 46.2000 96.8000 47.4000 97.1000 ;
	    RECT 52.6000 96.8000 53.0000 97.2000 ;
	    RECT 52.6000 96.2000 52.9000 96.8000 ;
	    RECT 55.8000 96.2000 56.1000 104.8000 ;
	    RECT 58.2000 104.2000 58.5000 104.8000 ;
	    RECT 56.6000 104.1000 57.0000 104.2000 ;
	    RECT 57.4000 104.1000 57.8000 104.2000 ;
	    RECT 56.6000 103.8000 57.8000 104.1000 ;
	    RECT 58.2000 103.8000 58.6000 104.2000 ;
	    RECT 59.0000 99.1000 59.3000 104.8000 ;
	    RECT 62.2000 104.1000 62.5000 106.8000 ;
	    RECT 67.0000 106.2000 67.3000 108.8000 ;
	    RECT 63.0000 106.1000 63.4000 106.2000 ;
	    RECT 63.8000 106.1000 64.2000 106.2000 ;
	    RECT 63.0000 105.8000 64.2000 106.1000 ;
	    RECT 64.6000 105.8000 65.0000 106.2000 ;
	    RECT 67.0000 105.8000 67.4000 106.2000 ;
	    RECT 67.8000 105.8000 68.2000 106.2000 ;
	    RECT 70.2000 105.8000 70.6000 106.2000 ;
	    RECT 73.4000 105.8000 73.8000 106.2000 ;
	    RECT 75.8000 105.8000 76.2000 106.2000 ;
	    RECT 79.0000 105.8000 79.4000 106.2000 ;
	    RECT 64.6000 105.2000 64.9000 105.8000 ;
	    RECT 67.8000 105.2000 68.1000 105.8000 ;
	    RECT 63.8000 104.8000 64.2000 105.2000 ;
	    RECT 64.6000 104.8000 65.0000 105.2000 ;
	    RECT 67.8000 105.1000 68.2000 105.2000 ;
	    RECT 68.6000 105.1000 69.0000 105.2000 ;
	    RECT 67.8000 104.8000 69.0000 105.1000 ;
	    RECT 63.0000 104.1000 63.4000 104.2000 ;
	    RECT 62.2000 103.8000 63.4000 104.1000 ;
	    RECT 63.8000 103.2000 64.1000 104.8000 ;
	    RECT 66.2000 103.8000 66.6000 104.2000 ;
	    RECT 67.0000 103.8000 67.4000 104.2000 ;
	    RECT 69.4000 104.1000 69.8000 104.2000 ;
	    RECT 68.6000 103.8000 69.8000 104.1000 ;
	    RECT 66.2000 103.2000 66.5000 103.8000 ;
	    RECT 67.0000 103.2000 67.3000 103.8000 ;
	    RECT 63.8000 102.8000 64.2000 103.2000 ;
	    RECT 66.2000 102.8000 66.6000 103.2000 ;
	    RECT 67.0000 102.8000 67.4000 103.2000 ;
	    RECT 59.8000 99.1000 60.2000 99.2000 ;
	    RECT 59.0000 98.8000 60.2000 99.1000 ;
	    RECT 57.4000 97.1000 57.8000 97.2000 ;
	    RECT 58.2000 97.1000 58.6000 97.2000 ;
	    RECT 57.4000 96.8000 58.6000 97.1000 ;
	    RECT 59.8000 97.1000 60.2000 97.2000 ;
	    RECT 60.6000 97.1000 61.0000 97.2000 ;
	    RECT 59.8000 96.8000 61.0000 97.1000 ;
	    RECT 66.2000 96.8000 66.6000 97.2000 ;
	    RECT 66.2000 96.2000 66.5000 96.8000 ;
	    RECT 45.4000 95.8000 45.8000 96.2000 ;
	    RECT 47.8000 96.1000 48.2000 96.2000 ;
	    RECT 48.6000 96.1000 49.0000 96.2000 ;
	    RECT 47.8000 95.8000 49.0000 96.1000 ;
	    RECT 52.6000 95.8000 53.0000 96.2000 ;
	    RECT 55.8000 96.1000 56.2000 96.2000 ;
	    RECT 56.6000 96.1000 57.0000 96.2000 ;
	    RECT 55.8000 95.8000 57.0000 96.1000 ;
	    RECT 66.2000 95.8000 66.6000 96.2000 ;
	    RECT 45.4000 95.2000 45.7000 95.8000 ;
	    RECT 43.8000 94.8000 44.2000 95.2000 ;
	    RECT 45.4000 94.8000 45.8000 95.2000 ;
	    RECT 47.0000 95.1000 47.4000 95.2000 ;
	    RECT 47.8000 95.1000 48.2000 95.2000 ;
	    RECT 47.0000 94.8000 48.2000 95.1000 ;
	    RECT 55.8000 94.8000 56.2000 95.2000 ;
	    RECT 56.6000 95.1000 57.0000 95.2000 ;
	    RECT 57.4000 95.1000 57.8000 95.2000 ;
	    RECT 56.6000 94.8000 57.8000 95.1000 ;
	    RECT 43.8000 94.2000 44.1000 94.8000 ;
	    RECT 55.8000 94.2000 56.1000 94.8000 ;
	    RECT 43.0000 94.1000 43.4000 94.2000 ;
	    RECT 43.8000 94.1000 44.2000 94.2000 ;
	    RECT 43.0000 93.8000 44.2000 94.1000 ;
	    RECT 51.8000 94.1000 52.2000 94.2000 ;
	    RECT 52.6000 94.1000 53.0000 94.2000 ;
	    RECT 51.8000 93.8000 53.0000 94.1000 ;
	    RECT 55.8000 93.8000 56.2000 94.2000 ;
	    RECT 66.2000 93.8000 66.6000 94.2000 ;
	    RECT 66.2000 88.2000 66.5000 93.8000 ;
	    RECT 68.6000 89.2000 68.9000 103.8000 ;
	    RECT 70.2000 103.1000 70.5000 105.8000 ;
	    RECT 69.4000 102.8000 70.5000 103.1000 ;
	    RECT 69.4000 97.2000 69.7000 102.8000 ;
	    RECT 70.2000 102.1000 70.6000 102.2000 ;
	    RECT 71.0000 102.1000 71.4000 102.2000 ;
	    RECT 70.2000 101.8000 71.4000 102.1000 ;
	    RECT 71.8000 97.8000 72.2000 98.2000 ;
	    RECT 71.8000 97.2000 72.1000 97.8000 ;
	    RECT 69.4000 96.8000 69.8000 97.2000 ;
	    RECT 71.0000 96.8000 71.4000 97.2000 ;
	    RECT 71.8000 96.8000 72.2000 97.2000 ;
	    RECT 71.0000 96.2000 71.3000 96.8000 ;
	    RECT 71.0000 95.8000 71.4000 96.2000 ;
	    RECT 71.8000 94.8000 72.2000 95.2000 ;
	    RECT 71.8000 94.2000 72.1000 94.8000 ;
	    RECT 69.4000 94.1000 69.8000 94.2000 ;
	    RECT 70.2000 94.1000 70.6000 94.2000 ;
	    RECT 69.4000 93.8000 70.6000 94.1000 ;
	    RECT 71.8000 93.8000 72.2000 94.2000 ;
	    RECT 68.6000 88.8000 69.0000 89.2000 ;
	    RECT 26.2000 87.8000 26.6000 88.2000 ;
	    RECT 31.0000 87.8000 31.4000 88.2000 ;
	    RECT 34.2000 87.8000 34.6000 88.2000 ;
	    RECT 35.8000 87.8000 36.2000 88.2000 ;
	    RECT 36.6000 88.1000 37.0000 88.2000 ;
	    RECT 37.4000 88.1000 37.8000 88.2000 ;
	    RECT 36.6000 87.8000 37.8000 88.1000 ;
	    RECT 38.2000 87.8000 38.6000 88.2000 ;
	    RECT 43.8000 87.8000 44.2000 88.2000 ;
	    RECT 48.6000 87.8000 49.0000 88.2000 ;
	    RECT 51.0000 88.1000 51.4000 88.2000 ;
	    RECT 51.8000 88.1000 52.2000 88.2000 ;
	    RECT 51.0000 87.8000 52.2000 88.1000 ;
	    RECT 57.4000 88.1000 57.8000 88.2000 ;
	    RECT 58.2000 88.1000 58.6000 88.2000 ;
	    RECT 57.4000 87.8000 58.6000 88.1000 ;
	    RECT 66.2000 87.8000 66.6000 88.2000 ;
	    RECT 72.6000 87.8000 73.0000 88.2000 ;
	    RECT 31.0000 87.2000 31.3000 87.8000 ;
	    RECT 34.2000 87.2000 34.5000 87.8000 ;
	    RECT 24.6000 86.8000 25.0000 87.2000 ;
	    RECT 31.0000 86.8000 31.4000 87.2000 ;
	    RECT 34.2000 86.8000 34.6000 87.2000 ;
	    RECT 23.8000 85.8000 24.2000 86.2000 ;
	    RECT 24.6000 86.1000 24.9000 86.8000 ;
	    RECT 25.4000 86.1000 25.8000 86.2000 ;
	    RECT 24.6000 85.8000 25.8000 86.1000 ;
	    RECT 27.0000 86.1000 27.4000 86.2000 ;
	    RECT 27.8000 86.1000 28.2000 86.2000 ;
	    RECT 27.0000 85.8000 28.2000 86.1000 ;
	    RECT 30.2000 85.8000 30.6000 86.2000 ;
	    RECT 31.0000 86.1000 31.4000 86.2000 ;
	    RECT 31.8000 86.1000 32.2000 86.2000 ;
	    RECT 31.0000 85.8000 32.2000 86.1000 ;
	    RECT 34.2000 85.8000 34.6000 86.2000 ;
	    RECT 15.0000 84.8000 15.4000 85.2000 ;
	    RECT 17.4000 84.8000 17.8000 85.2000 ;
	    RECT 18.2000 85.1000 18.6000 85.2000 ;
	    RECT 19.0000 85.1000 19.4000 85.2000 ;
	    RECT 18.2000 84.8000 19.4000 85.1000 ;
	    RECT 23.0000 84.8000 23.4000 85.2000 ;
	    RECT 9.4000 84.1000 9.8000 84.2000 ;
	    RECT 10.2000 84.1000 10.6000 84.2000 ;
	    RECT 9.4000 83.8000 10.6000 84.1000 ;
	    RECT 13.4000 83.8000 13.8000 84.2000 ;
	    RECT 13.4000 82.2000 13.7000 83.8000 ;
	    RECT 10.2000 82.1000 10.6000 82.2000 ;
	    RECT 11.0000 82.1000 11.4000 82.2000 ;
	    RECT 10.2000 81.8000 11.4000 82.1000 ;
	    RECT 13.4000 81.8000 13.8000 82.2000 ;
	    RECT 14.2000 81.8000 14.6000 82.2000 ;
	    RECT 4.6000 76.8000 5.0000 77.2000 ;
	    RECT 14.2000 75.2000 14.5000 81.8000 ;
	    RECT 14.2000 74.8000 14.6000 75.2000 ;
	    RECT 2.2000 73.8000 2.6000 74.2000 ;
	    RECT 10.2000 73.8000 10.6000 74.2000 ;
	    RECT 13.4000 74.1000 13.8000 74.2000 ;
	    RECT 14.2000 74.1000 14.6000 74.2000 ;
	    RECT 13.4000 73.8000 14.6000 74.1000 ;
	    RECT 2.2000 73.2000 2.5000 73.8000 ;
	    RECT 10.2000 73.2000 10.5000 73.8000 ;
	    RECT 2.2000 72.8000 2.6000 73.2000 ;
	    RECT 4.6000 73.1000 5.0000 73.2000 ;
	    RECT 5.4000 73.1000 5.8000 73.2000 ;
	    RECT 4.6000 72.8000 5.8000 73.1000 ;
	    RECT 10.2000 72.8000 10.6000 73.2000 ;
	    RECT 1.4000 71.8000 1.8000 72.2000 ;
	    RECT 3.0000 71.8000 3.4000 72.2000 ;
	    RECT 4.6000 71.8000 5.0000 72.2000 ;
	    RECT 7.8000 71.8000 8.2000 72.2000 ;
	    RECT 1.4000 64.2000 1.7000 71.8000 ;
	    RECT 2.2000 66.1000 2.6000 66.2000 ;
	    RECT 3.0000 66.1000 3.3000 71.8000 ;
	    RECT 4.6000 69.2000 4.9000 71.8000 ;
	    RECT 5.4000 70.8000 5.8000 71.2000 ;
	    RECT 4.6000 68.8000 5.0000 69.2000 ;
	    RECT 5.4000 68.2000 5.7000 70.8000 ;
	    RECT 7.8000 68.2000 8.1000 71.8000 ;
	    RECT 10.2000 71.2000 10.5000 72.8000 ;
	    RECT 15.0000 72.2000 15.3000 84.8000 ;
	    RECT 30.2000 84.2000 30.5000 85.8000 ;
	    RECT 34.2000 85.2000 34.5000 85.8000 ;
	    RECT 31.0000 85.1000 31.4000 85.2000 ;
	    RECT 31.8000 85.1000 32.2000 85.2000 ;
	    RECT 31.0000 84.8000 32.2000 85.1000 ;
	    RECT 32.6000 85.1000 33.0000 85.2000 ;
	    RECT 32.6000 84.8000 33.7000 85.1000 ;
	    RECT 34.2000 84.8000 34.6000 85.2000 ;
	    RECT 24.6000 84.1000 25.0000 84.2000 ;
	    RECT 24.6000 83.8000 25.7000 84.1000 ;
	    RECT 25.4000 83.1000 25.7000 83.8000 ;
	    RECT 27.8000 83.8000 28.2000 84.2000 ;
	    RECT 30.2000 83.8000 30.6000 84.2000 ;
	    RECT 27.0000 83.1000 27.4000 83.2000 ;
	    RECT 25.4000 82.8000 27.4000 83.1000 ;
	    RECT 27.8000 75.2000 28.1000 83.8000 ;
	    RECT 33.4000 79.2000 33.7000 84.8000 ;
	    RECT 33.4000 78.8000 33.8000 79.2000 ;
	    RECT 35.8000 75.2000 36.1000 87.8000 ;
	    RECT 41.4000 86.8000 41.8000 87.2000 ;
	    RECT 41.4000 86.2000 41.7000 86.8000 ;
	    RECT 41.4000 85.8000 41.8000 86.2000 ;
	    RECT 43.8000 85.2000 44.1000 87.8000 ;
	    RECT 48.6000 87.2000 48.9000 87.8000 ;
	    RECT 66.2000 87.2000 66.5000 87.8000 ;
	    RECT 72.6000 87.2000 72.9000 87.8000 ;
	    RECT 48.6000 86.8000 49.0000 87.2000 ;
	    RECT 53.4000 86.8000 53.8000 87.2000 ;
	    RECT 66.2000 86.8000 66.6000 87.2000 ;
	    RECT 72.6000 86.8000 73.0000 87.2000 ;
	    RECT 53.4000 86.2000 53.7000 86.8000 ;
	    RECT 44.6000 85.8000 45.0000 86.2000 ;
	    RECT 48.6000 85.8000 49.0000 86.2000 ;
	    RECT 53.4000 85.8000 53.8000 86.2000 ;
	    RECT 55.0000 86.1000 55.4000 86.2000 ;
	    RECT 55.8000 86.1000 56.2000 86.2000 ;
	    RECT 55.0000 85.8000 56.2000 86.1000 ;
	    RECT 61.4000 86.1000 61.8000 86.2000 ;
	    RECT 62.2000 86.1000 62.6000 86.2000 ;
	    RECT 61.4000 85.8000 62.6000 86.1000 ;
	    RECT 71.8000 86.1000 72.2000 86.2000 ;
	    RECT 72.6000 86.1000 73.0000 86.2000 ;
	    RECT 71.8000 85.8000 73.0000 86.1000 ;
	    RECT 44.6000 85.2000 44.9000 85.8000 ;
	    RECT 48.6000 85.2000 48.9000 85.8000 ;
	    RECT 73.4000 85.2000 73.7000 105.8000 ;
	    RECT 75.8000 105.2000 76.1000 105.8000 ;
	    RECT 75.8000 104.8000 76.2000 105.2000 ;
	    RECT 77.4000 104.1000 77.8000 104.2000 ;
	    RECT 78.2000 104.1000 78.6000 104.2000 ;
	    RECT 77.4000 103.8000 78.6000 104.1000 ;
	    RECT 79.0000 103.2000 79.3000 105.8000 ;
	    RECT 79.8000 105.1000 80.2000 105.2000 ;
	    RECT 80.6000 105.1000 81.0000 105.2000 ;
	    RECT 79.8000 104.8000 81.0000 105.1000 ;
	    RECT 81.4000 104.2000 81.7000 109.8000 ;
	    RECT 82.2000 106.8000 82.6000 107.2000 ;
	    RECT 89.4000 106.8000 89.8000 107.2000 ;
	    RECT 82.2000 106.2000 82.5000 106.8000 ;
	    RECT 89.4000 106.2000 89.7000 106.8000 ;
	    RECT 82.2000 105.8000 82.6000 106.2000 ;
	    RECT 83.8000 105.8000 84.2000 106.2000 ;
	    RECT 84.6000 105.8000 85.0000 106.2000 ;
	    RECT 87.0000 105.8000 87.4000 106.2000 ;
	    RECT 87.8000 105.8000 88.2000 106.2000 ;
	    RECT 89.4000 105.8000 89.8000 106.2000 ;
	    RECT 91.0000 106.1000 91.4000 106.2000 ;
	    RECT 91.8000 106.1000 92.2000 106.2000 ;
	    RECT 91.0000 105.8000 92.2000 106.1000 ;
	    RECT 83.8000 105.2000 84.1000 105.8000 ;
	    RECT 82.2000 105.1000 82.6000 105.2000 ;
	    RECT 83.0000 105.1000 83.4000 105.2000 ;
	    RECT 82.2000 104.8000 83.4000 105.1000 ;
	    RECT 83.8000 104.8000 84.2000 105.2000 ;
	    RECT 84.6000 104.2000 84.9000 105.8000 ;
	    RECT 87.0000 105.2000 87.3000 105.8000 ;
	    RECT 87.0000 104.8000 87.4000 105.2000 ;
	    RECT 81.4000 103.8000 81.8000 104.2000 ;
	    RECT 84.6000 103.8000 85.0000 104.2000 ;
	    RECT 85.4000 103.8000 85.8000 104.2000 ;
	    RECT 87.8000 104.1000 88.1000 105.8000 ;
	    RECT 92.6000 104.8000 93.0000 105.2000 ;
	    RECT 93.4000 105.1000 93.8000 107.9000 ;
	    RECT 92.6000 104.2000 92.9000 104.8000 ;
	    RECT 87.0000 103.8000 88.1000 104.1000 ;
	    RECT 88.6000 103.8000 89.0000 104.2000 ;
	    RECT 91.0000 103.8000 91.4000 104.2000 ;
	    RECT 92.6000 103.8000 93.0000 104.2000 ;
	    RECT 85.4000 103.2000 85.7000 103.8000 ;
	    RECT 79.0000 102.8000 79.4000 103.2000 ;
	    RECT 85.4000 102.8000 85.8000 103.2000 ;
	    RECT 75.0000 101.8000 75.4000 102.2000 ;
	    RECT 79.0000 101.8000 79.4000 102.2000 ;
	    RECT 82.2000 101.8000 82.6000 102.2000 ;
	    RECT 86.2000 101.8000 86.6000 102.2000 ;
	    RECT 74.2000 97.8000 74.6000 98.2000 ;
	    RECT 74.2000 97.2000 74.5000 97.8000 ;
	    RECT 74.2000 96.8000 74.6000 97.2000 ;
	    RECT 75.0000 96.2000 75.3000 101.8000 ;
	    RECT 79.0000 100.2000 79.3000 101.8000 ;
	    RECT 82.2000 101.2000 82.5000 101.8000 ;
	    RECT 82.2000 100.8000 82.6000 101.2000 ;
	    RECT 79.0000 99.8000 79.4000 100.2000 ;
	    RECT 83.8000 99.1000 84.2000 99.2000 ;
	    RECT 84.6000 99.1000 85.0000 99.2000 ;
	    RECT 83.8000 98.8000 85.0000 99.1000 ;
	    RECT 85.4000 97.8000 85.8000 98.2000 ;
	    RECT 85.4000 97.2000 85.7000 97.8000 ;
	    RECT 81.4000 96.8000 81.8000 97.2000 ;
	    RECT 83.0000 97.1000 83.4000 97.2000 ;
	    RECT 83.8000 97.1000 84.2000 97.2000 ;
	    RECT 83.0000 96.8000 84.2000 97.1000 ;
	    RECT 85.4000 96.8000 85.8000 97.2000 ;
	    RECT 81.4000 96.2000 81.7000 96.8000 ;
	    RECT 75.0000 95.8000 75.4000 96.2000 ;
	    RECT 79.8000 96.1000 80.2000 96.2000 ;
	    RECT 80.6000 96.1000 81.0000 96.2000 ;
	    RECT 79.8000 95.8000 81.0000 96.1000 ;
	    RECT 81.4000 95.8000 81.8000 96.2000 ;
	    RECT 83.8000 96.1000 84.2000 96.2000 ;
	    RECT 84.6000 96.1000 85.0000 96.2000 ;
	    RECT 83.8000 95.8000 85.0000 96.1000 ;
	    RECT 86.2000 95.2000 86.5000 101.8000 ;
	    RECT 87.0000 99.2000 87.3000 103.8000 ;
	    RECT 87.8000 102.8000 88.2000 103.2000 ;
	    RECT 87.8000 99.2000 88.1000 102.8000 ;
	    RECT 88.6000 100.2000 88.9000 103.8000 ;
	    RECT 91.0000 103.2000 91.3000 103.8000 ;
	    RECT 91.0000 102.8000 91.4000 103.2000 ;
	    RECT 95.0000 103.1000 95.4000 108.9000 ;
	    RECT 99.0000 106.2000 99.3000 113.8000 ;
	    RECT 99.8000 113.1000 100.2000 115.9000 ;
	    RECT 100.6000 111.8000 101.0000 112.2000 ;
	    RECT 103.0000 112.1000 103.4000 117.9000 ;
	    RECT 107.0000 115.1000 107.3000 142.8000 ;
	    RECT 108.6000 134.8000 109.0000 135.2000 ;
	    RECT 109.4000 134.8000 109.8000 135.2000 ;
	    RECT 108.6000 134.2000 108.9000 134.8000 ;
	    RECT 109.4000 134.2000 109.7000 134.8000 ;
	    RECT 111.0000 134.2000 111.3000 145.8000 ;
	    RECT 113.4000 145.2000 113.7000 145.8000 ;
	    RECT 113.4000 144.8000 113.8000 145.2000 ;
	    RECT 112.6000 143.8000 113.0000 144.2000 ;
	    RECT 113.4000 144.1000 113.7000 144.8000 ;
	    RECT 115.0000 144.2000 115.3000 145.8000 ;
	    RECT 116.6000 145.2000 116.9000 147.8000 ;
	    RECT 117.4000 147.2000 117.7000 149.8000 ;
	    RECT 119.8000 149.2000 120.1000 149.8000 ;
	    RECT 119.8000 148.8000 120.2000 149.2000 ;
	    RECT 120.6000 148.1000 120.9000 151.8000 ;
	    RECT 119.8000 147.8000 120.9000 148.1000 ;
	    RECT 121.4000 148.2000 121.7000 153.8000 ;
	    RECT 122.2000 153.2000 122.5000 154.8000 ;
	    RECT 123.0000 153.8000 123.4000 154.2000 ;
	    RECT 123.8000 153.8000 124.2000 154.2000 ;
	    RECT 131.0000 153.8000 131.4000 154.2000 ;
	    RECT 123.0000 153.2000 123.3000 153.8000 ;
	    RECT 122.2000 152.8000 122.6000 153.2000 ;
	    RECT 123.0000 152.8000 123.4000 153.2000 ;
	    RECT 122.2000 151.8000 122.6000 152.2000 ;
	    RECT 121.4000 147.8000 121.8000 148.2000 ;
	    RECT 117.4000 146.8000 117.8000 147.2000 ;
	    RECT 118.2000 145.8000 118.6000 146.2000 ;
	    RECT 118.2000 145.2000 118.5000 145.8000 ;
	    RECT 119.8000 145.2000 120.1000 147.8000 ;
	    RECT 120.6000 146.8000 121.0000 147.2000 ;
	    RECT 120.6000 146.2000 120.9000 146.8000 ;
	    RECT 122.2000 146.2000 122.5000 151.8000 ;
	    RECT 123.0000 147.2000 123.3000 152.8000 ;
	    RECT 123.8000 152.2000 124.1000 153.8000 ;
	    RECT 124.6000 153.1000 125.0000 153.2000 ;
	    RECT 125.4000 153.1000 125.8000 153.2000 ;
	    RECT 124.6000 152.8000 125.8000 153.1000 ;
	    RECT 128.6000 152.8000 129.0000 153.2000 ;
	    RECT 130.2000 153.1000 130.6000 153.2000 ;
	    RECT 131.0000 153.1000 131.3000 153.8000 ;
	    RECT 130.2000 152.8000 131.3000 153.1000 ;
	    RECT 131.8000 153.2000 132.1000 154.8000 ;
	    RECT 132.6000 154.2000 132.9000 154.8000 ;
	    RECT 132.6000 153.8000 133.0000 154.2000 ;
	    RECT 135.0000 153.8000 135.4000 154.2000 ;
	    RECT 131.8000 152.8000 132.2000 153.2000 ;
	    RECT 132.6000 153.1000 133.0000 153.2000 ;
	    RECT 133.4000 153.1000 133.8000 153.2000 ;
	    RECT 132.6000 152.8000 133.8000 153.1000 ;
	    RECT 134.2000 152.8000 134.6000 153.2000 ;
	    RECT 123.8000 151.8000 124.2000 152.2000 ;
	    RECT 127.0000 150.8000 127.4000 151.2000 ;
	    RECT 123.8000 148.8000 124.2000 149.2000 ;
	    RECT 123.0000 146.8000 123.4000 147.2000 ;
	    RECT 120.6000 145.8000 121.0000 146.2000 ;
	    RECT 122.2000 145.8000 122.6000 146.2000 ;
	    RECT 115.8000 144.8000 116.2000 145.2000 ;
	    RECT 116.6000 144.8000 117.0000 145.2000 ;
	    RECT 118.2000 144.8000 118.6000 145.2000 ;
	    RECT 119.8000 144.8000 120.2000 145.2000 ;
	    RECT 120.6000 144.8000 121.0000 145.2000 ;
	    RECT 113.4000 143.8000 114.5000 144.1000 ;
	    RECT 115.0000 143.8000 115.4000 144.2000 ;
	    RECT 112.6000 139.2000 112.9000 143.8000 ;
	    RECT 113.4000 139.8000 113.8000 140.2000 ;
	    RECT 113.4000 139.2000 113.7000 139.8000 ;
	    RECT 112.6000 138.8000 113.0000 139.2000 ;
	    RECT 113.4000 138.8000 113.8000 139.2000 ;
	    RECT 107.8000 133.8000 108.2000 134.2000 ;
	    RECT 108.6000 133.8000 109.0000 134.2000 ;
	    RECT 109.4000 133.8000 109.8000 134.2000 ;
	    RECT 111.0000 133.8000 111.4000 134.2000 ;
	    RECT 107.8000 133.2000 108.1000 133.8000 ;
	    RECT 111.0000 133.2000 111.3000 133.8000 ;
	    RECT 107.8000 132.8000 108.2000 133.2000 ;
	    RECT 111.0000 132.8000 111.4000 133.2000 ;
	    RECT 110.2000 126.8000 110.6000 127.2000 ;
	    RECT 110.2000 126.3000 110.5000 126.8000 ;
	    RECT 110.2000 125.9000 110.6000 126.3000 ;
	    RECT 111.0000 123.1000 111.4000 128.9000 ;
	    RECT 111.8000 127.8000 112.2000 128.2000 ;
	    RECT 111.8000 127.2000 112.1000 127.8000 ;
	    RECT 111.8000 126.8000 112.2000 127.2000 ;
	    RECT 112.6000 125.1000 113.0000 127.9000 ;
	    RECT 114.2000 122.2000 114.5000 143.8000 ;
	    RECT 115.8000 143.2000 116.1000 144.8000 ;
	    RECT 120.6000 144.2000 120.9000 144.8000 ;
	    RECT 120.6000 143.8000 121.0000 144.2000 ;
	    RECT 115.8000 142.8000 116.2000 143.2000 ;
	    RECT 120.6000 135.2000 120.9000 143.8000 ;
	    RECT 122.2000 142.2000 122.5000 145.8000 ;
	    RECT 123.8000 145.2000 124.1000 148.8000 ;
	    RECT 127.0000 148.2000 127.3000 150.8000 ;
	    RECT 128.6000 148.2000 128.9000 152.8000 ;
	    RECT 134.2000 152.2000 134.5000 152.8000 ;
	    RECT 134.2000 151.8000 134.6000 152.2000 ;
	    RECT 127.0000 147.8000 127.4000 148.2000 ;
	    RECT 128.6000 147.8000 129.0000 148.2000 ;
	    RECT 125.4000 146.8000 125.8000 147.2000 ;
	    RECT 129.4000 146.8000 129.8000 147.2000 ;
	    RECT 132.6000 146.8000 133.0000 147.2000 ;
	    RECT 125.4000 146.2000 125.7000 146.8000 ;
	    RECT 124.6000 145.8000 125.0000 146.2000 ;
	    RECT 125.4000 145.8000 125.8000 146.2000 ;
	    RECT 127.0000 145.8000 127.4000 146.2000 ;
	    RECT 123.8000 144.8000 124.2000 145.2000 ;
	    RECT 122.2000 141.8000 122.6000 142.2000 ;
	    RECT 124.6000 136.2000 124.9000 145.8000 ;
	    RECT 127.0000 145.2000 127.3000 145.8000 ;
	    RECT 127.0000 144.8000 127.4000 145.2000 ;
	    RECT 125.4000 143.8000 125.8000 144.2000 ;
	    RECT 125.4000 137.1000 125.7000 143.8000 ;
	    RECT 128.6000 141.8000 129.0000 142.2000 ;
	    RECT 128.6000 141.2000 128.9000 141.8000 ;
	    RECT 128.6000 140.8000 129.0000 141.2000 ;
	    RECT 128.6000 139.2000 128.9000 140.8000 ;
	    RECT 127.0000 139.1000 127.4000 139.2000 ;
	    RECT 127.8000 139.1000 128.2000 139.2000 ;
	    RECT 127.0000 138.8000 128.2000 139.1000 ;
	    RECT 128.6000 138.8000 129.0000 139.2000 ;
	    RECT 129.4000 138.2000 129.7000 146.8000 ;
	    RECT 132.6000 146.2000 132.9000 146.8000 ;
	    RECT 131.8000 145.8000 132.2000 146.2000 ;
	    RECT 132.6000 145.8000 133.0000 146.2000 ;
	    RECT 130.2000 144.8000 130.6000 145.2000 ;
	    RECT 130.2000 140.2000 130.5000 144.8000 ;
	    RECT 131.8000 144.2000 132.1000 145.8000 ;
	    RECT 131.8000 143.8000 132.2000 144.2000 ;
	    RECT 132.6000 141.8000 133.0000 142.2000 ;
	    RECT 130.2000 139.8000 130.6000 140.2000 ;
	    RECT 132.6000 139.2000 132.9000 141.8000 ;
	    RECT 135.0000 139.2000 135.3000 153.8000 ;
	    RECT 136.6000 149.2000 136.9000 155.8000 ;
	    RECT 143.0000 155.2000 143.3000 155.8000 ;
	    RECT 138.2000 154.8000 138.6000 155.2000 ;
	    RECT 141.4000 154.8000 141.8000 155.2000 ;
	    RECT 143.0000 154.8000 143.4000 155.2000 ;
	    RECT 144.6000 154.8000 145.0000 155.2000 ;
	    RECT 137.4000 151.8000 137.8000 152.2000 ;
	    RECT 137.4000 151.2000 137.7000 151.8000 ;
	    RECT 137.4000 150.8000 137.8000 151.2000 ;
	    RECT 137.4000 149.2000 137.7000 150.8000 ;
	    RECT 136.6000 148.8000 137.0000 149.2000 ;
	    RECT 137.4000 148.8000 137.8000 149.2000 ;
	    RECT 136.6000 145.8000 137.0000 146.2000 ;
	    RECT 135.8000 144.8000 136.2000 145.2000 ;
	    RECT 135.8000 139.2000 136.1000 144.8000 ;
	    RECT 136.6000 140.2000 136.9000 145.8000 ;
	    RECT 138.2000 141.2000 138.5000 154.8000 ;
	    RECT 139.0000 153.8000 139.4000 154.2000 ;
	    RECT 139.0000 142.2000 139.3000 153.8000 ;
	    RECT 141.4000 153.2000 141.7000 154.8000 ;
	    RECT 142.2000 153.8000 142.6000 154.2000 ;
	    RECT 143.8000 153.8000 144.2000 154.2000 ;
	    RECT 142.2000 153.2000 142.5000 153.8000 ;
	    RECT 143.8000 153.2000 144.1000 153.8000 ;
	    RECT 141.4000 152.8000 141.8000 153.2000 ;
	    RECT 142.2000 152.8000 142.6000 153.2000 ;
	    RECT 143.8000 152.8000 144.2000 153.2000 ;
	    RECT 144.6000 152.2000 144.9000 154.8000 ;
	    RECT 144.6000 151.8000 145.0000 152.2000 ;
	    RECT 145.4000 151.1000 145.7000 155.8000 ;
	    RECT 144.6000 150.8000 145.7000 151.1000 ;
	    RECT 144.6000 149.2000 144.9000 150.8000 ;
	    RECT 146.2000 150.2000 146.5000 156.8000 ;
	    RECT 147.8000 156.2000 148.1000 156.8000 ;
	    RECT 147.0000 155.8000 147.4000 156.2000 ;
	    RECT 147.8000 155.8000 148.2000 156.2000 ;
	    RECT 147.0000 155.2000 147.3000 155.8000 ;
	    RECT 151.8000 155.2000 152.1000 156.8000 ;
	    RECT 159.0000 156.2000 159.3000 156.8000 ;
	    RECT 153.4000 155.8000 153.8000 156.2000 ;
	    RECT 155.0000 156.1000 155.4000 156.2000 ;
	    RECT 155.8000 156.1000 156.2000 156.2000 ;
	    RECT 155.0000 155.8000 156.2000 156.1000 ;
	    RECT 159.0000 155.8000 159.4000 156.2000 ;
	    RECT 161.4000 155.8000 161.8000 156.2000 ;
	    RECT 147.0000 154.8000 147.4000 155.2000 ;
	    RECT 147.8000 155.1000 148.2000 155.2000 ;
	    RECT 148.6000 155.1000 149.0000 155.2000 ;
	    RECT 147.8000 154.8000 149.0000 155.1000 ;
	    RECT 149.4000 154.8000 149.8000 155.2000 ;
	    RECT 151.8000 154.8000 152.2000 155.2000 ;
	    RECT 152.6000 154.8000 153.0000 155.2000 ;
	    RECT 147.0000 153.8000 147.4000 154.2000 ;
	    RECT 147.0000 153.2000 147.3000 153.8000 ;
	    RECT 147.0000 152.8000 147.4000 153.2000 ;
	    RECT 148.6000 151.2000 148.9000 154.8000 ;
	    RECT 148.6000 150.8000 149.0000 151.2000 ;
	    RECT 146.2000 149.8000 146.6000 150.2000 ;
	    RECT 149.4000 150.1000 149.7000 154.8000 ;
	    RECT 151.0000 154.1000 151.4000 154.2000 ;
	    RECT 151.8000 154.1000 152.2000 154.2000 ;
	    RECT 151.0000 153.8000 152.2000 154.1000 ;
	    RECT 152.6000 153.2000 152.9000 154.8000 ;
	    RECT 152.6000 152.8000 153.0000 153.2000 ;
	    RECT 153.4000 152.2000 153.7000 155.8000 ;
	    RECT 157.4000 154.8000 157.8000 155.2000 ;
	    RECT 159.0000 155.1000 159.4000 155.2000 ;
	    RECT 159.8000 155.1000 160.2000 155.2000 ;
	    RECT 159.0000 154.8000 160.2000 155.1000 ;
	    RECT 154.2000 154.1000 154.6000 154.2000 ;
	    RECT 155.0000 154.1000 155.4000 154.2000 ;
	    RECT 154.2000 153.8000 155.4000 154.1000 ;
	    RECT 156.6000 153.8000 157.0000 154.2000 ;
	    RECT 155.0000 152.8000 155.4000 153.2000 ;
	    RECT 153.4000 151.8000 153.8000 152.2000 ;
	    RECT 148.6000 149.8000 149.7000 150.1000 ;
	    RECT 154.2000 150.8000 154.6000 151.2000 ;
	    RECT 144.6000 148.8000 145.0000 149.2000 ;
	    RECT 146.2000 147.2000 146.5000 149.8000 ;
	    RECT 148.6000 149.2000 148.9000 149.8000 ;
	    RECT 148.6000 148.8000 149.0000 149.2000 ;
	    RECT 151.0000 147.8000 151.4000 148.2000 ;
	    RECT 139.8000 146.8000 140.2000 147.2000 ;
	    RECT 142.2000 147.1000 142.6000 147.2000 ;
	    RECT 143.0000 147.1000 143.4000 147.2000 ;
	    RECT 142.2000 146.8000 143.4000 147.1000 ;
	    RECT 143.8000 146.8000 144.2000 147.2000 ;
	    RECT 144.6000 147.1000 145.0000 147.2000 ;
	    RECT 145.4000 147.1000 145.8000 147.2000 ;
	    RECT 144.6000 146.8000 145.8000 147.1000 ;
	    RECT 146.2000 146.8000 146.6000 147.2000 ;
	    RECT 149.4000 146.8000 149.8000 147.2000 ;
	    RECT 139.8000 146.2000 140.1000 146.8000 ;
	    RECT 139.8000 145.8000 140.2000 146.2000 ;
	    RECT 140.6000 145.8000 141.0000 146.2000 ;
	    RECT 143.0000 145.8000 143.4000 146.2000 ;
	    RECT 140.6000 144.2000 140.9000 145.8000 ;
	    RECT 143.0000 145.2000 143.3000 145.8000 ;
	    RECT 142.2000 144.8000 142.6000 145.2000 ;
	    RECT 143.0000 144.8000 143.4000 145.2000 ;
	    RECT 140.6000 143.8000 141.0000 144.2000 ;
	    RECT 142.2000 143.2000 142.5000 144.8000 ;
	    RECT 142.2000 142.8000 142.6000 143.2000 ;
	    RECT 139.0000 141.8000 139.4000 142.2000 ;
	    RECT 143.8000 141.2000 144.1000 146.8000 ;
	    RECT 146.2000 145.8000 146.6000 146.2000 ;
	    RECT 138.2000 140.8000 138.6000 141.2000 ;
	    RECT 143.8000 140.8000 144.2000 141.2000 ;
	    RECT 136.6000 139.8000 137.0000 140.2000 ;
	    RECT 146.2000 139.2000 146.5000 145.8000 ;
	    RECT 149.4000 142.2000 149.7000 146.8000 ;
	    RECT 150.2000 145.8000 150.6000 146.2000 ;
	    RECT 149.4000 141.8000 149.8000 142.2000 ;
	    RECT 147.8000 139.8000 148.2000 140.2000 ;
	    RECT 132.6000 138.8000 133.0000 139.2000 ;
	    RECT 135.0000 138.8000 135.4000 139.2000 ;
	    RECT 135.8000 138.8000 136.2000 139.2000 ;
	    RECT 139.0000 138.8000 139.4000 139.2000 ;
	    RECT 146.2000 138.8000 146.6000 139.2000 ;
	    RECT 139.0000 138.2000 139.3000 138.8000 ;
	    RECT 129.4000 137.8000 129.8000 138.2000 ;
	    RECT 139.0000 137.8000 139.4000 138.2000 ;
	    RECT 126.2000 137.1000 126.6000 137.2000 ;
	    RECT 127.0000 137.1000 127.4000 137.2000 ;
	    RECT 125.4000 136.8000 127.4000 137.1000 ;
	    RECT 137.4000 136.8000 137.8000 137.2000 ;
	    RECT 147.0000 136.8000 147.4000 137.2000 ;
	    RECT 137.4000 136.2000 137.7000 136.8000 ;
	    RECT 123.8000 135.8000 124.2000 136.2000 ;
	    RECT 124.6000 135.8000 125.0000 136.2000 ;
	    RECT 130.2000 136.1000 130.6000 136.2000 ;
	    RECT 131.0000 136.1000 131.4000 136.2000 ;
	    RECT 130.2000 135.8000 131.4000 136.1000 ;
	    RECT 137.4000 135.8000 137.8000 136.2000 ;
	    RECT 140.6000 136.1000 141.0000 136.2000 ;
	    RECT 141.4000 136.1000 141.8000 136.2000 ;
	    RECT 140.6000 135.8000 141.8000 136.1000 ;
	    RECT 115.0000 134.8000 115.4000 135.2000 ;
	    RECT 115.8000 135.1000 116.2000 135.2000 ;
	    RECT 116.6000 135.1000 117.0000 135.2000 ;
	    RECT 115.8000 134.8000 117.0000 135.1000 ;
	    RECT 120.6000 134.8000 121.0000 135.2000 ;
	    RECT 115.0000 134.2000 115.3000 134.8000 ;
	    RECT 115.0000 133.8000 115.4000 134.2000 ;
	    RECT 118.2000 133.8000 118.6000 134.2000 ;
	    RECT 118.2000 133.2000 118.5000 133.8000 ;
	    RECT 115.8000 133.1000 116.2000 133.2000 ;
	    RECT 116.6000 133.1000 117.0000 133.2000 ;
	    RECT 115.8000 132.8000 117.0000 133.1000 ;
	    RECT 117.4000 132.8000 117.8000 133.2000 ;
	    RECT 118.2000 132.8000 118.6000 133.2000 ;
	    RECT 119.8000 132.8000 120.2000 133.2000 ;
	    RECT 121.4000 133.1000 121.8000 133.2000 ;
	    RECT 122.2000 133.1000 122.6000 133.2000 ;
	    RECT 121.4000 132.8000 122.6000 133.1000 ;
	    RECT 116.6000 131.8000 117.0000 132.2000 ;
	    RECT 115.8000 129.8000 116.2000 130.2000 ;
	    RECT 115.8000 129.2000 116.1000 129.8000 ;
	    RECT 115.8000 128.8000 116.2000 129.2000 ;
	    RECT 115.0000 126.8000 115.4000 127.2000 ;
	    RECT 115.0000 124.2000 115.3000 126.8000 ;
	    RECT 116.6000 125.2000 116.9000 131.8000 ;
	    RECT 117.4000 128.2000 117.7000 132.8000 ;
	    RECT 119.8000 132.2000 120.1000 132.8000 ;
	    RECT 119.8000 131.8000 120.2000 132.2000 ;
	    RECT 123.8000 130.2000 124.1000 135.8000 ;
	    RECT 124.6000 135.1000 125.0000 135.2000 ;
	    RECT 125.4000 135.1000 125.8000 135.2000 ;
	    RECT 124.6000 134.8000 125.8000 135.1000 ;
	    RECT 128.6000 134.8000 129.0000 135.2000 ;
	    RECT 132.6000 135.1000 133.0000 135.2000 ;
	    RECT 133.4000 135.1000 133.8000 135.2000 ;
	    RECT 132.6000 134.8000 133.8000 135.1000 ;
	    RECT 134.2000 134.8000 134.6000 135.2000 ;
	    RECT 135.8000 135.1000 136.2000 135.2000 ;
	    RECT 139.0000 135.1000 139.4000 135.2000 ;
	    RECT 135.8000 134.8000 139.4000 135.1000 ;
	    RECT 142.2000 134.8000 142.6000 135.2000 ;
	    RECT 143.8000 135.1000 144.2000 135.2000 ;
	    RECT 143.8000 134.8000 144.9000 135.1000 ;
	    RECT 127.8000 133.8000 128.2000 134.2000 ;
	    RECT 127.0000 131.8000 127.4000 132.2000 ;
	    RECT 124.6000 130.8000 125.0000 131.2000 ;
	    RECT 123.8000 129.8000 124.2000 130.2000 ;
	    RECT 124.6000 129.2000 124.9000 130.8000 ;
	    RECT 118.2000 128.8000 118.6000 129.2000 ;
	    RECT 124.6000 128.8000 125.0000 129.2000 ;
	    RECT 118.2000 128.2000 118.5000 128.8000 ;
	    RECT 117.4000 127.8000 117.8000 128.2000 ;
	    RECT 118.2000 127.8000 118.6000 128.2000 ;
	    RECT 116.6000 124.8000 117.0000 125.2000 ;
	    RECT 115.0000 123.8000 115.4000 124.2000 ;
	    RECT 114.2000 121.8000 114.6000 122.2000 ;
	    RECT 107.0000 114.7000 107.4000 115.1000 ;
	    RECT 107.8000 112.1000 108.2000 117.9000 ;
	    RECT 109.4000 113.1000 109.8000 115.9000 ;
	    RECT 111.8000 113.1000 112.2000 115.9000 ;
	    RECT 113.4000 112.1000 113.8000 117.9000 ;
	    RECT 115.8000 115.1000 116.2000 115.2000 ;
	    RECT 116.6000 115.1000 117.0000 115.2000 ;
	    RECT 115.8000 114.8000 117.0000 115.1000 ;
	    RECT 114.2000 112.8000 114.6000 113.2000 ;
	    RECT 96.6000 105.8000 97.0000 106.2000 ;
	    RECT 99.0000 105.8000 99.4000 106.2000 ;
	    RECT 96.6000 103.2000 96.9000 105.8000 ;
	    RECT 99.0000 105.2000 99.3000 105.8000 ;
	    RECT 99.0000 104.8000 99.4000 105.2000 ;
	    RECT 99.0000 103.8000 99.4000 104.2000 ;
	    RECT 96.6000 102.8000 97.0000 103.2000 ;
	    RECT 91.8000 101.8000 92.2000 102.2000 ;
	    RECT 97.4000 101.8000 97.8000 102.2000 ;
	    RECT 88.6000 99.8000 89.0000 100.2000 ;
	    RECT 91.0000 99.8000 91.4000 100.2000 ;
	    RECT 91.0000 99.2000 91.3000 99.8000 ;
	    RECT 87.0000 98.8000 87.4000 99.2000 ;
	    RECT 87.8000 98.8000 88.2000 99.2000 ;
	    RECT 91.0000 98.8000 91.4000 99.2000 ;
	    RECT 91.8000 97.2000 92.1000 101.8000 ;
	    RECT 97.4000 97.2000 97.7000 101.8000 ;
	    RECT 88.6000 96.8000 89.0000 97.2000 ;
	    RECT 91.0000 96.8000 91.4000 97.2000 ;
	    RECT 91.8000 96.8000 92.2000 97.2000 ;
	    RECT 97.4000 96.8000 97.8000 97.2000 ;
	    RECT 74.2000 95.1000 74.6000 95.2000 ;
	    RECT 75.0000 95.1000 75.4000 95.2000 ;
	    RECT 74.2000 94.8000 75.4000 95.1000 ;
	    RECT 79.8000 94.8000 80.2000 95.2000 ;
	    RECT 81.4000 95.1000 81.8000 95.2000 ;
	    RECT 82.2000 95.1000 82.6000 95.2000 ;
	    RECT 81.4000 94.8000 82.6000 95.1000 ;
	    RECT 86.2000 94.8000 86.6000 95.2000 ;
	    RECT 87.8000 94.8000 88.2000 95.2000 ;
	    RECT 79.8000 94.2000 80.1000 94.8000 ;
	    RECT 79.8000 93.8000 80.2000 94.2000 ;
	    RECT 86.2000 93.8000 86.6000 94.2000 ;
	    RECT 86.2000 93.2000 86.5000 93.8000 ;
	    RECT 75.8000 93.1000 76.2000 93.2000 ;
	    RECT 76.6000 93.1000 77.0000 93.2000 ;
	    RECT 75.8000 92.8000 77.0000 93.1000 ;
	    RECT 83.8000 92.8000 84.2000 93.2000 ;
	    RECT 86.2000 93.1000 86.6000 93.2000 ;
	    RECT 86.2000 92.8000 87.3000 93.1000 ;
	    RECT 75.0000 91.8000 75.4000 92.2000 ;
	    RECT 75.0000 88.2000 75.3000 91.8000 ;
	    RECT 83.8000 88.2000 84.1000 92.8000 ;
	    RECT 86.2000 91.8000 86.6000 92.2000 ;
	    RECT 86.2000 89.2000 86.5000 91.8000 ;
	    RECT 86.2000 88.8000 86.6000 89.2000 ;
	    RECT 75.0000 87.8000 75.4000 88.2000 ;
	    RECT 83.8000 87.8000 84.2000 88.2000 ;
	    RECT 87.0000 87.2000 87.3000 92.8000 ;
	    RECT 87.8000 92.2000 88.1000 94.8000 ;
	    RECT 87.8000 91.8000 88.2000 92.2000 ;
	    RECT 88.6000 89.2000 88.9000 96.8000 ;
	    RECT 91.0000 95.1000 91.3000 96.8000 ;
	    RECT 99.0000 96.2000 99.3000 103.8000 ;
	    RECT 99.8000 103.1000 100.2000 108.9000 ;
	    RECT 100.6000 105.2000 100.9000 111.8000 ;
	    RECT 103.0000 110.8000 103.4000 111.2000 ;
	    RECT 103.0000 109.2000 103.3000 110.8000 ;
	    RECT 102.2000 108.8000 102.6000 109.2000 ;
	    RECT 103.0000 108.8000 103.4000 109.2000 ;
	    RECT 104.6000 108.8000 105.0000 109.2000 ;
	    RECT 111.0000 109.1000 111.4000 109.2000 ;
	    RECT 111.8000 109.1000 112.2000 109.2000 ;
	    RECT 111.0000 108.8000 112.2000 109.1000 ;
	    RECT 102.2000 108.2000 102.5000 108.8000 ;
	    RECT 102.2000 107.8000 102.6000 108.2000 ;
	    RECT 104.6000 107.0000 104.9000 108.8000 ;
	    RECT 106.2000 107.1000 106.6000 107.2000 ;
	    RECT 107.0000 107.1000 107.4000 107.2000 ;
	    RECT 104.6000 106.6000 105.0000 107.0000 ;
	    RECT 106.2000 106.8000 107.4000 107.1000 ;
	    RECT 107.0000 105.8000 107.4000 106.2000 ;
	    RECT 109.4000 106.1000 109.8000 106.2000 ;
	    RECT 110.2000 106.1000 110.6000 106.2000 ;
	    RECT 109.4000 105.8000 110.6000 106.1000 ;
	    RECT 107.0000 105.2000 107.3000 105.8000 ;
	    RECT 100.6000 104.8000 101.0000 105.2000 ;
	    RECT 107.0000 104.8000 107.4000 105.2000 ;
	    RECT 108.6000 102.8000 109.0000 103.2000 ;
	    RECT 113.4000 103.1000 113.8000 108.9000 ;
	    RECT 114.2000 107.2000 114.5000 112.8000 ;
	    RECT 117.4000 109.2000 117.7000 127.8000 ;
	    RECT 127.0000 127.2000 127.3000 131.8000 ;
	    RECT 127.8000 130.2000 128.1000 133.8000 ;
	    RECT 127.8000 129.8000 128.2000 130.2000 ;
	    RECT 127.8000 127.8000 128.2000 128.2000 ;
	    RECT 127.0000 126.8000 127.4000 127.2000 ;
	    RECT 127.8000 126.2000 128.1000 127.8000 ;
	    RECT 119.0000 126.1000 119.4000 126.2000 ;
	    RECT 119.8000 126.1000 120.2000 126.2000 ;
	    RECT 119.0000 125.8000 120.2000 126.1000 ;
	    RECT 120.6000 126.1000 121.0000 126.2000 ;
	    RECT 121.4000 126.1000 121.8000 126.2000 ;
	    RECT 120.6000 125.8000 121.8000 126.1000 ;
	    RECT 126.2000 125.8000 126.6000 126.2000 ;
	    RECT 127.8000 125.8000 128.2000 126.2000 ;
	    RECT 121.4000 124.8000 121.8000 125.2000 ;
	    RECT 123.8000 125.1000 124.2000 125.2000 ;
	    RECT 124.6000 125.1000 125.0000 125.2000 ;
	    RECT 123.8000 124.8000 125.0000 125.1000 ;
	    RECT 121.4000 124.2000 121.7000 124.8000 ;
	    RECT 120.6000 123.8000 121.0000 124.2000 ;
	    RECT 121.4000 123.8000 121.8000 124.2000 ;
	    RECT 120.6000 119.2000 120.9000 123.8000 ;
	    RECT 120.6000 118.8000 121.0000 119.2000 ;
	    RECT 118.2000 112.1000 118.6000 117.9000 ;
	    RECT 121.4000 116.2000 121.7000 123.8000 ;
	    RECT 126.2000 123.2000 126.5000 125.8000 ;
	    RECT 126.2000 122.8000 126.6000 123.2000 ;
	    RECT 128.6000 122.2000 128.9000 134.8000 ;
	    RECT 130.2000 133.8000 130.6000 134.2000 ;
	    RECT 129.4000 130.8000 129.8000 131.2000 ;
	    RECT 130.2000 131.1000 130.5000 133.8000 ;
	    RECT 131.0000 133.1000 131.4000 133.2000 ;
	    RECT 131.0000 132.8000 132.1000 133.1000 ;
	    RECT 131.0000 131.1000 131.4000 131.2000 ;
	    RECT 130.2000 130.8000 131.4000 131.1000 ;
	    RECT 129.4000 130.1000 129.7000 130.8000 ;
	    RECT 129.4000 129.8000 130.5000 130.1000 ;
	    RECT 129.4000 128.8000 129.8000 129.2000 ;
	    RECT 129.4000 128.2000 129.7000 128.8000 ;
	    RECT 130.2000 128.2000 130.5000 129.8000 ;
	    RECT 131.0000 128.2000 131.3000 130.8000 ;
	    RECT 131.8000 128.2000 132.1000 132.8000 ;
	    RECT 129.4000 127.8000 129.8000 128.2000 ;
	    RECT 130.2000 127.8000 130.6000 128.2000 ;
	    RECT 131.0000 127.8000 131.4000 128.2000 ;
	    RECT 131.8000 127.8000 132.2000 128.2000 ;
	    RECT 132.6000 127.2000 132.9000 134.8000 ;
	    RECT 133.4000 133.8000 133.8000 134.2000 ;
	    RECT 133.4000 133.2000 133.7000 133.8000 ;
	    RECT 133.4000 132.8000 133.8000 133.2000 ;
	    RECT 134.2000 132.2000 134.5000 134.8000 ;
	    RECT 136.6000 134.1000 137.0000 134.2000 ;
	    RECT 137.4000 134.1000 137.8000 134.2000 ;
	    RECT 136.6000 133.8000 137.8000 134.1000 ;
	    RECT 139.8000 134.1000 140.2000 134.2000 ;
	    RECT 140.6000 134.1000 141.0000 134.2000 ;
	    RECT 139.8000 133.8000 141.0000 134.1000 ;
	    RECT 142.2000 132.2000 142.5000 134.8000 ;
	    RECT 143.0000 133.8000 143.4000 134.2000 ;
	    RECT 143.8000 133.8000 144.2000 134.2000 ;
	    RECT 134.2000 131.8000 134.6000 132.2000 ;
	    RECT 142.2000 131.8000 142.6000 132.2000 ;
	    RECT 143.0000 130.2000 143.3000 133.8000 ;
	    RECT 143.8000 133.2000 144.1000 133.8000 ;
	    RECT 143.8000 132.8000 144.2000 133.2000 ;
	    RECT 143.0000 129.8000 143.4000 130.2000 ;
	    RECT 138.2000 128.8000 138.6000 129.2000 ;
	    RECT 141.4000 128.8000 141.8000 129.2000 ;
	    RECT 135.8000 128.1000 136.2000 128.2000 ;
	    RECT 136.6000 128.1000 137.0000 128.2000 ;
	    RECT 135.8000 127.8000 137.0000 128.1000 ;
	    RECT 137.4000 127.8000 137.8000 128.2000 ;
	    RECT 131.0000 126.8000 131.4000 127.2000 ;
	    RECT 132.6000 126.8000 133.0000 127.2000 ;
	    RECT 135.8000 126.8000 136.2000 127.2000 ;
	    RECT 131.0000 126.2000 131.3000 126.8000 ;
	    RECT 135.8000 126.2000 136.1000 126.8000 ;
	    RECT 131.0000 125.8000 131.4000 126.2000 ;
	    RECT 134.2000 126.1000 134.6000 126.2000 ;
	    RECT 135.0000 126.1000 135.4000 126.2000 ;
	    RECT 134.2000 125.8000 135.4000 126.1000 ;
	    RECT 135.8000 125.8000 136.2000 126.2000 ;
	    RECT 134.2000 122.8000 134.6000 123.2000 ;
	    RECT 122.2000 121.8000 122.6000 122.2000 ;
	    RECT 124.6000 121.8000 125.0000 122.2000 ;
	    RECT 128.6000 121.8000 129.0000 122.2000 ;
	    RECT 121.4000 115.8000 121.8000 116.2000 ;
	    RECT 122.2000 115.2000 122.5000 121.8000 ;
	    RECT 123.8000 115.8000 124.2000 116.2000 ;
	    RECT 123.8000 115.2000 124.1000 115.8000 ;
	    RECT 124.6000 115.2000 124.9000 121.8000 ;
	    RECT 127.8000 115.8000 128.2000 116.2000 ;
	    RECT 130.2000 115.8000 130.6000 116.2000 ;
	    RECT 127.8000 115.2000 128.1000 115.8000 ;
	    RECT 130.2000 115.2000 130.5000 115.8000 ;
	    RECT 120.6000 114.8000 121.0000 115.2000 ;
	    RECT 122.2000 114.8000 122.6000 115.2000 ;
	    RECT 123.8000 114.8000 124.2000 115.2000 ;
	    RECT 124.6000 114.8000 125.0000 115.2000 ;
	    RECT 127.8000 114.8000 128.2000 115.2000 ;
	    RECT 129.4000 114.8000 129.8000 115.2000 ;
	    RECT 130.2000 114.8000 130.6000 115.2000 ;
	    RECT 132.6000 115.1000 133.0000 115.2000 ;
	    RECT 133.4000 115.1000 133.8000 115.2000 ;
	    RECT 132.6000 114.8000 133.8000 115.1000 ;
	    RECT 120.6000 109.2000 120.9000 114.8000 ;
	    RECT 123.8000 113.8000 124.2000 114.2000 ;
	    RECT 123.8000 112.2000 124.1000 113.8000 ;
	    RECT 123.8000 111.8000 124.2000 112.2000 ;
	    RECT 117.4000 108.8000 117.8000 109.2000 ;
	    RECT 114.2000 106.8000 114.6000 107.2000 ;
	    RECT 116.6000 105.8000 117.0000 106.2000 ;
	    RECT 116.6000 105.2000 116.9000 105.8000 ;
	    RECT 116.6000 104.8000 117.0000 105.2000 ;
	    RECT 118.2000 103.1000 118.6000 108.9000 ;
	    RECT 120.6000 108.8000 121.0000 109.2000 ;
	    RECT 119.0000 106.8000 119.4000 107.2000 ;
	    RECT 119.0000 105.2000 119.3000 106.8000 ;
	    RECT 119.0000 104.8000 119.4000 105.2000 ;
	    RECT 119.8000 105.1000 120.2000 107.9000 ;
	    RECT 123.0000 106.8000 123.4000 107.2000 ;
	    RECT 123.8000 106.8000 124.2000 107.2000 ;
	    RECT 122.2000 105.8000 122.6000 106.2000 ;
	    RECT 108.6000 99.2000 108.9000 102.8000 ;
	    RECT 114.2000 100.8000 114.6000 101.2000 ;
	    RECT 108.6000 98.8000 109.0000 99.2000 ;
	    RECT 109.4000 98.8000 109.8000 99.2000 ;
	    RECT 106.2000 96.8000 106.6000 97.2000 ;
	    RECT 99.0000 95.8000 99.4000 96.2000 ;
	    RECT 99.8000 95.8000 100.2000 96.2000 ;
	    RECT 90.2000 94.8000 91.3000 95.1000 ;
	    RECT 91.8000 95.1000 92.2000 95.2000 ;
	    RECT 95.8000 95.1000 96.2000 95.2000 ;
	    RECT 91.8000 94.8000 96.2000 95.1000 ;
	    RECT 97.4000 95.1000 97.8000 95.2000 ;
	    RECT 98.2000 95.1000 98.6000 95.2000 ;
	    RECT 97.4000 94.8000 98.6000 95.1000 ;
	    RECT 90.2000 89.2000 90.5000 94.8000 ;
	    RECT 91.0000 92.8000 91.4000 93.2000 ;
	    RECT 92.6000 93.1000 93.0000 93.2000 ;
	    RECT 93.4000 93.1000 93.8000 93.2000 ;
	    RECT 92.6000 92.8000 93.8000 93.1000 ;
	    RECT 88.6000 88.8000 89.0000 89.2000 ;
	    RECT 90.2000 88.8000 90.6000 89.2000 ;
	    RECT 91.0000 87.2000 91.3000 92.8000 ;
	    RECT 99.0000 92.2000 99.3000 95.8000 ;
	    RECT 99.8000 95.2000 100.1000 95.8000 ;
	    RECT 106.2000 95.2000 106.5000 96.8000 ;
	    RECT 109.4000 95.2000 109.7000 98.8000 ;
	    RECT 114.2000 95.2000 114.5000 100.8000 ;
	    RECT 122.2000 100.2000 122.5000 105.8000 ;
	    RECT 122.2000 99.8000 122.6000 100.2000 ;
	    RECT 99.8000 94.8000 100.2000 95.2000 ;
	    RECT 102.2000 94.8000 102.6000 95.2000 ;
	    RECT 105.4000 94.8000 105.8000 95.2000 ;
	    RECT 106.2000 94.8000 106.6000 95.2000 ;
	    RECT 109.4000 94.8000 109.8000 95.2000 ;
	    RECT 114.2000 94.8000 114.6000 95.2000 ;
	    RECT 102.2000 94.2000 102.5000 94.8000 ;
	    RECT 105.4000 94.2000 105.7000 94.8000 ;
	    RECT 100.6000 93.8000 101.0000 94.2000 ;
	    RECT 102.2000 93.8000 102.6000 94.2000 ;
	    RECT 104.6000 93.8000 105.0000 94.2000 ;
	    RECT 105.4000 93.8000 105.8000 94.2000 ;
	    RECT 107.0000 93.8000 107.4000 94.2000 ;
	    RECT 109.4000 94.1000 109.8000 94.2000 ;
	    RECT 110.2000 94.1000 110.6000 94.2000 ;
	    RECT 109.4000 93.8000 110.6000 94.1000 ;
	    RECT 115.0000 93.8000 115.4000 94.2000 ;
	    RECT 115.8000 94.1000 116.2000 94.2000 ;
	    RECT 116.6000 94.1000 117.0000 94.2000 ;
	    RECT 115.8000 93.8000 117.0000 94.1000 ;
	    RECT 98.2000 91.8000 98.6000 92.2000 ;
	    RECT 99.0000 91.8000 99.4000 92.2000 ;
	    RECT 93.4000 87.8000 93.8000 88.2000 ;
	    RECT 75.0000 86.8000 75.4000 87.2000 ;
	    RECT 75.8000 86.8000 76.2000 87.2000 ;
	    RECT 82.2000 87.1000 82.6000 87.2000 ;
	    RECT 83.0000 87.1000 83.4000 87.2000 ;
	    RECT 82.2000 86.8000 83.4000 87.1000 ;
	    RECT 87.0000 86.8000 87.4000 87.2000 ;
	    RECT 91.0000 86.8000 91.4000 87.2000 ;
	    RECT 74.2000 86.1000 74.6000 86.2000 ;
	    RECT 75.0000 86.1000 75.3000 86.8000 ;
	    RECT 74.2000 85.8000 75.3000 86.1000 ;
	    RECT 75.8000 86.2000 76.1000 86.8000 ;
	    RECT 93.4000 86.2000 93.7000 87.8000 ;
	    RECT 75.8000 85.8000 76.2000 86.2000 ;
	    RECT 76.6000 85.8000 77.0000 86.2000 ;
	    RECT 78.2000 86.1000 78.6000 86.2000 ;
	    RECT 79.0000 86.1000 79.4000 86.2000 ;
	    RECT 78.2000 85.8000 79.4000 86.1000 ;
	    RECT 81.4000 85.8000 81.8000 86.2000 ;
	    RECT 83.0000 85.8000 83.4000 86.2000 ;
	    RECT 93.4000 85.8000 93.8000 86.2000 ;
	    RECT 95.8000 86.1000 96.2000 86.2000 ;
	    RECT 96.6000 86.1000 97.0000 86.2000 ;
	    RECT 95.8000 85.8000 97.0000 86.1000 ;
	    RECT 76.6000 85.2000 76.9000 85.8000 ;
	    RECT 81.4000 85.2000 81.7000 85.8000 ;
	    RECT 39.8000 84.8000 40.2000 85.2000 ;
	    RECT 43.8000 84.8000 44.2000 85.2000 ;
	    RECT 44.6000 84.8000 45.0000 85.2000 ;
	    RECT 48.6000 84.8000 49.0000 85.2000 ;
	    RECT 49.4000 85.1000 49.8000 85.2000 ;
	    RECT 50.2000 85.1000 50.6000 85.2000 ;
	    RECT 49.4000 84.8000 50.6000 85.1000 ;
	    RECT 51.0000 84.8000 51.4000 85.2000 ;
	    RECT 56.6000 85.1000 57.0000 85.2000 ;
	    RECT 57.4000 85.1000 57.8000 85.2000 ;
	    RECT 56.6000 84.8000 57.8000 85.1000 ;
	    RECT 67.8000 84.8000 68.2000 85.2000 ;
	    RECT 68.6000 84.8000 69.0000 85.2000 ;
	    RECT 73.4000 84.8000 73.8000 85.2000 ;
	    RECT 76.6000 84.8000 77.0000 85.2000 ;
	    RECT 79.0000 85.1000 79.4000 85.2000 ;
	    RECT 79.8000 85.1000 80.2000 85.2000 ;
	    RECT 79.0000 84.8000 80.2000 85.1000 ;
	    RECT 81.4000 84.8000 81.8000 85.2000 ;
	    RECT 39.8000 82.2000 40.1000 84.8000 ;
	    RECT 42.2000 83.8000 42.6000 84.2000 ;
	    RECT 37.4000 81.8000 37.8000 82.2000 ;
	    RECT 39.0000 81.8000 39.4000 82.2000 ;
	    RECT 39.8000 81.8000 40.2000 82.2000 ;
	    RECT 37.4000 79.2000 37.7000 81.8000 ;
	    RECT 39.0000 81.2000 39.3000 81.8000 ;
	    RECT 42.2000 81.2000 42.5000 83.8000 ;
	    RECT 39.0000 80.8000 39.4000 81.2000 ;
	    RECT 42.2000 80.8000 42.6000 81.2000 ;
	    RECT 43.8000 80.2000 44.1000 84.8000 ;
	    RECT 48.6000 84.1000 49.0000 84.2000 ;
	    RECT 49.4000 84.1000 49.8000 84.2000 ;
	    RECT 48.6000 83.8000 49.8000 84.1000 ;
	    RECT 46.2000 81.8000 46.6000 82.2000 ;
	    RECT 50.2000 81.8000 50.6000 82.2000 ;
	    RECT 46.2000 80.2000 46.5000 81.8000 ;
	    RECT 39.8000 79.8000 40.2000 80.2000 ;
	    RECT 43.8000 79.8000 44.2000 80.2000 ;
	    RECT 46.2000 79.8000 46.6000 80.2000 ;
	    RECT 39.8000 79.2000 40.1000 79.8000 ;
	    RECT 50.2000 79.2000 50.5000 81.8000 ;
	    RECT 37.4000 78.8000 37.8000 79.2000 ;
	    RECT 39.8000 78.8000 40.2000 79.2000 ;
	    RECT 50.2000 78.8000 50.6000 79.2000 ;
	    RECT 44.6000 76.8000 45.0000 77.2000 ;
	    RECT 48.6000 77.1000 49.0000 77.2000 ;
	    RECT 49.4000 77.1000 49.8000 77.2000 ;
	    RECT 48.6000 76.8000 49.8000 77.1000 ;
	    RECT 44.6000 76.2000 44.9000 76.8000 ;
	    RECT 51.0000 76.2000 51.3000 84.8000 ;
	    RECT 67.8000 84.2000 68.1000 84.8000 ;
	    RECT 55.0000 84.1000 55.4000 84.2000 ;
	    RECT 55.8000 84.1000 56.2000 84.2000 ;
	    RECT 55.0000 83.8000 56.2000 84.1000 ;
	    RECT 62.2000 84.1000 62.6000 84.2000 ;
	    RECT 63.0000 84.1000 63.4000 84.2000 ;
	    RECT 62.2000 83.8000 63.4000 84.1000 ;
	    RECT 67.8000 83.8000 68.2000 84.2000 ;
	    RECT 67.0000 82.8000 67.4000 83.2000 ;
	    RECT 67.0000 82.2000 67.3000 82.8000 ;
	    RECT 68.6000 82.2000 68.9000 84.8000 ;
	    RECT 71.8000 83.8000 72.2000 84.2000 ;
	    RECT 72.6000 83.8000 73.0000 84.2000 ;
	    RECT 71.8000 83.2000 72.1000 83.8000 ;
	    RECT 71.8000 82.8000 72.2000 83.2000 ;
	    RECT 55.8000 81.8000 56.2000 82.2000 ;
	    RECT 67.0000 81.8000 67.4000 82.2000 ;
	    RECT 68.6000 81.8000 69.0000 82.2000 ;
	    RECT 69.4000 81.8000 69.8000 82.2000 ;
	    RECT 55.8000 77.2000 56.1000 81.8000 ;
	    RECT 69.4000 79.2000 69.7000 81.8000 ;
	    RECT 72.6000 79.2000 72.9000 83.8000 ;
	    RECT 73.4000 79.2000 73.7000 84.8000 ;
	    RECT 75.0000 83.8000 75.4000 84.2000 ;
	    RECT 78.2000 83.8000 78.6000 84.2000 ;
	    RECT 81.4000 83.8000 81.8000 84.2000 ;
	    RECT 75.0000 80.2000 75.3000 83.8000 ;
	    RECT 78.2000 83.2000 78.5000 83.8000 ;
	    RECT 78.2000 82.8000 78.6000 83.2000 ;
	    RECT 79.0000 81.8000 79.4000 82.2000 ;
	    RECT 75.0000 79.8000 75.4000 80.2000 ;
	    RECT 59.0000 79.1000 59.4000 79.2000 ;
	    RECT 59.8000 79.1000 60.2000 79.2000 ;
	    RECT 59.0000 78.8000 60.2000 79.1000 ;
	    RECT 63.8000 79.1000 64.2000 79.2000 ;
	    RECT 64.6000 79.1000 65.0000 79.2000 ;
	    RECT 63.8000 78.8000 65.0000 79.1000 ;
	    RECT 69.4000 78.8000 69.8000 79.2000 ;
	    RECT 70.2000 78.8000 70.6000 79.2000 ;
	    RECT 72.6000 78.8000 73.0000 79.2000 ;
	    RECT 73.4000 78.8000 73.8000 79.2000 ;
	    RECT 55.8000 76.8000 56.2000 77.2000 ;
	    RECT 58.2000 76.8000 58.6000 77.2000 ;
	    RECT 63.0000 76.8000 63.4000 77.2000 ;
	    RECT 63.8000 76.8000 64.2000 77.2000 ;
	    RECT 67.8000 76.8000 68.2000 77.2000 ;
	    RECT 68.6000 76.8000 69.0000 77.2000 ;
	    RECT 39.0000 75.8000 39.4000 76.2000 ;
	    RECT 44.6000 75.8000 45.0000 76.2000 ;
	    RECT 47.8000 75.8000 48.2000 76.2000 ;
	    RECT 51.0000 75.8000 51.4000 76.2000 ;
	    RECT 54.2000 76.1000 54.6000 76.2000 ;
	    RECT 55.0000 76.1000 55.4000 76.2000 ;
	    RECT 54.2000 75.8000 55.4000 76.1000 ;
	    RECT 16.6000 74.8000 17.0000 75.2000 ;
	    RECT 27.8000 74.8000 28.2000 75.2000 ;
	    RECT 29.4000 74.8000 29.8000 75.2000 ;
	    RECT 35.8000 74.8000 36.2000 75.2000 ;
	    RECT 37.4000 74.8000 37.8000 75.2000 ;
	    RECT 12.6000 71.8000 13.0000 72.2000 ;
	    RECT 15.0000 71.8000 15.4000 72.2000 ;
	    RECT 10.2000 70.8000 10.6000 71.2000 ;
	    RECT 5.4000 67.8000 5.8000 68.2000 ;
	    RECT 7.8000 67.8000 8.2000 68.2000 ;
	    RECT 11.0000 67.8000 11.4000 68.2000 ;
	    RECT 7.8000 67.1000 8.2000 67.2000 ;
	    RECT 8.6000 67.1000 9.0000 67.2000 ;
	    RECT 7.8000 66.8000 9.0000 67.1000 ;
	    RECT 9.4000 66.8000 9.8000 67.2000 ;
	    RECT 10.2000 66.8000 10.6000 67.2000 ;
	    RECT 2.2000 65.8000 3.3000 66.1000 ;
	    RECT 9.4000 66.2000 9.7000 66.8000 ;
	    RECT 9.4000 65.8000 9.8000 66.2000 ;
	    RECT 3.0000 65.1000 3.4000 65.2000 ;
	    RECT 3.8000 65.1000 4.2000 65.2000 ;
	    RECT 3.0000 64.8000 4.2000 65.1000 ;
	    RECT 8.6000 65.1000 9.0000 65.2000 ;
	    RECT 9.4000 65.1000 9.8000 65.2000 ;
	    RECT 8.6000 64.8000 9.8000 65.1000 ;
	    RECT 10.2000 64.2000 10.5000 66.8000 ;
	    RECT 1.4000 63.8000 1.8000 64.2000 ;
	    RECT 10.2000 63.8000 10.6000 64.2000 ;
	    RECT 2.2000 61.8000 2.6000 62.2000 ;
	    RECT 3.0000 61.8000 3.4000 62.2000 ;
	    RECT 3.8000 62.1000 4.2000 62.2000 ;
	    RECT 4.6000 62.1000 5.0000 62.2000 ;
	    RECT 3.8000 61.8000 5.0000 62.1000 ;
	    RECT 1.4000 56.8000 1.8000 57.2000 ;
	    RECT 1.4000 49.2000 1.7000 56.8000 ;
	    RECT 2.2000 55.2000 2.5000 61.8000 ;
	    RECT 3.0000 56.2000 3.3000 61.8000 ;
	    RECT 5.4000 57.8000 5.8000 58.2000 ;
	    RECT 6.2000 57.8000 6.6000 58.2000 ;
	    RECT 7.8000 58.1000 8.2000 58.2000 ;
	    RECT 8.6000 58.1000 9.0000 58.2000 ;
	    RECT 7.8000 57.8000 9.0000 58.1000 ;
	    RECT 5.4000 57.2000 5.7000 57.8000 ;
	    RECT 3.8000 57.1000 4.2000 57.2000 ;
	    RECT 4.6000 57.1000 5.0000 57.2000 ;
	    RECT 3.8000 56.8000 5.0000 57.1000 ;
	    RECT 5.4000 56.8000 5.8000 57.2000 ;
	    RECT 6.2000 56.2000 6.5000 57.8000 ;
	    RECT 3.0000 55.8000 3.4000 56.2000 ;
	    RECT 6.2000 55.8000 6.6000 56.2000 ;
	    RECT 3.0000 55.2000 3.3000 55.8000 ;
	    RECT 11.0000 55.2000 11.3000 67.8000 ;
	    RECT 12.6000 67.2000 12.9000 71.8000 ;
	    RECT 13.4000 67.8000 13.8000 68.2000 ;
	    RECT 12.6000 66.8000 13.0000 67.2000 ;
	    RECT 13.4000 65.1000 13.7000 67.8000 ;
	    RECT 16.6000 66.2000 16.9000 74.8000 ;
	    RECT 29.4000 74.2000 29.7000 74.8000 ;
	    RECT 17.4000 74.1000 17.8000 74.2000 ;
	    RECT 18.2000 74.1000 18.6000 74.2000 ;
	    RECT 17.4000 73.8000 18.6000 74.1000 ;
	    RECT 22.2000 74.1000 22.6000 74.2000 ;
	    RECT 23.0000 74.1000 23.4000 74.2000 ;
	    RECT 22.2000 73.8000 23.4000 74.1000 ;
	    RECT 29.4000 73.8000 29.8000 74.2000 ;
	    RECT 31.8000 73.8000 32.2000 74.2000 ;
	    RECT 17.4000 71.8000 17.8000 72.2000 ;
	    RECT 19.0000 71.8000 19.4000 72.2000 ;
	    RECT 17.4000 66.2000 17.7000 71.8000 ;
	    RECT 12.6000 64.8000 13.7000 65.1000 ;
	    RECT 15.8000 65.8000 16.2000 66.2000 ;
	    RECT 16.6000 65.8000 17.0000 66.2000 ;
	    RECT 17.4000 65.8000 17.8000 66.2000 ;
	    RECT 11.8000 60.8000 12.2000 61.2000 ;
	    RECT 2.2000 54.8000 2.6000 55.2000 ;
	    RECT 3.0000 54.8000 3.4000 55.2000 ;
	    RECT 5.4000 54.8000 5.8000 55.2000 ;
	    RECT 11.0000 55.1000 11.4000 55.2000 ;
	    RECT 10.2000 54.8000 11.4000 55.1000 ;
	    RECT 5.4000 54.2000 5.7000 54.8000 ;
	    RECT 2.2000 53.8000 2.6000 54.2000 ;
	    RECT 5.4000 53.8000 5.8000 54.2000 ;
	    RECT 2.2000 53.2000 2.5000 53.8000 ;
	    RECT 2.2000 52.8000 2.6000 53.2000 ;
	    RECT 9.4000 49.8000 9.8000 50.2000 ;
	    RECT 1.4000 48.8000 1.8000 49.2000 ;
	    RECT 6.2000 48.1000 6.6000 48.2000 ;
	    RECT 7.0000 48.1000 7.4000 48.2000 ;
	    RECT 6.2000 47.8000 7.4000 48.1000 ;
	    RECT 3.8000 46.8000 4.2000 47.2000 ;
	    RECT 3.8000 46.2000 4.1000 46.8000 ;
	    RECT 1.4000 46.1000 1.8000 46.2000 ;
	    RECT 2.2000 46.1000 2.6000 46.2000 ;
	    RECT 1.4000 45.8000 2.6000 46.1000 ;
	    RECT 3.8000 45.8000 4.2000 46.2000 ;
	    RECT 7.8000 45.8000 8.2000 46.2000 ;
	    RECT 7.8000 44.2000 8.1000 45.8000 ;
	    RECT 2.2000 44.1000 2.6000 44.2000 ;
	    RECT 3.0000 44.1000 3.4000 44.2000 ;
	    RECT 2.2000 43.8000 3.4000 44.1000 ;
	    RECT 7.8000 43.8000 8.2000 44.2000 ;
	    RECT 4.6000 41.8000 5.0000 42.2000 ;
	    RECT 4.6000 37.2000 4.9000 41.8000 ;
	    RECT 9.4000 39.2000 9.7000 49.8000 ;
	    RECT 10.2000 48.2000 10.5000 54.8000 ;
	    RECT 11.8000 49.2000 12.1000 60.8000 ;
	    RECT 12.6000 56.2000 12.9000 64.8000 ;
	    RECT 15.8000 64.2000 16.1000 65.8000 ;
	    RECT 17.4000 64.8000 17.8000 65.2000 ;
	    RECT 13.4000 63.8000 13.8000 64.2000 ;
	    RECT 15.8000 63.8000 16.2000 64.2000 ;
	    RECT 13.4000 61.2000 13.7000 63.8000 ;
	    RECT 14.2000 61.8000 14.6000 62.2000 ;
	    RECT 16.6000 61.8000 17.0000 62.2000 ;
	    RECT 13.4000 60.8000 13.8000 61.2000 ;
	    RECT 14.2000 57.2000 14.5000 61.8000 ;
	    RECT 15.0000 57.8000 15.4000 58.2000 ;
	    RECT 15.8000 57.8000 16.2000 58.2000 ;
	    RECT 15.0000 57.2000 15.3000 57.8000 ;
	    RECT 14.2000 56.8000 14.6000 57.2000 ;
	    RECT 15.0000 56.8000 15.4000 57.2000 ;
	    RECT 15.8000 56.2000 16.1000 57.8000 ;
	    RECT 16.6000 57.2000 16.9000 61.8000 ;
	    RECT 17.4000 58.2000 17.7000 64.8000 ;
	    RECT 19.0000 64.2000 19.3000 71.8000 ;
	    RECT 23.0000 68.2000 23.3000 73.8000 ;
	    RECT 31.8000 73.2000 32.1000 73.8000 ;
	    RECT 31.8000 72.8000 32.2000 73.2000 ;
	    RECT 33.4000 72.8000 33.8000 73.2000 ;
	    RECT 23.8000 72.1000 24.2000 72.2000 ;
	    RECT 23.8000 71.8000 24.9000 72.1000 ;
	    RECT 21.4000 67.8000 21.8000 68.2000 ;
	    RECT 23.0000 67.8000 23.4000 68.2000 ;
	    RECT 21.4000 67.2000 21.7000 67.8000 ;
	    RECT 23.0000 67.2000 23.3000 67.8000 ;
	    RECT 19.8000 66.8000 20.2000 67.2000 ;
	    RECT 21.4000 66.8000 21.8000 67.2000 ;
	    RECT 23.0000 66.8000 23.4000 67.2000 ;
	    RECT 19.8000 66.2000 20.1000 66.8000 ;
	    RECT 19.8000 65.8000 20.2000 66.2000 ;
	    RECT 24.6000 65.2000 24.9000 71.8000 ;
	    RECT 30.2000 71.8000 30.6000 72.2000 ;
	    RECT 30.2000 71.2000 30.5000 71.8000 ;
	    RECT 25.4000 70.8000 25.8000 71.2000 ;
	    RECT 30.2000 70.8000 30.6000 71.2000 ;
	    RECT 25.4000 66.2000 25.7000 70.8000 ;
	    RECT 26.2000 68.1000 26.6000 68.2000 ;
	    RECT 27.0000 68.1000 27.4000 68.2000 ;
	    RECT 26.2000 67.8000 27.4000 68.1000 ;
	    RECT 33.4000 67.2000 33.7000 72.8000 ;
	    RECT 37.4000 67.2000 37.7000 74.8000 ;
	    RECT 39.0000 69.2000 39.3000 75.8000 ;
	    RECT 47.8000 75.2000 48.1000 75.8000 ;
	    RECT 47.8000 74.8000 48.2000 75.2000 ;
	    RECT 49.4000 75.1000 49.8000 75.2000 ;
	    RECT 50.2000 75.1000 50.6000 75.2000 ;
	    RECT 49.4000 74.8000 50.6000 75.1000 ;
	    RECT 46.2000 73.8000 46.6000 74.2000 ;
	    RECT 58.2000 74.1000 58.5000 76.8000 ;
	    RECT 59.0000 75.8000 59.4000 76.2000 ;
	    RECT 59.0000 75.2000 59.3000 75.8000 ;
	    RECT 59.0000 74.8000 59.4000 75.2000 ;
	    RECT 57.4000 73.8000 58.5000 74.1000 ;
	    RECT 46.2000 73.2000 46.5000 73.8000 ;
	    RECT 46.2000 72.8000 46.6000 73.2000 ;
	    RECT 48.6000 72.8000 49.0000 73.2000 ;
	    RECT 51.8000 73.1000 52.2000 73.2000 ;
	    RECT 52.6000 73.1000 53.0000 73.2000 ;
	    RECT 51.8000 72.8000 53.0000 73.1000 ;
	    RECT 55.0000 72.8000 55.4000 73.2000 ;
	    RECT 46.2000 70.8000 46.6000 71.2000 ;
	    RECT 46.2000 69.2000 46.5000 70.8000 ;
	    RECT 39.0000 68.8000 39.4000 69.2000 ;
	    RECT 46.2000 68.8000 46.6000 69.2000 ;
	    RECT 48.6000 67.2000 48.9000 72.8000 ;
	    RECT 29.4000 66.8000 29.8000 67.2000 ;
	    RECT 33.4000 66.8000 33.8000 67.2000 ;
	    RECT 37.4000 66.8000 37.8000 67.2000 ;
	    RECT 41.4000 67.1000 41.8000 67.2000 ;
	    RECT 42.2000 67.1000 42.6000 67.2000 ;
	    RECT 41.4000 66.8000 42.6000 67.1000 ;
	    RECT 44.6000 66.8000 45.0000 67.2000 ;
	    RECT 48.6000 66.8000 49.0000 67.2000 ;
	    RECT 49.4000 67.1000 49.8000 67.2000 ;
	    RECT 50.2000 67.1000 50.6000 67.2000 ;
	    RECT 49.4000 66.8000 50.6000 67.1000 ;
	    RECT 29.4000 66.2000 29.7000 66.8000 ;
	    RECT 25.4000 65.8000 25.8000 66.2000 ;
	    RECT 29.4000 65.8000 29.8000 66.2000 ;
	    RECT 30.2000 66.1000 30.6000 66.2000 ;
	    RECT 31.0000 66.1000 31.4000 66.2000 ;
	    RECT 30.2000 65.8000 31.4000 66.1000 ;
	    RECT 24.6000 64.8000 25.0000 65.2000 ;
	    RECT 25.4000 65.1000 25.8000 65.2000 ;
	    RECT 26.2000 65.1000 26.6000 65.2000 ;
	    RECT 25.4000 64.8000 26.6000 65.1000 ;
	    RECT 29.4000 65.1000 29.8000 65.2000 ;
	    RECT 30.2000 65.1000 30.6000 65.2000 ;
	    RECT 29.4000 64.8000 30.6000 65.1000 ;
	    RECT 31.8000 64.8000 32.2000 65.2000 ;
	    RECT 31.8000 64.2000 32.1000 64.8000 ;
	    RECT 19.0000 63.8000 19.4000 64.2000 ;
	    RECT 31.0000 63.8000 31.4000 64.2000 ;
	    RECT 31.8000 63.8000 32.2000 64.2000 ;
	    RECT 31.0000 63.2000 31.3000 63.8000 ;
	    RECT 33.4000 63.2000 33.7000 66.8000 ;
	    RECT 44.6000 66.2000 44.9000 66.8000 ;
	    RECT 52.6000 66.2000 52.9000 72.8000 ;
	    RECT 55.0000 72.2000 55.3000 72.8000 ;
	    RECT 55.0000 72.1000 55.4000 72.2000 ;
	    RECT 55.0000 71.8000 56.1000 72.1000 ;
	    RECT 55.8000 67.2000 56.1000 71.8000 ;
	    RECT 57.4000 69.2000 57.7000 73.8000 ;
	    RECT 63.0000 73.2000 63.3000 76.8000 ;
	    RECT 63.8000 75.2000 64.1000 76.8000 ;
	    RECT 63.8000 74.8000 64.2000 75.2000 ;
	    RECT 59.0000 72.8000 59.4000 73.2000 ;
	    RECT 63.0000 72.8000 63.4000 73.2000 ;
	    RECT 64.6000 72.8000 65.0000 73.2000 ;
	    RECT 59.0000 69.2000 59.3000 72.8000 ;
	    RECT 64.6000 69.2000 64.9000 72.8000 ;
	    RECT 67.0000 71.8000 67.4000 72.2000 ;
	    RECT 57.4000 68.8000 57.8000 69.2000 ;
	    RECT 59.0000 68.8000 59.4000 69.2000 ;
	    RECT 64.6000 68.8000 65.0000 69.2000 ;
	    RECT 67.0000 68.2000 67.3000 71.8000 ;
	    RECT 67.8000 69.2000 68.1000 76.8000 ;
	    RECT 68.6000 73.2000 68.9000 76.8000 ;
	    RECT 70.2000 76.2000 70.5000 78.8000 ;
	    RECT 71.8000 77.1000 72.2000 77.2000 ;
	    RECT 72.6000 77.1000 73.0000 77.2000 ;
	    RECT 71.8000 76.8000 73.0000 77.1000 ;
	    RECT 70.2000 75.8000 70.6000 76.2000 ;
	    RECT 79.0000 75.2000 79.3000 81.8000 ;
	    RECT 81.4000 79.2000 81.7000 83.8000 ;
	    RECT 81.4000 78.8000 81.8000 79.2000 ;
	    RECT 82.2000 76.8000 82.6000 77.2000 ;
	    RECT 69.4000 75.1000 69.8000 75.2000 ;
	    RECT 72.6000 75.1000 73.0000 75.2000 ;
	    RECT 73.4000 75.1000 73.8000 75.2000 ;
	    RECT 69.4000 74.8000 70.5000 75.1000 ;
	    RECT 72.6000 74.8000 73.8000 75.1000 ;
	    RECT 74.2000 75.1000 74.6000 75.2000 ;
	    RECT 75.0000 75.1000 75.4000 75.2000 ;
	    RECT 74.2000 74.8000 75.4000 75.1000 ;
	    RECT 79.0000 74.8000 79.4000 75.2000 ;
	    RECT 79.8000 75.1000 80.2000 75.2000 ;
	    RECT 81.4000 75.1000 81.8000 75.2000 ;
	    RECT 79.8000 74.8000 81.8000 75.1000 ;
	    RECT 68.6000 72.8000 69.0000 73.2000 ;
	    RECT 70.2000 69.2000 70.5000 74.8000 ;
	    RECT 76.6000 72.8000 77.0000 73.2000 ;
	    RECT 79.8000 72.8000 80.2000 73.2000 ;
	    RECT 75.8000 71.8000 76.2000 72.2000 ;
	    RECT 75.8000 69.2000 76.1000 71.8000 ;
	    RECT 67.8000 68.8000 68.2000 69.2000 ;
	    RECT 70.2000 68.8000 70.6000 69.2000 ;
	    RECT 75.8000 68.8000 76.2000 69.2000 ;
	    RECT 76.6000 68.2000 76.9000 72.8000 ;
	    RECT 79.8000 69.2000 80.1000 72.8000 ;
	    RECT 82.2000 72.2000 82.5000 76.8000 ;
	    RECT 82.2000 71.8000 82.6000 72.2000 ;
	    RECT 83.0000 69.2000 83.3000 85.8000 ;
	    RECT 87.0000 84.8000 87.4000 85.2000 ;
	    RECT 88.6000 84.8000 89.0000 85.2000 ;
	    RECT 89.4000 84.8000 89.8000 85.2000 ;
	    RECT 92.6000 84.8000 93.0000 85.2000 ;
	    RECT 94.2000 85.1000 94.6000 85.2000 ;
	    RECT 95.0000 85.1000 95.4000 85.2000 ;
	    RECT 94.2000 84.8000 95.4000 85.1000 ;
	    RECT 97.4000 84.8000 97.8000 85.2000 ;
	    RECT 84.6000 83.8000 85.0000 84.2000 ;
	    RECT 84.6000 79.2000 84.9000 83.8000 ;
	    RECT 86.2000 82.8000 86.6000 83.2000 ;
	    RECT 86.2000 79.2000 86.5000 82.8000 ;
	    RECT 87.0000 79.2000 87.3000 84.8000 ;
	    RECT 88.6000 84.2000 88.9000 84.8000 ;
	    RECT 88.6000 83.8000 89.0000 84.2000 ;
	    RECT 89.4000 83.2000 89.7000 84.8000 ;
	    RECT 92.6000 84.2000 92.9000 84.8000 ;
	    RECT 92.6000 83.8000 93.0000 84.2000 ;
	    RECT 95.0000 84.1000 95.4000 84.2000 ;
	    RECT 95.8000 84.1000 96.2000 84.2000 ;
	    RECT 95.0000 83.8000 96.2000 84.1000 ;
	    RECT 89.4000 82.8000 89.8000 83.2000 ;
	    RECT 92.6000 82.8000 93.0000 83.2000 ;
	    RECT 92.6000 79.2000 92.9000 82.8000 ;
	    RECT 93.4000 81.8000 93.8000 82.2000 ;
	    RECT 96.6000 81.8000 97.0000 82.2000 ;
	    RECT 93.4000 80.2000 93.7000 81.8000 ;
	    RECT 93.4000 79.8000 93.8000 80.2000 ;
	    RECT 84.6000 78.8000 85.0000 79.2000 ;
	    RECT 86.2000 78.8000 86.6000 79.2000 ;
	    RECT 87.0000 78.8000 87.4000 79.2000 ;
	    RECT 92.6000 78.8000 93.0000 79.2000 ;
	    RECT 95.0000 77.8000 95.4000 78.2000 ;
	    RECT 95.0000 77.2000 95.3000 77.8000 ;
	    RECT 93.4000 77.1000 93.8000 77.2000 ;
	    RECT 94.2000 77.1000 94.6000 77.2000 ;
	    RECT 93.4000 76.8000 94.6000 77.1000 ;
	    RECT 95.0000 76.8000 95.4000 77.2000 ;
	    RECT 95.8000 76.8000 96.2000 77.2000 ;
	    RECT 95.8000 76.2000 96.1000 76.8000 ;
	    RECT 96.6000 76.2000 96.9000 81.8000 ;
	    RECT 97.4000 77.2000 97.7000 84.8000 ;
	    RECT 98.2000 79.2000 98.5000 91.8000 ;
	    RECT 99.0000 87.8000 99.4000 88.2000 ;
	    RECT 99.0000 84.2000 99.3000 87.8000 ;
	    RECT 100.6000 87.2000 100.9000 93.8000 ;
	    RECT 104.6000 93.2000 104.9000 93.8000 ;
	    RECT 102.2000 92.8000 102.6000 93.2000 ;
	    RECT 104.6000 92.8000 105.0000 93.2000 ;
	    RECT 99.8000 86.8000 100.2000 87.2000 ;
	    RECT 100.6000 86.8000 101.0000 87.2000 ;
	    RECT 99.8000 86.2000 100.1000 86.8000 ;
	    RECT 99.8000 85.8000 100.2000 86.2000 ;
	    RECT 100.6000 84.8000 101.0000 85.2000 ;
	    RECT 101.4000 85.1000 101.8000 87.9000 ;
	    RECT 99.0000 83.8000 99.4000 84.2000 ;
	    RECT 99.8000 81.8000 100.2000 82.2000 ;
	    RECT 99.8000 81.2000 100.1000 81.8000 ;
	    RECT 99.8000 80.8000 100.2000 81.2000 ;
	    RECT 98.2000 78.8000 98.6000 79.2000 ;
	    RECT 99.8000 78.8000 100.2000 79.2000 ;
	    RECT 97.4000 76.8000 97.8000 77.2000 ;
	    RECT 95.8000 75.8000 96.2000 76.2000 ;
	    RECT 96.6000 75.8000 97.0000 76.2000 ;
	    RECT 99.8000 75.2000 100.1000 78.8000 ;
	    RECT 100.6000 77.2000 100.9000 84.8000 ;
	    RECT 100.6000 76.8000 101.0000 77.2000 ;
	    RECT 91.0000 74.8000 91.4000 75.2000 ;
	    RECT 94.2000 75.1000 94.6000 75.2000 ;
	    RECT 95.0000 75.1000 95.4000 75.2000 ;
	    RECT 94.2000 74.8000 95.4000 75.1000 ;
	    RECT 95.8000 75.1000 96.2000 75.2000 ;
	    RECT 96.6000 75.1000 97.0000 75.2000 ;
	    RECT 95.8000 74.8000 97.0000 75.1000 ;
	    RECT 98.2000 75.1000 98.6000 75.2000 ;
	    RECT 99.0000 75.1000 99.4000 75.2000 ;
	    RECT 98.2000 74.8000 99.4000 75.1000 ;
	    RECT 99.8000 74.8000 100.2000 75.2000 ;
	    RECT 88.6000 74.0000 89.0000 74.4000 ;
	    RECT 79.8000 68.8000 80.2000 69.2000 ;
	    RECT 83.0000 68.8000 83.4000 69.2000 ;
	    RECT 67.0000 67.8000 67.4000 68.2000 ;
	    RECT 71.8000 68.1000 72.2000 68.2000 ;
	    RECT 72.6000 68.1000 73.0000 68.2000 ;
	    RECT 71.8000 67.8000 73.0000 68.1000 ;
	    RECT 76.6000 67.8000 77.0000 68.2000 ;
	    RECT 77.4000 67.8000 77.8000 68.2000 ;
	    RECT 80.6000 67.8000 81.0000 68.2000 ;
	    RECT 53.4000 66.8000 53.8000 67.2000 ;
	    RECT 55.8000 66.8000 56.2000 67.2000 ;
	    RECT 66.2000 67.1000 66.6000 67.2000 ;
	    RECT 67.0000 67.1000 67.3000 67.8000 ;
	    RECT 76.6000 67.2000 76.9000 67.8000 ;
	    RECT 77.4000 67.2000 77.7000 67.8000 ;
	    RECT 80.6000 67.2000 80.9000 67.8000 ;
	    RECT 66.2000 66.8000 67.3000 67.1000 ;
	    RECT 72.6000 66.8000 73.0000 67.2000 ;
	    RECT 76.6000 66.8000 77.0000 67.2000 ;
	    RECT 77.4000 66.8000 77.8000 67.2000 ;
	    RECT 80.6000 66.8000 81.0000 67.2000 ;
	    RECT 53.4000 66.2000 53.7000 66.8000 ;
	    RECT 34.2000 65.8000 34.6000 66.2000 ;
	    RECT 44.6000 65.8000 45.0000 66.2000 ;
	    RECT 52.6000 65.8000 53.0000 66.2000 ;
	    RECT 53.4000 65.8000 53.8000 66.2000 ;
	    RECT 58.2000 65.8000 58.6000 66.2000 ;
	    RECT 34.2000 65.2000 34.5000 65.8000 ;
	    RECT 58.2000 65.2000 58.5000 65.8000 ;
	    RECT 34.2000 64.8000 34.6000 65.2000 ;
	    RECT 46.2000 64.8000 46.6000 65.2000 ;
	    RECT 48.6000 65.1000 49.0000 65.2000 ;
	    RECT 49.4000 65.1000 49.8000 65.2000 ;
	    RECT 48.6000 64.8000 49.8000 65.1000 ;
	    RECT 50.2000 65.1000 50.6000 65.2000 ;
	    RECT 51.0000 65.1000 51.4000 65.2000 ;
	    RECT 50.2000 64.8000 51.4000 65.1000 ;
	    RECT 52.6000 64.8000 53.0000 65.2000 ;
	    RECT 55.8000 64.8000 56.2000 65.2000 ;
	    RECT 57.4000 64.8000 57.8000 65.2000 ;
	    RECT 58.2000 64.8000 58.6000 65.2000 ;
	    RECT 46.2000 64.2000 46.5000 64.8000 ;
	    RECT 52.6000 64.2000 52.9000 64.8000 ;
	    RECT 41.4000 64.1000 41.8000 64.2000 ;
	    RECT 42.2000 64.1000 42.6000 64.2000 ;
	    RECT 41.4000 63.8000 42.6000 64.1000 ;
	    RECT 46.2000 63.8000 46.6000 64.2000 ;
	    RECT 52.6000 63.8000 53.0000 64.2000 ;
	    RECT 54.2000 64.1000 54.6000 64.2000 ;
	    RECT 55.0000 64.1000 55.4000 64.2000 ;
	    RECT 54.2000 63.8000 55.4000 64.1000 ;
	    RECT 31.0000 62.8000 31.4000 63.2000 ;
	    RECT 31.8000 62.8000 32.2000 63.2000 ;
	    RECT 33.4000 62.8000 33.8000 63.2000 ;
	    RECT 19.0000 61.8000 19.4000 62.2000 ;
	    RECT 23.8000 61.8000 24.2000 62.2000 ;
	    RECT 17.4000 57.8000 17.8000 58.2000 ;
	    RECT 19.0000 57.2000 19.3000 61.8000 ;
	    RECT 23.8000 61.2000 24.1000 61.8000 ;
	    RECT 23.8000 60.8000 24.2000 61.2000 ;
	    RECT 20.6000 58.8000 21.0000 59.2000 ;
	    RECT 23.0000 59.1000 23.4000 59.2000 ;
	    RECT 23.8000 59.1000 24.2000 59.2000 ;
	    RECT 23.0000 58.8000 24.2000 59.1000 ;
	    RECT 24.6000 58.8000 25.0000 59.2000 ;
	    RECT 27.0000 59.1000 27.4000 59.2000 ;
	    RECT 27.8000 59.1000 28.2000 59.2000 ;
	    RECT 27.0000 58.8000 28.2000 59.1000 ;
	    RECT 19.8000 57.8000 20.2000 58.2000 ;
	    RECT 16.6000 56.8000 17.0000 57.2000 ;
	    RECT 19.0000 56.8000 19.4000 57.2000 ;
	    RECT 19.8000 56.2000 20.1000 57.8000 ;
	    RECT 12.6000 55.8000 13.0000 56.2000 ;
	    RECT 15.8000 55.8000 16.2000 56.2000 ;
	    RECT 19.8000 55.8000 20.2000 56.2000 ;
	    RECT 20.6000 55.2000 20.9000 58.8000 ;
	    RECT 21.4000 57.8000 21.8000 58.2000 ;
	    RECT 21.4000 57.2000 21.7000 57.8000 ;
	    RECT 24.6000 57.2000 24.9000 58.8000 ;
	    RECT 21.4000 56.8000 21.8000 57.2000 ;
	    RECT 24.6000 56.8000 25.0000 57.2000 ;
	    RECT 27.0000 57.1000 27.4000 57.2000 ;
	    RECT 27.8000 57.1000 28.2000 57.2000 ;
	    RECT 27.0000 56.8000 28.2000 57.1000 ;
	    RECT 23.0000 55.8000 23.4000 56.2000 ;
	    RECT 29.4000 55.8000 29.8000 56.2000 ;
	    RECT 23.0000 55.2000 23.3000 55.8000 ;
	    RECT 29.4000 55.2000 29.7000 55.8000 ;
	    RECT 15.0000 54.8000 15.4000 55.2000 ;
	    RECT 18.2000 54.8000 18.6000 55.2000 ;
	    RECT 19.0000 55.1000 19.4000 55.2000 ;
	    RECT 19.8000 55.1000 20.2000 55.2000 ;
	    RECT 19.0000 54.8000 20.2000 55.1000 ;
	    RECT 20.6000 54.8000 21.0000 55.2000 ;
	    RECT 23.0000 54.8000 23.4000 55.2000 ;
	    RECT 23.8000 55.1000 24.2000 55.2000 ;
	    RECT 24.6000 55.1000 25.0000 55.2000 ;
	    RECT 23.8000 54.8000 25.0000 55.1000 ;
	    RECT 27.0000 55.1000 27.4000 55.2000 ;
	    RECT 27.8000 55.1000 28.2000 55.2000 ;
	    RECT 27.0000 54.8000 28.2000 55.1000 ;
	    RECT 29.4000 54.8000 29.8000 55.2000 ;
	    RECT 15.0000 54.2000 15.3000 54.8000 ;
	    RECT 18.2000 54.2000 18.5000 54.8000 ;
	    RECT 15.0000 53.8000 15.4000 54.2000 ;
	    RECT 16.6000 54.1000 17.0000 54.2000 ;
	    RECT 17.4000 54.1000 17.8000 54.2000 ;
	    RECT 16.6000 53.8000 17.8000 54.1000 ;
	    RECT 18.2000 53.8000 18.6000 54.2000 ;
	    RECT 26.2000 53.8000 26.6000 54.2000 ;
	    RECT 21.4000 53.1000 21.8000 53.2000 ;
	    RECT 22.2000 53.1000 22.6000 53.2000 ;
	    RECT 21.4000 52.8000 22.6000 53.1000 ;
	    RECT 12.6000 51.8000 13.0000 52.2000 ;
	    RECT 15.0000 51.8000 15.4000 52.2000 ;
	    RECT 11.8000 48.8000 12.2000 49.2000 ;
	    RECT 10.2000 47.8000 10.6000 48.2000 ;
	    RECT 10.2000 47.2000 10.5000 47.8000 ;
	    RECT 10.2000 46.8000 10.6000 47.2000 ;
	    RECT 10.2000 46.2000 10.5000 46.8000 ;
	    RECT 10.2000 45.8000 10.6000 46.2000 ;
	    RECT 12.6000 45.2000 12.9000 51.8000 ;
	    RECT 15.0000 47.2000 15.3000 51.8000 ;
	    RECT 26.2000 49.2000 26.5000 53.8000 ;
	    RECT 31.8000 53.2000 32.1000 62.8000 ;
	    RECT 55.8000 59.2000 56.1000 64.8000 ;
	    RECT 57.4000 64.2000 57.7000 64.8000 ;
	    RECT 57.4000 63.8000 57.8000 64.2000 ;
	    RECT 58.2000 63.8000 58.6000 64.2000 ;
	    RECT 70.2000 63.8000 70.6000 64.2000 ;
	    RECT 58.2000 59.2000 58.5000 63.8000 ;
	    RECT 70.2000 59.2000 70.5000 63.8000 ;
	    RECT 72.6000 59.2000 72.9000 66.8000 ;
	    RECT 75.8000 62.8000 76.2000 63.2000 ;
	    RECT 75.8000 59.2000 76.1000 62.8000 ;
	    RECT 77.4000 59.2000 77.7000 66.8000 ;
	    RECT 78.2000 65.8000 78.6000 66.2000 ;
	    RECT 81.4000 65.8000 81.8000 66.2000 ;
	    RECT 78.2000 65.2000 78.5000 65.8000 ;
	    RECT 78.2000 64.8000 78.6000 65.2000 ;
	    RECT 81.4000 64.2000 81.7000 65.8000 ;
	    RECT 83.8000 65.1000 84.2000 67.9000 ;
	    RECT 81.4000 63.8000 81.8000 64.2000 ;
	    RECT 85.4000 63.1000 85.8000 68.9000 ;
	    RECT 88.6000 67.1000 88.9000 74.0000 ;
	    RECT 89.4000 73.8000 89.8000 74.2000 ;
	    RECT 89.4000 68.2000 89.7000 73.8000 ;
	    RECT 89.4000 67.8000 89.8000 68.2000 ;
	    RECT 88.6000 66.8000 89.7000 67.1000 ;
	    RECT 86.2000 65.9000 86.6000 66.3000 ;
	    RECT 79.8000 61.8000 80.2000 62.2000 ;
	    RECT 79.8000 59.2000 80.1000 61.8000 ;
	    RECT 86.2000 60.2000 86.5000 65.9000 ;
	    RECT 88.6000 65.8000 89.0000 66.2000 ;
	    RECT 86.2000 59.8000 86.6000 60.2000 ;
	    RECT 44.6000 59.1000 45.0000 59.2000 ;
	    RECT 45.4000 59.1000 45.8000 59.2000 ;
	    RECT 44.6000 58.8000 45.8000 59.1000 ;
	    RECT 46.2000 58.8000 46.6000 59.2000 ;
	    RECT 55.8000 58.8000 56.2000 59.2000 ;
	    RECT 58.2000 58.8000 58.6000 59.2000 ;
	    RECT 70.2000 58.8000 70.6000 59.2000 ;
	    RECT 72.6000 58.8000 73.0000 59.2000 ;
	    RECT 75.8000 58.8000 76.2000 59.2000 ;
	    RECT 77.4000 58.8000 77.8000 59.2000 ;
	    RECT 79.8000 58.8000 80.2000 59.2000 ;
	    RECT 35.8000 57.8000 36.2000 58.2000 ;
	    RECT 35.0000 56.8000 35.4000 57.2000 ;
	    RECT 35.0000 56.2000 35.3000 56.8000 ;
	    RECT 35.0000 55.8000 35.4000 56.2000 ;
	    RECT 35.8000 55.2000 36.1000 57.8000 ;
	    RECT 38.2000 56.8000 38.6000 57.2000 ;
	    RECT 41.4000 56.8000 41.8000 57.2000 ;
	    RECT 38.2000 56.2000 38.5000 56.8000 ;
	    RECT 41.4000 56.2000 41.7000 56.8000 ;
	    RECT 38.2000 55.8000 38.6000 56.2000 ;
	    RECT 41.4000 55.8000 41.8000 56.2000 ;
	    RECT 32.6000 54.8000 33.0000 55.2000 ;
	    RECT 35.8000 54.8000 36.2000 55.2000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 39.0000 55.1000 39.4000 55.2000 ;
	    RECT 38.2000 54.8000 39.4000 55.1000 ;
	    RECT 41.4000 55.1000 41.8000 55.2000 ;
	    RECT 42.2000 55.1000 42.6000 55.2000 ;
	    RECT 41.4000 54.8000 42.6000 55.1000 ;
	    RECT 32.6000 53.2000 32.9000 54.8000 ;
	    RECT 46.2000 54.2000 46.5000 58.8000 ;
	    RECT 33.4000 53.8000 33.8000 54.2000 ;
	    RECT 36.6000 53.8000 37.0000 54.2000 ;
	    RECT 39.0000 54.1000 39.4000 54.2000 ;
	    RECT 39.8000 54.1000 40.2000 54.2000 ;
	    RECT 39.0000 53.8000 40.2000 54.1000 ;
	    RECT 41.4000 53.8000 41.8000 54.2000 ;
	    RECT 43.0000 53.8000 43.4000 54.2000 ;
	    RECT 46.2000 53.8000 46.6000 54.2000 ;
	    RECT 31.8000 52.8000 32.2000 53.2000 ;
	    RECT 32.6000 52.8000 33.0000 53.2000 ;
	    RECT 31.8000 52.2000 32.1000 52.8000 ;
	    RECT 31.8000 51.8000 32.2000 52.2000 ;
	    RECT 33.4000 51.2000 33.7000 53.8000 ;
	    RECT 35.0000 53.1000 35.4000 53.2000 ;
	    RECT 35.8000 53.1000 36.2000 53.2000 ;
	    RECT 35.0000 52.8000 36.2000 53.1000 ;
	    RECT 33.4000 50.8000 33.8000 51.2000 ;
	    RECT 15.8000 49.1000 16.2000 49.2000 ;
	    RECT 16.6000 49.1000 17.0000 49.2000 ;
	    RECT 15.8000 48.8000 17.0000 49.1000 ;
	    RECT 26.2000 48.8000 26.6000 49.2000 ;
	    RECT 19.8000 47.8000 20.2000 48.2000 ;
	    RECT 23.0000 47.8000 23.4000 48.2000 ;
	    RECT 27.8000 48.1000 28.2000 48.2000 ;
	    RECT 28.6000 48.1000 29.0000 48.2000 ;
	    RECT 27.8000 47.8000 29.0000 48.1000 ;
	    RECT 15.0000 46.8000 15.4000 47.2000 ;
	    RECT 15.0000 46.2000 15.3000 46.8000 ;
	    RECT 15.0000 45.8000 15.4000 46.2000 ;
	    RECT 18.2000 46.1000 18.6000 46.2000 ;
	    RECT 19.0000 46.1000 19.4000 46.2000 ;
	    RECT 18.2000 45.8000 19.4000 46.1000 ;
	    RECT 12.6000 44.8000 13.0000 45.2000 ;
	    RECT 15.0000 44.8000 15.4000 45.2000 ;
	    RECT 15.8000 45.1000 16.2000 45.2000 ;
	    RECT 16.6000 45.1000 17.0000 45.2000 ;
	    RECT 15.8000 44.8000 17.0000 45.1000 ;
	    RECT 15.0000 44.2000 15.3000 44.8000 ;
	    RECT 11.8000 43.8000 12.2000 44.2000 ;
	    RECT 15.0000 43.8000 15.4000 44.2000 ;
	    RECT 19.0000 44.1000 19.4000 44.2000 ;
	    RECT 19.8000 44.1000 20.1000 47.8000 ;
	    RECT 23.0000 47.2000 23.3000 47.8000 ;
	    RECT 23.0000 46.8000 23.4000 47.2000 ;
	    RECT 27.0000 46.8000 27.4000 47.2000 ;
	    RECT 20.6000 46.1000 21.0000 46.2000 ;
	    RECT 21.4000 46.1000 21.8000 46.2000 ;
	    RECT 20.6000 45.8000 21.8000 46.1000 ;
	    RECT 24.6000 45.8000 25.0000 46.2000 ;
	    RECT 19.0000 43.8000 20.1000 44.1000 ;
	    RECT 11.8000 39.2000 12.1000 43.8000 ;
	    RECT 18.2000 42.8000 18.6000 43.2000 ;
	    RECT 18.2000 42.2000 18.5000 42.8000 ;
	    RECT 24.6000 42.2000 24.9000 45.8000 ;
	    RECT 25.4000 43.8000 25.8000 44.2000 ;
	    RECT 25.4000 43.2000 25.7000 43.8000 ;
	    RECT 25.4000 42.8000 25.8000 43.2000 ;
	    RECT 18.2000 41.8000 18.6000 42.2000 ;
	    RECT 24.6000 41.8000 25.0000 42.2000 ;
	    RECT 15.0000 39.8000 15.4000 40.2000 ;
	    RECT 15.0000 39.2000 15.3000 39.8000 ;
	    RECT 9.4000 38.8000 9.8000 39.2000 ;
	    RECT 11.8000 38.8000 12.2000 39.2000 ;
	    RECT 15.0000 38.8000 15.4000 39.2000 ;
	    RECT 17.4000 37.8000 17.8000 38.2000 ;
	    RECT 23.0000 37.8000 23.4000 38.2000 ;
	    RECT 1.4000 37.1000 1.8000 37.2000 ;
	    RECT 2.2000 37.1000 2.6000 37.2000 ;
	    RECT 1.4000 36.8000 2.6000 37.1000 ;
	    RECT 4.6000 36.8000 5.0000 37.2000 ;
	    RECT 8.6000 36.8000 9.0000 37.2000 ;
	    RECT 11.0000 36.8000 11.4000 37.2000 ;
	    RECT 3.0000 35.8000 3.4000 36.2000 ;
	    RECT 5.4000 36.1000 5.8000 36.2000 ;
	    RECT 6.2000 36.1000 6.6000 36.2000 ;
	    RECT 5.4000 35.8000 6.6000 36.1000 ;
	    RECT 2.2000 34.8000 2.6000 35.2000 ;
	    RECT 0.6000 34.1000 1.0000 34.2000 ;
	    RECT 1.4000 34.1000 1.8000 34.2000 ;
	    RECT 0.6000 33.8000 1.8000 34.1000 ;
	    RECT 1.4000 32.8000 1.8000 33.2000 ;
	    RECT 1.4000 19.2000 1.7000 32.8000 ;
	    RECT 2.2000 32.2000 2.5000 34.8000 ;
	    RECT 3.0000 33.2000 3.3000 35.8000 ;
	    RECT 4.6000 34.8000 5.0000 35.2000 ;
	    RECT 5.4000 34.8000 5.8000 35.2000 ;
	    RECT 7.0000 35.1000 7.4000 35.2000 ;
	    RECT 7.8000 35.1000 8.2000 35.2000 ;
	    RECT 7.0000 34.8000 8.2000 35.1000 ;
	    RECT 4.6000 34.2000 4.9000 34.8000 ;
	    RECT 5.4000 34.2000 5.7000 34.8000 ;
	    RECT 4.6000 33.8000 5.0000 34.2000 ;
	    RECT 5.4000 33.8000 5.8000 34.2000 ;
	    RECT 3.0000 32.8000 3.4000 33.2000 ;
	    RECT 2.2000 31.8000 2.6000 32.2000 ;
	    RECT 4.6000 31.8000 5.0000 32.2000 ;
	    RECT 2.2000 30.8000 2.6000 31.2000 ;
	    RECT 2.2000 29.2000 2.5000 30.8000 ;
	    RECT 4.6000 29.2000 4.9000 31.8000 ;
	    RECT 8.6000 29.2000 8.9000 36.8000 ;
	    RECT 11.0000 35.2000 11.3000 36.8000 ;
	    RECT 16.6000 35.8000 17.0000 36.2000 ;
	    RECT 16.6000 35.2000 16.9000 35.8000 ;
	    RECT 17.4000 35.2000 17.7000 37.8000 ;
	    RECT 23.0000 37.2000 23.3000 37.8000 ;
	    RECT 18.2000 36.8000 18.6000 37.2000 ;
	    RECT 19.8000 36.8000 20.2000 37.2000 ;
	    RECT 23.0000 36.8000 23.4000 37.2000 ;
	    RECT 23.8000 37.1000 24.2000 37.2000 ;
	    RECT 23.8000 36.8000 24.9000 37.1000 ;
	    RECT 18.2000 36.2000 18.5000 36.8000 ;
	    RECT 19.8000 36.2000 20.1000 36.8000 ;
	    RECT 18.2000 35.8000 18.6000 36.2000 ;
	    RECT 19.8000 35.8000 20.2000 36.2000 ;
	    RECT 21.4000 35.8000 21.8000 36.2000 ;
	    RECT 22.2000 36.1000 22.6000 36.2000 ;
	    RECT 23.0000 36.1000 23.4000 36.2000 ;
	    RECT 22.2000 35.8000 23.4000 36.1000 ;
	    RECT 21.4000 35.2000 21.7000 35.8000 ;
	    RECT 11.0000 34.8000 11.4000 35.2000 ;
	    RECT 11.8000 35.1000 12.2000 35.2000 ;
	    RECT 12.6000 35.1000 13.0000 35.2000 ;
	    RECT 11.8000 34.8000 13.0000 35.1000 ;
	    RECT 15.0000 34.8000 15.4000 35.2000 ;
	    RECT 16.6000 34.8000 17.0000 35.2000 ;
	    RECT 17.4000 34.8000 17.8000 35.2000 ;
	    RECT 18.2000 34.8000 18.6000 35.2000 ;
	    RECT 21.4000 34.8000 21.8000 35.2000 ;
	    RECT 15.0000 29.2000 15.3000 34.8000 ;
	    RECT 18.2000 29.2000 18.5000 34.8000 ;
	    RECT 22.2000 33.2000 22.5000 35.8000 ;
	    RECT 23.0000 35.1000 23.4000 35.2000 ;
	    RECT 23.8000 35.1000 24.2000 35.2000 ;
	    RECT 23.0000 34.8000 24.2000 35.1000 ;
	    RECT 24.6000 33.2000 24.9000 36.8000 ;
	    RECT 25.4000 34.8000 25.8000 35.2000 ;
	    RECT 25.4000 34.2000 25.7000 34.8000 ;
	    RECT 25.4000 33.8000 25.8000 34.2000 ;
	    RECT 22.2000 32.8000 22.6000 33.2000 ;
	    RECT 24.6000 32.8000 25.0000 33.2000 ;
	    RECT 21.4000 31.8000 21.8000 32.2000 ;
	    RECT 21.4000 29.2000 21.7000 31.8000 ;
	    RECT 2.2000 28.8000 2.6000 29.2000 ;
	    RECT 4.6000 28.8000 5.0000 29.2000 ;
	    RECT 8.6000 28.8000 9.0000 29.2000 ;
	    RECT 11.0000 28.8000 11.4000 29.2000 ;
	    RECT 15.0000 28.8000 15.4000 29.2000 ;
	    RECT 18.2000 28.8000 18.6000 29.2000 ;
	    RECT 21.4000 28.8000 21.8000 29.2000 ;
	    RECT 11.0000 28.2000 11.3000 28.8000 ;
	    RECT 3.8000 27.8000 4.2000 28.2000 ;
	    RECT 6.2000 27.8000 6.6000 28.2000 ;
	    RECT 11.0000 27.8000 11.4000 28.2000 ;
	    RECT 3.8000 27.2000 4.1000 27.8000 ;
	    RECT 6.2000 27.2000 6.5000 27.8000 ;
	    RECT 3.8000 26.8000 4.2000 27.2000 ;
	    RECT 6.2000 26.8000 6.6000 27.2000 ;
	    RECT 1.4000 18.8000 1.8000 19.2000 ;
	    RECT 5.4000 18.8000 5.8000 19.2000 ;
	    RECT 1.4000 16.8000 1.8000 17.2000 ;
	    RECT 3.0000 17.1000 3.4000 17.2000 ;
	    RECT 3.8000 17.1000 4.2000 17.2000 ;
	    RECT 3.0000 16.8000 4.2000 17.1000 ;
	    RECT 1.4000 9.2000 1.7000 16.8000 ;
	    RECT 5.4000 16.2000 5.7000 18.8000 ;
	    RECT 6.2000 17.2000 6.5000 26.8000 ;
	    RECT 9.4000 25.8000 9.8000 26.2000 ;
	    RECT 11.0000 25.8000 11.4000 26.2000 ;
	    RECT 14.2000 25.8000 14.6000 26.2000 ;
	    RECT 17.4000 25.8000 17.8000 26.2000 ;
	    RECT 7.0000 23.8000 7.4000 24.2000 ;
	    RECT 7.8000 24.1000 8.2000 24.2000 ;
	    RECT 8.6000 24.1000 9.0000 24.2000 ;
	    RECT 7.8000 23.8000 9.0000 24.1000 ;
	    RECT 6.2000 16.8000 6.6000 17.2000 ;
	    RECT 5.4000 15.8000 5.8000 16.2000 ;
	    RECT 6.2000 15.8000 6.6000 16.2000 ;
	    RECT 6.2000 15.2000 6.5000 15.8000 ;
	    RECT 4.6000 15.1000 5.0000 15.2000 ;
	    RECT 5.4000 15.1000 5.8000 15.2000 ;
	    RECT 4.6000 14.8000 5.8000 15.1000 ;
	    RECT 6.2000 14.8000 6.6000 15.2000 ;
	    RECT 4.6000 13.8000 5.0000 14.2000 ;
	    RECT 4.6000 13.2000 4.9000 13.8000 ;
	    RECT 4.6000 12.8000 5.0000 13.2000 ;
	    RECT 7.0000 9.2000 7.3000 23.8000 ;
	    RECT 9.4000 23.2000 9.7000 25.8000 ;
	    RECT 9.4000 22.8000 9.8000 23.2000 ;
	    RECT 11.0000 19.2000 11.3000 25.8000 ;
	    RECT 14.2000 24.2000 14.5000 25.8000 ;
	    RECT 14.2000 23.8000 14.6000 24.2000 ;
	    RECT 15.0000 23.8000 15.4000 24.2000 ;
	    RECT 15.0000 19.2000 15.3000 23.8000 ;
	    RECT 17.4000 22.2000 17.7000 25.8000 ;
	    RECT 22.2000 25.2000 22.5000 32.8000 ;
	    RECT 27.0000 32.2000 27.3000 46.8000 ;
	    RECT 28.6000 45.8000 29.0000 46.2000 ;
	    RECT 30.2000 45.8000 30.6000 46.2000 ;
	    RECT 34.2000 46.1000 34.6000 46.2000 ;
	    RECT 35.8000 46.1000 36.2000 46.2000 ;
	    RECT 34.2000 45.8000 36.2000 46.1000 ;
	    RECT 28.6000 45.2000 28.9000 45.8000 ;
	    RECT 28.6000 44.8000 29.0000 45.2000 ;
	    RECT 30.2000 43.1000 30.5000 45.8000 ;
	    RECT 31.0000 44.1000 31.4000 44.2000 ;
	    RECT 31.8000 44.1000 32.2000 44.2000 ;
	    RECT 31.0000 43.8000 32.2000 44.1000 ;
	    RECT 33.4000 43.8000 33.8000 44.2000 ;
	    RECT 34.2000 44.1000 34.6000 44.2000 ;
	    RECT 35.0000 44.1000 35.4000 44.2000 ;
	    RECT 34.2000 43.8000 35.4000 44.1000 ;
	    RECT 33.4000 43.2000 33.7000 43.8000 ;
	    RECT 30.2000 42.8000 31.3000 43.1000 ;
	    RECT 33.4000 42.8000 33.8000 43.2000 ;
	    RECT 30.2000 41.8000 30.6000 42.2000 ;
	    RECT 30.2000 41.2000 30.5000 41.8000 ;
	    RECT 30.2000 40.8000 30.6000 41.2000 ;
	    RECT 31.0000 39.2000 31.3000 42.8000 ;
	    RECT 36.6000 40.2000 36.9000 53.8000 ;
	    RECT 41.4000 53.2000 41.7000 53.8000 ;
	    RECT 38.2000 53.1000 38.6000 53.2000 ;
	    RECT 39.0000 53.1000 39.4000 53.2000 ;
	    RECT 38.2000 52.8000 39.4000 53.1000 ;
	    RECT 41.4000 52.8000 41.8000 53.2000 ;
	    RECT 43.0000 50.2000 43.3000 53.8000 ;
	    RECT 43.8000 53.1000 44.2000 53.2000 ;
	    RECT 44.6000 53.1000 45.0000 53.2000 ;
	    RECT 47.0000 53.1000 47.4000 55.9000 ;
	    RECT 43.8000 52.8000 45.0000 53.1000 ;
	    RECT 48.6000 52.1000 49.0000 57.9000 ;
	    RECT 52.6000 57.8000 53.0000 58.2000 ;
	    RECT 52.6000 55.2000 52.9000 57.8000 ;
	    RECT 49.4000 54.7000 49.8000 55.1000 ;
	    RECT 52.6000 54.8000 53.0000 55.2000 ;
	    RECT 49.4000 54.2000 49.7000 54.7000 ;
	    RECT 49.4000 53.8000 49.8000 54.2000 ;
	    RECT 53.4000 52.1000 53.8000 57.9000 ;
	    RECT 57.4000 57.1000 57.8000 57.2000 ;
	    RECT 56.6000 56.8000 57.8000 57.1000 ;
	    RECT 43.0000 49.8000 43.4000 50.2000 ;
	    RECT 38.2000 47.8000 38.6000 48.2000 ;
	    RECT 41.4000 47.8000 41.8000 48.2000 ;
	    RECT 43.8000 47.8000 44.2000 48.2000 ;
	    RECT 38.2000 47.2000 38.5000 47.8000 ;
	    RECT 41.4000 47.2000 41.7000 47.8000 ;
	    RECT 43.8000 47.2000 44.1000 47.8000 ;
	    RECT 38.2000 46.8000 38.6000 47.2000 ;
	    RECT 40.6000 46.8000 41.0000 47.2000 ;
	    RECT 41.4000 46.8000 41.8000 47.2000 ;
	    RECT 43.8000 46.8000 44.2000 47.2000 ;
	    RECT 45.4000 46.8000 45.8000 47.2000 ;
	    RECT 53.4000 46.8000 53.8000 47.2000 ;
	    RECT 40.6000 45.2000 40.9000 46.8000 ;
	    RECT 45.4000 46.2000 45.7000 46.8000 ;
	    RECT 45.4000 45.8000 45.8000 46.2000 ;
	    RECT 47.0000 45.8000 47.4000 46.2000 ;
	    RECT 47.0000 45.2000 47.3000 45.8000 ;
	    RECT 40.6000 44.8000 41.0000 45.2000 ;
	    RECT 45.4000 45.1000 45.8000 45.2000 ;
	    RECT 46.2000 45.1000 46.6000 45.2000 ;
	    RECT 45.4000 44.8000 46.6000 45.1000 ;
	    RECT 47.0000 44.8000 47.4000 45.2000 ;
	    RECT 43.8000 44.1000 44.2000 44.2000 ;
	    RECT 44.6000 44.1000 45.0000 44.2000 ;
	    RECT 43.8000 43.8000 45.0000 44.1000 ;
	    RECT 51.8000 43.8000 52.2000 44.2000 ;
	    RECT 51.8000 43.2000 52.1000 43.8000 ;
	    RECT 51.8000 42.8000 52.2000 43.2000 ;
	    RECT 52.6000 42.8000 53.0000 43.2000 ;
	    RECT 39.8000 41.8000 40.2000 42.2000 ;
	    RECT 42.2000 41.8000 42.6000 42.2000 ;
	    RECT 36.6000 39.8000 37.0000 40.2000 ;
	    RECT 31.0000 38.8000 31.4000 39.2000 ;
	    RECT 39.8000 38.2000 40.1000 41.8000 ;
	    RECT 30.2000 37.8000 30.6000 38.2000 ;
	    RECT 39.8000 37.8000 40.2000 38.2000 ;
	    RECT 30.2000 37.2000 30.5000 37.8000 ;
	    RECT 30.2000 36.8000 30.6000 37.2000 ;
	    RECT 42.2000 36.2000 42.5000 41.8000 ;
	    RECT 52.6000 39.2000 52.9000 42.8000 ;
	    RECT 52.6000 38.8000 53.0000 39.2000 ;
	    RECT 49.4000 37.8000 49.8000 38.2000 ;
	    RECT 51.0000 37.8000 51.4000 38.2000 ;
	    RECT 47.8000 37.1000 48.2000 37.2000 ;
	    RECT 47.0000 36.8000 48.2000 37.1000 ;
	    RECT 28.6000 36.1000 29.0000 36.2000 ;
	    RECT 29.4000 36.1000 29.8000 36.2000 ;
	    RECT 28.6000 35.8000 29.8000 36.1000 ;
	    RECT 31.8000 35.8000 32.2000 36.2000 ;
	    RECT 39.0000 36.1000 39.4000 36.2000 ;
	    RECT 39.8000 36.1000 40.2000 36.2000 ;
	    RECT 39.0000 35.8000 40.2000 36.1000 ;
	    RECT 42.2000 35.8000 42.6000 36.2000 ;
	    RECT 43.8000 35.8000 44.2000 36.2000 ;
	    RECT 31.8000 35.2000 32.1000 35.8000 ;
	    RECT 28.6000 35.1000 29.0000 35.2000 ;
	    RECT 29.4000 35.1000 29.8000 35.2000 ;
	    RECT 28.6000 34.8000 29.8000 35.1000 ;
	    RECT 31.8000 34.8000 32.2000 35.2000 ;
	    RECT 39.0000 34.8000 39.4000 35.2000 ;
	    RECT 40.6000 34.8000 41.0000 35.2000 ;
	    RECT 39.0000 34.2000 39.3000 34.8000 ;
	    RECT 39.0000 33.8000 39.4000 34.2000 ;
	    RECT 27.8000 32.8000 28.2000 33.2000 ;
	    RECT 34.2000 32.8000 34.6000 33.2000 ;
	    RECT 35.8000 33.1000 36.2000 33.2000 ;
	    RECT 36.6000 33.1000 37.0000 33.2000 ;
	    RECT 35.8000 32.8000 37.0000 33.1000 ;
	    RECT 27.0000 31.8000 27.4000 32.2000 ;
	    RECT 27.8000 28.2000 28.1000 32.8000 ;
	    RECT 34.2000 29.2000 34.5000 32.8000 ;
	    RECT 40.6000 29.2000 40.9000 34.8000 ;
	    RECT 43.8000 33.2000 44.1000 35.8000 ;
	    RECT 46.2000 34.8000 46.6000 35.2000 ;
	    RECT 46.2000 34.2000 46.5000 34.8000 ;
	    RECT 46.2000 33.8000 46.6000 34.2000 ;
	    RECT 43.8000 32.8000 44.2000 33.2000 ;
	    RECT 30.2000 28.8000 30.6000 29.2000 ;
	    RECT 34.2000 28.8000 34.6000 29.2000 ;
	    RECT 39.0000 28.8000 39.4000 29.2000 ;
	    RECT 40.6000 28.8000 41.0000 29.2000 ;
	    RECT 30.2000 28.2000 30.5000 28.8000 ;
	    RECT 39.0000 28.2000 39.3000 28.8000 ;
	    RECT 27.8000 28.1000 28.2000 28.2000 ;
	    RECT 28.6000 28.1000 29.0000 28.2000 ;
	    RECT 27.8000 27.8000 29.0000 28.1000 ;
	    RECT 30.2000 27.8000 30.6000 28.2000 ;
	    RECT 32.6000 27.8000 33.0000 28.2000 ;
	    RECT 39.0000 27.8000 39.4000 28.2000 ;
	    RECT 39.8000 27.8000 40.2000 28.2000 ;
	    RECT 23.0000 26.8000 23.4000 27.2000 ;
	    RECT 22.2000 24.8000 22.6000 25.2000 ;
	    RECT 23.0000 24.2000 23.3000 26.8000 ;
	    RECT 23.8000 26.1000 24.2000 26.2000 ;
	    RECT 25.4000 26.1000 25.8000 26.2000 ;
	    RECT 23.8000 25.8000 25.8000 26.1000 ;
	    RECT 32.6000 25.2000 32.9000 27.8000 ;
	    RECT 39.8000 27.2000 40.1000 27.8000 ;
	    RECT 36.6000 26.8000 37.0000 27.2000 ;
	    RECT 39.8000 26.8000 40.2000 27.2000 ;
	    RECT 43.8000 27.1000 44.1000 32.8000 ;
	    RECT 47.0000 29.2000 47.3000 36.8000 ;
	    RECT 49.4000 36.2000 49.7000 37.8000 ;
	    RECT 49.4000 35.8000 49.8000 36.2000 ;
	    RECT 47.8000 35.1000 48.2000 35.2000 ;
	    RECT 48.6000 35.1000 49.0000 35.2000 ;
	    RECT 47.8000 34.8000 49.0000 35.1000 ;
	    RECT 48.6000 33.8000 49.0000 34.2000 ;
	    RECT 48.6000 33.2000 48.9000 33.8000 ;
	    RECT 48.6000 32.8000 49.0000 33.2000 ;
	    RECT 47.0000 28.8000 47.4000 29.2000 ;
	    RECT 49.4000 28.1000 49.8000 28.2000 ;
	    RECT 50.2000 28.1000 50.6000 28.2000 ;
	    RECT 49.4000 27.8000 50.6000 28.1000 ;
	    RECT 44.6000 27.1000 45.0000 27.2000 ;
	    RECT 43.8000 26.8000 45.0000 27.1000 ;
	    RECT 36.6000 26.2000 36.9000 26.8000 ;
	    RECT 34.2000 26.1000 34.6000 26.2000 ;
	    RECT 35.0000 26.1000 35.4000 26.2000 ;
	    RECT 34.2000 25.8000 35.4000 26.1000 ;
	    RECT 36.6000 25.8000 37.0000 26.2000 ;
	    RECT 26.2000 24.8000 26.6000 25.2000 ;
	    RECT 31.0000 24.8000 31.4000 25.2000 ;
	    RECT 31.8000 24.8000 32.2000 25.2000 ;
	    RECT 32.6000 24.8000 33.0000 25.2000 ;
	    RECT 33.4000 25.1000 33.8000 25.2000 ;
	    RECT 34.2000 25.1000 34.6000 25.2000 ;
	    RECT 33.4000 24.8000 34.6000 25.1000 ;
	    RECT 44.6000 25.1000 45.0000 25.2000 ;
	    RECT 45.4000 25.1000 45.8000 25.2000 ;
	    RECT 44.6000 24.8000 45.8000 25.1000 ;
	    RECT 18.2000 23.8000 18.6000 24.2000 ;
	    RECT 19.8000 23.8000 20.2000 24.2000 ;
	    RECT 23.0000 23.8000 23.4000 24.2000 ;
	    RECT 17.4000 21.8000 17.8000 22.2000 ;
	    RECT 18.2000 21.2000 18.5000 23.8000 ;
	    RECT 18.2000 20.8000 18.6000 21.2000 ;
	    RECT 19.8000 19.2000 20.1000 23.8000 ;
	    RECT 23.0000 23.1000 23.4000 23.2000 ;
	    RECT 23.8000 23.1000 24.2000 23.2000 ;
	    RECT 23.0000 22.8000 24.2000 23.1000 ;
	    RECT 23.8000 20.8000 24.2000 21.2000 ;
	    RECT 23.8000 19.2000 24.1000 20.8000 ;
	    RECT 11.0000 18.8000 11.4000 19.2000 ;
	    RECT 15.0000 18.8000 15.4000 19.2000 ;
	    RECT 19.8000 18.8000 20.2000 19.2000 ;
	    RECT 23.8000 18.8000 24.2000 19.2000 ;
	    RECT 21.4000 17.8000 21.8000 18.2000 ;
	    RECT 21.4000 17.2000 21.7000 17.8000 ;
	    RECT 8.6000 16.8000 9.0000 17.2000 ;
	    RECT 10.2000 16.8000 10.6000 17.2000 ;
	    RECT 15.8000 16.8000 16.2000 17.2000 ;
	    RECT 19.0000 17.1000 19.4000 17.2000 ;
	    RECT 19.8000 17.1000 20.2000 17.2000 ;
	    RECT 19.0000 16.8000 20.2000 17.1000 ;
	    RECT 21.4000 16.8000 21.8000 17.2000 ;
	    RECT 22.2000 16.8000 22.6000 17.2000 ;
	    RECT 24.6000 16.8000 25.0000 17.2000 ;
	    RECT 8.6000 13.2000 8.9000 16.8000 ;
	    RECT 10.2000 13.2000 10.5000 16.8000 ;
	    RECT 12.6000 15.8000 13.0000 16.2000 ;
	    RECT 12.6000 15.2000 12.9000 15.8000 ;
	    RECT 11.0000 14.8000 11.4000 15.2000 ;
	    RECT 12.6000 14.8000 13.0000 15.2000 ;
	    RECT 15.0000 14.8000 15.4000 15.2000 ;
	    RECT 11.0000 14.2000 11.3000 14.8000 ;
	    RECT 11.0000 13.8000 11.4000 14.2000 ;
	    RECT 8.6000 12.8000 9.0000 13.2000 ;
	    RECT 10.2000 12.8000 10.6000 13.2000 ;
	    RECT 1.4000 8.8000 1.8000 9.2000 ;
	    RECT 7.0000 8.8000 7.4000 9.2000 ;
	    RECT 8.6000 8.2000 8.9000 12.8000 ;
	    RECT 15.0000 9.2000 15.3000 14.8000 ;
	    RECT 15.8000 14.2000 16.1000 16.8000 ;
	    RECT 22.2000 16.2000 22.5000 16.8000 ;
	    RECT 17.4000 16.1000 17.8000 16.2000 ;
	    RECT 18.2000 16.1000 18.6000 16.2000 ;
	    RECT 17.4000 15.8000 18.6000 16.1000 ;
	    RECT 22.2000 15.8000 22.6000 16.2000 ;
	    RECT 18.2000 15.1000 18.6000 15.2000 ;
	    RECT 19.0000 15.1000 19.4000 15.2000 ;
	    RECT 18.2000 14.8000 19.4000 15.1000 ;
	    RECT 23.8000 14.8000 24.2000 15.2000 ;
	    RECT 23.8000 14.2000 24.1000 14.8000 ;
	    RECT 24.6000 14.2000 24.9000 16.8000 ;
	    RECT 26.2000 16.2000 26.5000 24.8000 ;
	    RECT 31.0000 24.2000 31.3000 24.8000 ;
	    RECT 31.0000 23.8000 31.4000 24.2000 ;
	    RECT 27.0000 21.8000 27.4000 22.2000 ;
	    RECT 27.0000 19.2000 27.3000 21.8000 ;
	    RECT 27.0000 18.8000 27.4000 19.2000 ;
	    RECT 27.8000 17.1000 28.2000 17.2000 ;
	    RECT 28.6000 17.1000 29.0000 17.2000 ;
	    RECT 27.8000 16.8000 29.0000 17.1000 ;
	    RECT 30.2000 16.8000 30.6000 17.2000 ;
	    RECT 26.2000 15.8000 26.6000 16.2000 ;
	    RECT 27.0000 15.1000 27.4000 15.2000 ;
	    RECT 27.8000 15.1000 28.2000 15.2000 ;
	    RECT 27.0000 14.8000 28.2000 15.1000 ;
	    RECT 15.8000 13.8000 16.2000 14.2000 ;
	    RECT 23.0000 13.8000 23.4000 14.2000 ;
	    RECT 23.8000 13.8000 24.2000 14.2000 ;
	    RECT 24.6000 13.8000 25.0000 14.2000 ;
	    RECT 27.0000 13.8000 27.4000 14.2000 ;
	    RECT 17.4000 12.8000 17.8000 13.2000 ;
	    RECT 17.4000 9.2000 17.7000 12.8000 ;
	    RECT 23.0000 9.2000 23.3000 13.8000 ;
	    RECT 27.0000 9.2000 27.3000 13.8000 ;
	    RECT 30.2000 9.2000 30.5000 16.8000 ;
	    RECT 31.8000 16.2000 32.1000 24.8000 ;
	    RECT 34.2000 23.8000 34.6000 24.2000 ;
	    RECT 35.0000 24.1000 35.4000 24.2000 ;
	    RECT 35.0000 23.8000 36.1000 24.1000 ;
	    RECT 34.2000 23.2000 34.5000 23.8000 ;
	    RECT 34.2000 22.8000 34.6000 23.2000 ;
	    RECT 32.6000 18.8000 33.0000 19.2000 ;
	    RECT 32.6000 18.2000 32.9000 18.8000 ;
	    RECT 32.6000 17.8000 33.0000 18.2000 ;
	    RECT 33.4000 17.1000 33.8000 17.2000 ;
	    RECT 33.4000 16.8000 34.5000 17.1000 ;
	    RECT 31.8000 15.8000 32.2000 16.2000 ;
	    RECT 32.6000 15.1000 33.0000 15.2000 ;
	    RECT 33.4000 15.1000 33.8000 15.2000 ;
	    RECT 32.6000 14.8000 33.8000 15.1000 ;
	    RECT 31.0000 13.8000 31.4000 14.2000 ;
	    RECT 31.0000 13.2000 31.3000 13.8000 ;
	    RECT 31.0000 12.8000 31.4000 13.2000 ;
	    RECT 34.2000 9.2000 34.5000 16.8000 ;
	    RECT 35.0000 15.8000 35.4000 16.2000 ;
	    RECT 35.0000 15.2000 35.3000 15.8000 ;
	    RECT 35.0000 14.8000 35.4000 15.2000 ;
	    RECT 35.8000 9.2000 36.1000 23.8000 ;
	    RECT 49.4000 21.8000 49.8000 22.2000 ;
	    RECT 49.4000 19.2000 49.7000 21.8000 ;
	    RECT 49.4000 18.8000 49.8000 19.2000 ;
	    RECT 45.4000 17.1000 45.8000 17.2000 ;
	    RECT 46.2000 17.1000 46.6000 17.2000 ;
	    RECT 45.4000 16.8000 46.6000 17.1000 ;
	    RECT 50.2000 16.8000 50.6000 17.2000 ;
	    RECT 38.2000 15.8000 38.6000 16.2000 ;
	    RECT 47.0000 15.8000 47.4000 16.2000 ;
	    RECT 38.2000 15.2000 38.5000 15.8000 ;
	    RECT 38.2000 14.8000 38.6000 15.2000 ;
	    RECT 41.4000 14.8000 41.8000 15.2000 ;
	    RECT 44.6000 14.8000 45.0000 15.2000 ;
	    RECT 45.4000 14.8000 45.8000 15.2000 ;
	    RECT 41.4000 14.2000 41.7000 14.8000 ;
	    RECT 44.6000 14.2000 44.9000 14.8000 ;
	    RECT 41.4000 13.8000 41.8000 14.2000 ;
	    RECT 44.6000 13.8000 45.0000 14.2000 ;
	    RECT 45.4000 13.2000 45.7000 14.8000 ;
	    RECT 36.6000 13.1000 37.0000 13.2000 ;
	    RECT 37.4000 13.1000 37.8000 13.2000 ;
	    RECT 36.6000 12.8000 37.8000 13.1000 ;
	    RECT 39.8000 13.1000 40.2000 13.2000 ;
	    RECT 40.6000 13.1000 41.0000 13.2000 ;
	    RECT 39.8000 12.8000 41.0000 13.1000 ;
	    RECT 41.4000 12.8000 41.8000 13.2000 ;
	    RECT 43.0000 13.1000 43.4000 13.2000 ;
	    RECT 43.8000 13.1000 44.2000 13.2000 ;
	    RECT 43.0000 12.8000 44.2000 13.1000 ;
	    RECT 45.4000 13.1000 45.8000 13.2000 ;
	    RECT 45.4000 12.8000 46.5000 13.1000 ;
	    RECT 12.6000 8.8000 13.0000 9.2000 ;
	    RECT 15.0000 8.8000 15.4000 9.2000 ;
	    RECT 17.4000 8.8000 17.8000 9.2000 ;
	    RECT 23.0000 8.8000 23.4000 9.2000 ;
	    RECT 27.0000 8.8000 27.4000 9.2000 ;
	    RECT 30.2000 8.8000 30.6000 9.2000 ;
	    RECT 34.2000 8.8000 34.6000 9.2000 ;
	    RECT 35.8000 8.8000 36.2000 9.2000 ;
	    RECT 12.6000 8.2000 12.9000 8.8000 ;
	    RECT 8.6000 7.8000 9.0000 8.2000 ;
	    RECT 12.6000 7.8000 13.0000 8.2000 ;
	    RECT 8.6000 7.2000 8.9000 7.8000 ;
	    RECT 0.6000 7.1000 1.0000 7.2000 ;
	    RECT 1.4000 7.1000 1.8000 7.2000 ;
	    RECT 0.6000 6.8000 1.8000 7.1000 ;
	    RECT 3.0000 7.1000 3.4000 7.2000 ;
	    RECT 3.8000 7.1000 4.2000 7.2000 ;
	    RECT 3.0000 6.8000 4.2000 7.1000 ;
	    RECT 8.6000 6.8000 9.0000 7.2000 ;
	    RECT 22.2000 6.8000 22.6000 7.2000 ;
	    RECT 25.4000 7.1000 25.8000 7.2000 ;
	    RECT 26.2000 7.1000 26.6000 7.2000 ;
	    RECT 25.4000 6.8000 26.6000 7.1000 ;
	    RECT 27.8000 7.1000 28.2000 7.2000 ;
	    RECT 28.6000 7.1000 29.0000 7.2000 ;
	    RECT 27.8000 6.8000 29.0000 7.1000 ;
	    RECT 31.8000 7.1000 32.2000 7.2000 ;
	    RECT 32.6000 7.1000 33.0000 7.2000 ;
	    RECT 31.8000 6.8000 33.0000 7.1000 ;
	    RECT 34.2000 7.1000 34.6000 7.2000 ;
	    RECT 35.0000 7.1000 35.4000 7.2000 ;
	    RECT 34.2000 6.8000 35.4000 7.1000 ;
	    RECT 35.8000 7.1000 36.2000 7.2000 ;
	    RECT 36.6000 7.1000 37.0000 7.2000 ;
	    RECT 35.8000 6.8000 37.0000 7.1000 ;
	    RECT 37.4000 6.8000 37.8000 7.2000 ;
	    RECT 2.2000 5.8000 2.6000 6.2000 ;
	    RECT 8.6000 6.1000 8.9000 6.8000 ;
	    RECT 22.2000 6.2000 22.5000 6.8000 ;
	    RECT 9.4000 6.1000 9.8000 6.2000 ;
	    RECT 8.6000 5.8000 9.8000 6.1000 ;
	    RECT 15.8000 6.1000 16.2000 6.2000 ;
	    RECT 16.6000 6.1000 17.0000 6.2000 ;
	    RECT 15.8000 5.8000 17.0000 6.1000 ;
	    RECT 22.2000 5.8000 22.6000 6.2000 ;
	    RECT 2.2000 5.2000 2.5000 5.8000 ;
	    RECT 37.4000 5.2000 37.7000 6.8000 ;
	    RECT 41.4000 6.2000 41.7000 12.8000 ;
	    RECT 46.2000 7.2000 46.5000 12.8000 ;
	    RECT 47.0000 9.2000 47.3000 15.8000 ;
	    RECT 47.8000 14.8000 48.2000 15.2000 ;
	    RECT 47.8000 14.2000 48.1000 14.8000 ;
	    RECT 50.2000 14.2000 50.5000 16.8000 ;
	    RECT 51.0000 16.2000 51.3000 37.8000 ;
	    RECT 53.4000 36.2000 53.7000 46.8000 ;
	    RECT 55.8000 44.8000 56.2000 45.2000 ;
	    RECT 55.8000 44.2000 56.1000 44.8000 ;
	    RECT 55.8000 43.8000 56.2000 44.2000 ;
	    RECT 56.6000 43.1000 56.9000 56.8000 ;
	    RECT 57.4000 55.1000 57.8000 55.2000 ;
	    RECT 58.2000 55.1000 58.6000 55.2000 ;
	    RECT 57.4000 54.8000 58.6000 55.1000 ;
	    RECT 61.4000 53.1000 61.8000 55.9000 ;
	    RECT 63.0000 52.1000 63.4000 57.9000 ;
	    RECT 67.0000 57.8000 67.4000 58.2000 ;
	    RECT 67.0000 55.2000 67.3000 57.8000 ;
	    RECT 63.8000 54.7000 64.2000 55.1000 ;
	    RECT 67.0000 54.8000 67.4000 55.2000 ;
	    RECT 63.8000 54.2000 64.1000 54.7000 ;
	    RECT 63.8000 53.8000 64.2000 54.2000 ;
	    RECT 67.8000 52.1000 68.2000 57.9000 ;
	    RECT 71.0000 57.1000 71.4000 57.2000 ;
	    RECT 71.8000 57.1000 72.2000 57.2000 ;
	    RECT 71.0000 56.8000 72.2000 57.1000 ;
	    RECT 74.2000 57.1000 74.6000 57.2000 ;
	    RECT 75.0000 57.1000 75.4000 57.2000 ;
	    RECT 74.2000 56.8000 75.4000 57.1000 ;
	    RECT 79.0000 56.8000 79.4000 57.2000 ;
	    RECT 72.6000 54.8000 73.0000 55.2000 ;
	    RECT 75.8000 54.8000 76.2000 55.2000 ;
	    RECT 78.2000 54.8000 78.6000 55.2000 ;
	    RECT 70.2000 53.8000 70.6000 54.2000 ;
	    RECT 64.6000 49.8000 65.0000 50.2000 ;
	    RECT 61.4000 47.8000 61.8000 48.2000 ;
	    RECT 63.8000 47.8000 64.2000 48.2000 ;
	    RECT 61.4000 47.2000 61.7000 47.8000 ;
	    RECT 63.8000 47.2000 64.1000 47.8000 ;
	    RECT 61.4000 46.8000 61.8000 47.2000 ;
	    RECT 63.8000 46.8000 64.2000 47.2000 ;
	    RECT 58.2000 45.8000 58.6000 46.2000 ;
	    RECT 58.2000 45.2000 58.5000 45.8000 ;
	    RECT 58.2000 44.8000 58.6000 45.2000 ;
	    RECT 59.0000 44.8000 59.4000 45.2000 ;
	    RECT 60.6000 44.8000 61.0000 45.2000 ;
	    RECT 59.0000 44.2000 59.3000 44.8000 ;
	    RECT 60.6000 44.2000 60.9000 44.8000 ;
	    RECT 55.8000 42.8000 56.9000 43.1000 ;
	    RECT 57.4000 43.8000 57.8000 44.2000 ;
	    RECT 59.0000 43.8000 59.4000 44.2000 ;
	    RECT 60.6000 43.8000 61.0000 44.2000 ;
	    RECT 57.4000 43.2000 57.7000 43.8000 ;
	    RECT 57.4000 42.8000 57.8000 43.2000 ;
	    RECT 55.8000 39.2000 56.1000 42.8000 ;
	    RECT 55.8000 38.8000 56.2000 39.2000 ;
	    RECT 59.0000 38.2000 59.3000 43.8000 ;
	    RECT 64.6000 39.2000 64.9000 49.8000 ;
	    RECT 70.2000 49.2000 70.5000 53.8000 ;
	    RECT 72.6000 53.2000 72.9000 54.8000 ;
	    RECT 75.8000 54.2000 76.1000 54.8000 ;
	    RECT 78.2000 54.2000 78.5000 54.8000 ;
	    RECT 75.8000 53.8000 76.2000 54.2000 ;
	    RECT 78.2000 53.8000 78.6000 54.2000 ;
	    RECT 72.6000 52.8000 73.0000 53.2000 ;
	    RECT 79.0000 50.2000 79.3000 56.8000 ;
	    RECT 80.6000 53.1000 81.0000 55.9000 ;
	    RECT 82.2000 52.1000 82.6000 57.9000 ;
	    RECT 86.2000 56.8000 86.6000 57.2000 ;
	    RECT 83.0000 55.8000 83.4000 56.2000 ;
	    RECT 83.0000 55.1000 83.3000 55.8000 ;
	    RECT 86.2000 55.2000 86.5000 56.8000 ;
	    RECT 83.0000 54.7000 83.4000 55.1000 ;
	    RECT 86.2000 54.8000 86.6000 55.2000 ;
	    RECT 87.0000 52.1000 87.4000 57.9000 ;
	    RECT 88.6000 57.2000 88.9000 65.8000 ;
	    RECT 89.4000 59.2000 89.7000 66.8000 ;
	    RECT 90.2000 63.1000 90.6000 68.9000 ;
	    RECT 91.0000 68.2000 91.3000 74.8000 ;
	    RECT 102.2000 74.2000 102.5000 92.8000 ;
	    RECT 103.8000 91.8000 104.2000 92.2000 ;
	    RECT 103.8000 89.1000 104.1000 91.8000 ;
	    RECT 103.0000 83.1000 103.4000 88.9000 ;
	    RECT 103.8000 88.8000 104.9000 89.1000 ;
	    RECT 103.8000 87.8000 104.2000 88.2000 ;
	    RECT 103.8000 87.2000 104.1000 87.8000 ;
	    RECT 103.8000 86.8000 104.2000 87.2000 ;
	    RECT 103.8000 79.2000 104.1000 86.8000 ;
	    RECT 104.6000 86.2000 104.9000 88.8000 ;
	    RECT 104.6000 85.8000 105.0000 86.2000 ;
	    RECT 103.8000 78.8000 104.2000 79.2000 ;
	    RECT 97.4000 73.8000 97.8000 74.2000 ;
	    RECT 99.0000 73.8000 99.4000 74.2000 ;
	    RECT 100.6000 73.8000 101.0000 74.2000 ;
	    RECT 102.2000 73.8000 102.6000 74.2000 ;
	    RECT 97.4000 71.2000 97.7000 73.8000 ;
	    RECT 99.0000 73.2000 99.3000 73.8000 ;
	    RECT 99.0000 72.8000 99.4000 73.2000 ;
	    RECT 97.4000 70.8000 97.8000 71.2000 ;
	    RECT 95.0000 68.8000 95.4000 69.2000 ;
	    RECT 91.0000 67.8000 91.4000 68.2000 ;
	    RECT 93.4000 67.1000 93.8000 67.2000 ;
	    RECT 94.2000 67.1000 94.6000 67.2000 ;
	    RECT 93.4000 66.8000 94.6000 67.1000 ;
	    RECT 92.6000 66.1000 93.0000 66.2000 ;
	    RECT 93.4000 66.1000 93.8000 66.2000 ;
	    RECT 92.6000 65.8000 93.8000 66.1000 ;
	    RECT 89.4000 58.8000 89.8000 59.2000 ;
	    RECT 88.6000 56.8000 89.0000 57.2000 ;
	    RECT 90.2000 53.1000 90.6000 55.9000 ;
	    RECT 91.8000 52.1000 92.2000 57.9000 ;
	    RECT 95.0000 55.2000 95.3000 68.8000 ;
	    RECT 95.8000 67.8000 96.2000 68.2000 ;
	    RECT 96.6000 67.8000 97.0000 68.2000 ;
	    RECT 98.2000 67.8000 98.6000 68.2000 ;
	    RECT 95.8000 67.2000 96.1000 67.8000 ;
	    RECT 96.6000 67.2000 96.9000 67.8000 ;
	    RECT 98.2000 67.2000 98.5000 67.8000 ;
	    RECT 99.0000 67.2000 99.3000 72.8000 ;
	    RECT 100.6000 72.2000 100.9000 73.8000 ;
	    RECT 102.2000 73.1000 102.6000 73.2000 ;
	    RECT 103.0000 73.1000 103.4000 73.2000 ;
	    RECT 102.2000 72.8000 103.4000 73.1000 ;
	    RECT 100.6000 71.8000 101.0000 72.2000 ;
	    RECT 101.4000 71.8000 101.8000 72.2000 ;
	    RECT 101.4000 69.2000 101.7000 71.8000 ;
	    RECT 101.4000 68.8000 101.8000 69.2000 ;
	    RECT 95.8000 66.8000 96.2000 67.2000 ;
	    RECT 96.6000 66.8000 97.0000 67.2000 ;
	    RECT 97.4000 66.8000 97.8000 67.2000 ;
	    RECT 98.2000 66.8000 98.6000 67.2000 ;
	    RECT 99.0000 66.8000 99.4000 67.2000 ;
	    RECT 97.4000 66.2000 97.7000 66.8000 ;
	    RECT 95.8000 65.8000 96.2000 66.2000 ;
	    RECT 97.4000 65.8000 97.8000 66.2000 ;
	    RECT 99.0000 65.8000 99.4000 66.2000 ;
	    RECT 99.8000 66.1000 100.2000 66.2000 ;
	    RECT 100.6000 66.1000 101.0000 66.2000 ;
	    RECT 99.8000 65.8000 101.0000 66.1000 ;
	    RECT 95.8000 65.2000 96.1000 65.8000 ;
	    RECT 95.8000 64.8000 96.2000 65.2000 ;
	    RECT 99.0000 59.2000 99.3000 65.8000 ;
	    RECT 101.4000 65.1000 101.8000 67.9000 ;
	    RECT 102.2000 66.8000 102.6000 67.2000 ;
	    RECT 99.8000 63.8000 100.2000 64.2000 ;
	    RECT 99.8000 59.2000 100.1000 63.8000 ;
	    RECT 101.4000 62.8000 101.8000 63.2000 ;
	    RECT 99.0000 58.8000 99.4000 59.2000 ;
	    RECT 99.8000 58.8000 100.2000 59.2000 ;
	    RECT 95.8000 56.8000 96.2000 57.2000 ;
	    RECT 95.8000 55.2000 96.1000 56.8000 ;
	    RECT 95.0000 54.8000 95.4000 55.2000 ;
	    RECT 95.8000 54.8000 96.2000 55.2000 ;
	    RECT 96.6000 52.1000 97.0000 57.9000 ;
	    RECT 79.0000 49.8000 79.4000 50.2000 ;
	    RECT 101.4000 49.2000 101.7000 62.8000 ;
	    RECT 102.2000 59.2000 102.5000 66.8000 ;
	    RECT 103.0000 63.1000 103.4000 68.9000 ;
	    RECT 103.8000 66.2000 104.2000 66.3000 ;
	    RECT 104.6000 66.2000 105.0000 66.3000 ;
	    RECT 103.8000 65.9000 105.0000 66.2000 ;
	    RECT 102.2000 58.8000 102.6000 59.2000 ;
	    RECT 102.2000 57.2000 102.5000 58.8000 ;
	    RECT 102.2000 56.8000 102.6000 57.2000 ;
	    RECT 70.2000 48.8000 70.6000 49.2000 ;
	    RECT 101.4000 48.8000 101.8000 49.2000 ;
	    RECT 72.6000 47.8000 73.0000 48.2000 ;
	    RECT 78.2000 48.1000 78.6000 48.2000 ;
	    RECT 79.0000 48.1000 79.4000 48.2000 ;
	    RECT 78.2000 47.8000 79.4000 48.1000 ;
	    RECT 89.4000 47.8000 89.8000 48.2000 ;
	    RECT 66.2000 46.8000 66.6000 47.2000 ;
	    RECT 71.8000 46.8000 72.2000 47.2000 ;
	    RECT 66.2000 46.2000 66.5000 46.8000 ;
	    RECT 71.8000 46.2000 72.1000 46.8000 ;
	    RECT 66.2000 45.8000 66.6000 46.2000 ;
	    RECT 68.6000 46.1000 69.0000 46.2000 ;
	    RECT 67.8000 45.8000 69.0000 46.1000 ;
	    RECT 71.8000 45.8000 72.2000 46.2000 ;
	    RECT 67.8000 45.2000 68.1000 45.8000 ;
	    RECT 67.0000 44.8000 67.4000 45.2000 ;
	    RECT 67.8000 44.8000 68.2000 45.2000 ;
	    RECT 68.6000 44.8000 69.0000 45.2000 ;
	    RECT 67.0000 44.2000 67.3000 44.8000 ;
	    RECT 65.4000 43.8000 65.8000 44.2000 ;
	    RECT 67.0000 43.8000 67.4000 44.2000 ;
	    RECT 65.4000 43.2000 65.7000 43.8000 ;
	    RECT 65.4000 42.8000 65.8000 43.2000 ;
	    RECT 66.2000 41.8000 66.6000 42.2000 ;
	    RECT 64.6000 38.8000 65.0000 39.2000 ;
	    RECT 59.0000 37.8000 59.4000 38.2000 ;
	    RECT 65.4000 37.8000 65.8000 38.2000 ;
	    RECT 55.0000 36.8000 55.4000 37.2000 ;
	    RECT 63.8000 36.8000 64.2000 37.2000 ;
	    RECT 53.4000 35.8000 53.8000 36.2000 ;
	    RECT 53.4000 34.2000 53.7000 35.8000 ;
	    RECT 53.4000 33.8000 53.8000 34.2000 ;
	    RECT 53.4000 32.2000 53.7000 33.8000 ;
	    RECT 55.0000 33.2000 55.3000 36.8000 ;
	    RECT 55.8000 36.1000 56.2000 36.2000 ;
	    RECT 56.6000 36.1000 57.0000 36.2000 ;
	    RECT 55.8000 35.8000 57.0000 36.1000 ;
	    RECT 57.4000 35.8000 57.8000 36.2000 ;
	    RECT 62.2000 36.1000 62.6000 36.2000 ;
	    RECT 63.0000 36.1000 63.4000 36.2000 ;
	    RECT 62.2000 35.8000 63.4000 36.1000 ;
	    RECT 55.8000 34.8000 56.2000 35.2000 ;
	    RECT 56.6000 34.8000 57.0000 35.2000 ;
	    RECT 55.8000 34.2000 56.1000 34.8000 ;
	    RECT 55.8000 33.8000 56.2000 34.2000 ;
	    RECT 55.0000 32.8000 55.4000 33.2000 ;
	    RECT 53.4000 31.8000 53.8000 32.2000 ;
	    RECT 56.6000 29.2000 56.9000 34.8000 ;
	    RECT 57.4000 34.2000 57.7000 35.8000 ;
	    RECT 57.4000 33.8000 57.8000 34.2000 ;
	    RECT 57.4000 33.1000 57.8000 33.2000 ;
	    RECT 58.2000 33.1000 58.6000 33.2000 ;
	    RECT 57.4000 32.8000 58.6000 33.1000 ;
	    RECT 59.0000 31.8000 59.4000 32.2000 ;
	    RECT 59.0000 29.2000 59.3000 31.8000 ;
	    RECT 63.8000 29.2000 64.1000 36.8000 ;
	    RECT 65.4000 36.2000 65.7000 37.8000 ;
	    RECT 66.2000 36.2000 66.5000 41.8000 ;
	    RECT 67.0000 41.2000 67.3000 43.8000 ;
	    RECT 67.8000 42.8000 68.2000 43.2000 ;
	    RECT 67.0000 40.8000 67.4000 41.2000 ;
	    RECT 67.8000 39.2000 68.1000 42.8000 ;
	    RECT 67.8000 38.8000 68.2000 39.2000 ;
	    RECT 68.6000 38.2000 68.9000 44.8000 ;
	    RECT 72.6000 44.2000 72.9000 47.8000 ;
	    RECT 89.4000 47.2000 89.7000 47.8000 ;
	    RECT 74.2000 47.1000 74.6000 47.2000 ;
	    RECT 75.0000 47.1000 75.4000 47.2000 ;
	    RECT 74.2000 46.8000 75.4000 47.1000 ;
	    RECT 77.4000 46.8000 77.8000 47.2000 ;
	    RECT 82.2000 47.1000 82.6000 47.2000 ;
	    RECT 83.0000 47.1000 83.4000 47.2000 ;
	    RECT 82.2000 46.8000 83.4000 47.1000 ;
	    RECT 89.4000 46.8000 89.8000 47.2000 ;
	    RECT 91.8000 46.8000 92.2000 47.2000 ;
	    RECT 96.6000 46.8000 97.0000 47.2000 ;
	    RECT 102.2000 46.8000 102.6000 47.2000 ;
	    RECT 104.6000 46.8000 105.0000 47.2000 ;
	    RECT 69.4000 44.1000 69.8000 44.2000 ;
	    RECT 70.2000 44.1000 70.6000 44.2000 ;
	    RECT 69.4000 43.8000 70.6000 44.1000 ;
	    RECT 72.6000 43.8000 73.0000 44.2000 ;
	    RECT 74.2000 42.8000 74.6000 43.2000 ;
	    RECT 71.8000 41.8000 72.2000 42.2000 ;
	    RECT 71.8000 39.1000 72.1000 41.8000 ;
	    RECT 71.0000 38.8000 72.1000 39.1000 ;
	    RECT 74.2000 39.2000 74.5000 42.8000 ;
	    RECT 74.2000 38.8000 74.6000 39.2000 ;
	    RECT 68.6000 37.8000 69.0000 38.2000 ;
	    RECT 67.0000 36.8000 67.4000 37.2000 ;
	    RECT 64.6000 36.1000 65.0000 36.2000 ;
	    RECT 65.4000 36.1000 65.8000 36.2000 ;
	    RECT 64.6000 35.8000 65.8000 36.1000 ;
	    RECT 66.2000 35.8000 66.6000 36.2000 ;
	    RECT 64.6000 34.8000 65.0000 35.2000 ;
	    RECT 67.0000 35.1000 67.3000 36.8000 ;
	    RECT 68.6000 36.2000 68.9000 37.8000 ;
	    RECT 71.0000 37.2000 71.3000 38.8000 ;
	    RECT 71.8000 38.1000 72.2000 38.2000 ;
	    RECT 72.6000 38.1000 73.0000 38.2000 ;
	    RECT 71.8000 37.8000 73.0000 38.1000 ;
	    RECT 71.0000 36.8000 71.4000 37.2000 ;
	    RECT 73.4000 36.8000 73.8000 37.2000 ;
	    RECT 68.6000 35.8000 69.0000 36.2000 ;
	    RECT 70.2000 35.8000 70.6000 36.2000 ;
	    RECT 70.2000 35.2000 70.5000 35.8000 ;
	    RECT 66.2000 34.8000 67.3000 35.1000 ;
	    RECT 67.8000 34.8000 68.2000 35.2000 ;
	    RECT 70.2000 34.8000 70.6000 35.2000 ;
	    RECT 64.6000 34.2000 64.9000 34.8000 ;
	    RECT 64.6000 33.8000 65.0000 34.2000 ;
	    RECT 66.2000 29.2000 66.5000 34.8000 ;
	    RECT 67.8000 33.2000 68.1000 34.8000 ;
	    RECT 73.4000 34.2000 73.7000 36.8000 ;
	    RECT 75.8000 36.1000 76.2000 36.2000 ;
	    RECT 76.6000 36.1000 77.0000 36.2000 ;
	    RECT 75.8000 35.8000 77.0000 36.1000 ;
	    RECT 77.4000 35.2000 77.7000 46.8000 ;
	    RECT 91.8000 46.2000 92.1000 46.8000 ;
	    RECT 85.4000 46.1000 85.8000 46.2000 ;
	    RECT 87.0000 46.1000 87.4000 46.2000 ;
	    RECT 85.4000 45.8000 87.4000 46.1000 ;
	    RECT 91.8000 45.8000 92.2000 46.2000 ;
	    RECT 93.4000 45.8000 93.8000 46.2000 ;
	    RECT 93.4000 45.2000 93.7000 45.8000 ;
	    RECT 90.2000 44.8000 90.6000 45.2000 ;
	    RECT 91.8000 45.1000 92.2000 45.2000 ;
	    RECT 92.6000 45.1000 93.0000 45.2000 ;
	    RECT 91.8000 44.8000 93.0000 45.1000 ;
	    RECT 93.4000 44.8000 93.8000 45.2000 ;
	    RECT 90.2000 44.2000 90.5000 44.8000 ;
	    RECT 96.6000 44.2000 96.9000 46.8000 ;
	    RECT 102.2000 46.2000 102.5000 46.8000 ;
	    RECT 104.6000 46.2000 104.9000 46.8000 ;
	    RECT 97.4000 45.8000 97.8000 46.2000 ;
	    RECT 99.8000 46.1000 100.2000 46.2000 ;
	    RECT 100.6000 46.1000 101.0000 46.2000 ;
	    RECT 99.8000 45.8000 101.0000 46.1000 ;
	    RECT 101.4000 45.8000 101.8000 46.2000 ;
	    RECT 102.2000 45.8000 102.6000 46.2000 ;
	    RECT 104.6000 45.8000 105.0000 46.2000 ;
	    RECT 97.4000 44.2000 97.7000 45.8000 ;
	    RECT 98.2000 44.8000 98.6000 45.2000 ;
	    RECT 84.6000 43.8000 85.0000 44.2000 ;
	    RECT 85.4000 44.1000 85.8000 44.2000 ;
	    RECT 86.2000 44.1000 86.6000 44.2000 ;
	    RECT 85.4000 43.8000 86.6000 44.1000 ;
	    RECT 90.2000 43.8000 90.6000 44.2000 ;
	    RECT 95.8000 43.8000 96.2000 44.2000 ;
	    RECT 96.6000 43.8000 97.0000 44.2000 ;
	    RECT 97.4000 43.8000 97.8000 44.2000 ;
	    RECT 84.6000 43.2000 84.9000 43.8000 ;
	    RECT 84.6000 42.8000 85.0000 43.2000 ;
	    RECT 82.2000 41.8000 82.6000 42.2000 ;
	    RECT 81.4000 40.8000 81.8000 41.2000 ;
	    RECT 81.4000 39.2000 81.7000 40.8000 ;
	    RECT 81.4000 38.8000 81.8000 39.2000 ;
	    RECT 82.2000 36.2000 82.5000 41.8000 ;
	    RECT 89.4000 40.8000 89.8000 41.2000 ;
	    RECT 95.0000 40.8000 95.4000 41.2000 ;
	    RECT 89.4000 39.2000 89.7000 40.8000 ;
	    RECT 91.0000 39.8000 91.4000 40.2000 ;
	    RECT 89.4000 38.8000 89.8000 39.2000 ;
	    RECT 85.4000 38.1000 85.8000 38.2000 ;
	    RECT 86.2000 38.1000 86.6000 38.2000 ;
	    RECT 85.4000 37.8000 86.6000 38.1000 ;
	    RECT 88.6000 36.8000 89.0000 37.2000 ;
	    RECT 88.6000 36.2000 88.9000 36.8000 ;
	    RECT 82.2000 35.8000 82.6000 36.2000 ;
	    RECT 88.6000 35.8000 89.0000 36.2000 ;
	    RECT 89.4000 36.1000 89.8000 36.2000 ;
	    RECT 90.2000 36.1000 90.6000 36.2000 ;
	    RECT 89.4000 35.8000 90.6000 36.1000 ;
	    RECT 74.2000 34.8000 74.6000 35.2000 ;
	    RECT 75.8000 35.1000 76.2000 35.2000 ;
	    RECT 76.6000 35.1000 77.0000 35.2000 ;
	    RECT 75.8000 34.8000 77.0000 35.1000 ;
	    RECT 77.4000 35.1000 77.8000 35.2000 ;
	    RECT 77.4000 34.8000 79.3000 35.1000 ;
	    RECT 73.4000 33.8000 73.8000 34.2000 ;
	    RECT 67.8000 32.8000 68.2000 33.2000 ;
	    RECT 74.2000 32.2000 74.5000 34.8000 ;
	    RECT 76.6000 33.8000 77.0000 34.2000 ;
	    RECT 75.0000 32.8000 75.4000 33.2000 ;
	    RECT 74.2000 31.8000 74.6000 32.2000 ;
	    RECT 75.0000 29.2000 75.3000 32.8000 ;
	    RECT 76.6000 29.2000 76.9000 33.8000 ;
	    RECT 79.0000 29.2000 79.3000 34.8000 ;
	    RECT 82.2000 34.8000 82.6000 35.2000 ;
	    RECT 81.4000 31.8000 81.8000 32.2000 ;
	    RECT 56.6000 28.8000 57.0000 29.2000 ;
	    RECT 59.0000 28.8000 59.4000 29.2000 ;
	    RECT 63.8000 28.8000 64.2000 29.2000 ;
	    RECT 66.2000 28.8000 66.6000 29.2000 ;
	    RECT 67.8000 28.8000 68.2000 29.2000 ;
	    RECT 75.0000 28.8000 75.4000 29.2000 ;
	    RECT 75.8000 28.8000 76.2000 29.2000 ;
	    RECT 76.6000 28.8000 77.0000 29.2000 ;
	    RECT 79.0000 28.8000 79.4000 29.2000 ;
	    RECT 67.8000 28.2000 68.1000 28.8000 ;
	    RECT 63.8000 27.8000 64.2000 28.2000 ;
	    RECT 67.8000 27.8000 68.2000 28.2000 ;
	    RECT 69.4000 28.1000 69.8000 28.2000 ;
	    RECT 70.2000 28.1000 70.6000 28.2000 ;
	    RECT 69.4000 27.8000 70.6000 28.1000 ;
	    RECT 73.4000 27.8000 73.8000 28.2000 ;
	    RECT 51.8000 26.1000 52.2000 26.2000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 51.8000 25.8000 53.0000 26.1000 ;
	    RECT 53.4000 26.1000 53.8000 26.2000 ;
	    RECT 54.2000 26.1000 54.6000 26.2000 ;
	    RECT 53.4000 25.8000 54.6000 26.1000 ;
	    RECT 56.6000 26.1000 57.0000 26.2000 ;
	    RECT 57.4000 26.1000 57.8000 26.2000 ;
	    RECT 56.6000 25.8000 57.8000 26.1000 ;
	    RECT 53.4000 24.8000 53.8000 25.2000 ;
	    RECT 57.4000 24.8000 57.8000 25.2000 ;
	    RECT 60.6000 25.1000 61.0000 25.2000 ;
	    RECT 61.4000 25.1000 61.8000 25.2000 ;
	    RECT 60.6000 24.8000 61.8000 25.1000 ;
	    RECT 53.4000 24.2000 53.7000 24.8000 ;
	    RECT 53.4000 23.8000 53.8000 24.2000 ;
	    RECT 54.2000 23.8000 54.6000 24.2000 ;
	    RECT 56.6000 23.8000 57.0000 24.2000 ;
	    RECT 54.2000 23.2000 54.5000 23.8000 ;
	    RECT 56.6000 23.2000 56.9000 23.8000 ;
	    RECT 54.2000 22.8000 54.6000 23.2000 ;
	    RECT 56.6000 22.8000 57.0000 23.2000 ;
	    RECT 57.4000 19.2000 57.7000 24.8000 ;
	    RECT 57.4000 18.8000 57.8000 19.2000 ;
	    RECT 63.8000 17.2000 64.1000 27.8000 ;
	    RECT 73.4000 25.2000 73.7000 27.8000 ;
	    RECT 74.2000 25.8000 74.6000 26.2000 ;
	    RECT 65.4000 24.8000 65.8000 25.2000 ;
	    RECT 67.0000 24.8000 67.4000 25.2000 ;
	    RECT 73.4000 24.8000 73.8000 25.2000 ;
	    RECT 58.2000 16.8000 58.6000 17.2000 ;
	    RECT 63.8000 16.8000 64.2000 17.2000 ;
	    RECT 64.6000 16.8000 65.0000 17.2000 ;
	    RECT 51.0000 15.8000 51.4000 16.2000 ;
	    RECT 55.8000 15.8000 56.2000 16.2000 ;
	    RECT 51.0000 15.1000 51.4000 15.2000 ;
	    RECT 51.8000 15.1000 52.2000 15.2000 ;
	    RECT 51.0000 14.8000 52.2000 15.1000 ;
	    RECT 52.6000 14.8000 53.0000 15.2000 ;
	    RECT 52.6000 14.2000 52.9000 14.8000 ;
	    RECT 47.8000 13.8000 48.2000 14.2000 ;
	    RECT 50.2000 13.8000 50.6000 14.2000 ;
	    RECT 51.8000 13.8000 52.2000 14.2000 ;
	    RECT 52.6000 13.8000 53.0000 14.2000 ;
	    RECT 51.8000 9.2000 52.1000 13.8000 ;
	    RECT 55.0000 12.8000 55.4000 13.2000 ;
	    RECT 47.0000 8.8000 47.4000 9.2000 ;
	    RECT 51.8000 8.8000 52.2000 9.2000 ;
	    RECT 55.0000 8.2000 55.3000 12.8000 ;
	    RECT 55.8000 9.2000 56.1000 15.8000 ;
	    RECT 58.2000 15.2000 58.5000 16.8000 ;
	    RECT 63.8000 15.2000 64.1000 16.8000 ;
	    RECT 57.4000 14.8000 57.8000 15.2000 ;
	    RECT 58.2000 14.8000 58.6000 15.2000 ;
	    RECT 63.8000 14.8000 64.2000 15.2000 ;
	    RECT 57.4000 9.2000 57.7000 14.8000 ;
	    RECT 64.6000 9.2000 64.9000 16.8000 ;
	    RECT 65.4000 15.2000 65.7000 24.8000 ;
	    RECT 67.0000 19.2000 67.3000 24.8000 ;
	    RECT 73.4000 21.2000 73.7000 24.8000 ;
	    RECT 74.2000 24.2000 74.5000 25.8000 ;
	    RECT 74.2000 23.8000 74.6000 24.2000 ;
	    RECT 75.0000 23.8000 75.4000 24.2000 ;
	    RECT 75.0000 23.1000 75.3000 23.8000 ;
	    RECT 74.2000 22.8000 75.3000 23.1000 ;
	    RECT 69.4000 20.8000 69.8000 21.2000 ;
	    RECT 73.4000 20.8000 73.8000 21.2000 ;
	    RECT 67.0000 18.8000 67.4000 19.2000 ;
	    RECT 67.0000 17.1000 67.4000 17.2000 ;
	    RECT 67.8000 17.1000 68.2000 17.2000 ;
	    RECT 67.0000 16.8000 68.2000 17.1000 ;
	    RECT 68.6000 16.8000 69.0000 17.2000 ;
	    RECT 66.2000 15.8000 66.6000 16.2000 ;
	    RECT 66.2000 15.2000 66.5000 15.8000 ;
	    RECT 68.6000 15.2000 68.9000 16.8000 ;
	    RECT 69.4000 16.2000 69.7000 20.8000 ;
	    RECT 73.4000 17.2000 73.7000 20.8000 ;
	    RECT 72.6000 16.8000 73.0000 17.2000 ;
	    RECT 73.4000 16.8000 73.8000 17.2000 ;
	    RECT 72.6000 16.2000 72.9000 16.8000 ;
	    RECT 69.4000 15.8000 69.8000 16.2000 ;
	    RECT 72.6000 15.8000 73.0000 16.2000 ;
	    RECT 73.4000 15.8000 73.8000 16.2000 ;
	    RECT 73.4000 15.2000 73.7000 15.8000 ;
	    RECT 65.4000 14.8000 65.8000 15.2000 ;
	    RECT 66.2000 14.8000 66.6000 15.2000 ;
	    RECT 68.6000 14.8000 69.0000 15.2000 ;
	    RECT 69.4000 14.8000 69.8000 15.2000 ;
	    RECT 73.4000 14.8000 73.8000 15.2000 ;
	    RECT 67.0000 10.8000 67.4000 11.2000 ;
	    RECT 67.0000 9.2000 67.3000 10.8000 ;
	    RECT 69.4000 9.2000 69.7000 14.8000 ;
	    RECT 74.2000 13.2000 74.5000 22.8000 ;
	    RECT 75.0000 21.8000 75.4000 22.2000 ;
	    RECT 75.0000 19.2000 75.3000 21.8000 ;
	    RECT 75.0000 18.8000 75.4000 19.2000 ;
	    RECT 75.8000 15.2000 76.1000 28.8000 ;
	    RECT 81.4000 28.2000 81.7000 31.8000 ;
	    RECT 82.2000 29.2000 82.5000 34.8000 ;
	    RECT 91.0000 34.2000 91.3000 39.8000 ;
	    RECT 95.0000 37.2000 95.3000 40.8000 ;
	    RECT 95.8000 39.2000 96.1000 43.8000 ;
	    RECT 95.8000 38.8000 96.2000 39.2000 ;
	    RECT 98.2000 38.2000 98.5000 44.8000 ;
	    RECT 97.4000 37.8000 97.8000 38.2000 ;
	    RECT 98.2000 37.8000 98.6000 38.2000 ;
	    RECT 95.0000 36.8000 95.4000 37.2000 ;
	    RECT 97.4000 37.1000 97.7000 37.8000 ;
	    RECT 98.2000 37.1000 98.6000 37.2000 ;
	    RECT 97.4000 36.8000 98.6000 37.1000 ;
	    RECT 93.4000 35.8000 93.8000 36.2000 ;
	    RECT 96.6000 36.1000 97.0000 36.2000 ;
	    RECT 97.4000 36.1000 97.8000 36.2000 ;
	    RECT 96.6000 35.8000 97.8000 36.1000 ;
	    RECT 99.8000 35.8000 100.2000 36.2000 ;
	    RECT 100.6000 35.8000 101.0000 36.2000 ;
	    RECT 93.4000 35.2000 93.7000 35.8000 ;
	    RECT 93.4000 34.8000 93.8000 35.2000 ;
	    RECT 95.0000 35.1000 95.4000 35.2000 ;
	    RECT 95.8000 35.1000 96.2000 35.2000 ;
	    RECT 95.0000 34.8000 96.2000 35.1000 ;
	    RECT 99.0000 34.8000 99.4000 35.2000 ;
	    RECT 99.0000 34.2000 99.3000 34.8000 ;
	    RECT 86.2000 34.1000 86.6000 34.2000 ;
	    RECT 87.0000 34.1000 87.4000 34.2000 ;
	    RECT 86.2000 33.8000 87.4000 34.1000 ;
	    RECT 88.6000 34.1000 89.0000 34.2000 ;
	    RECT 89.4000 34.1000 89.8000 34.2000 ;
	    RECT 88.6000 33.8000 89.8000 34.1000 ;
	    RECT 91.0000 33.8000 91.4000 34.2000 ;
	    RECT 97.4000 34.1000 97.8000 34.2000 ;
	    RECT 98.2000 34.1000 98.6000 34.2000 ;
	    RECT 97.4000 33.8000 98.6000 34.1000 ;
	    RECT 99.0000 33.8000 99.4000 34.2000 ;
	    RECT 91.0000 33.2000 91.3000 33.8000 ;
	    RECT 91.0000 32.8000 91.4000 33.2000 ;
	    RECT 91.0000 31.8000 91.4000 32.2000 ;
	    RECT 91.0000 30.1000 91.3000 31.8000 ;
	    RECT 98.2000 30.8000 98.6000 31.2000 ;
	    RECT 91.0000 29.8000 92.1000 30.1000 ;
	    RECT 82.2000 28.8000 82.6000 29.2000 ;
	    RECT 81.4000 27.8000 81.8000 28.2000 ;
	    RECT 84.6000 28.1000 85.0000 28.2000 ;
	    RECT 85.4000 28.1000 85.8000 28.2000 ;
	    RECT 84.6000 27.8000 85.8000 28.1000 ;
	    RECT 89.4000 27.8000 89.8000 28.2000 ;
	    RECT 89.4000 27.2000 89.7000 27.8000 ;
	    RECT 88.6000 26.8000 89.0000 27.2000 ;
	    RECT 89.4000 26.8000 89.8000 27.2000 ;
	    RECT 88.6000 26.2000 88.9000 26.8000 ;
	    RECT 82.2000 25.8000 82.6000 26.2000 ;
	    RECT 87.0000 25.8000 87.4000 26.2000 ;
	    RECT 88.6000 25.8000 89.0000 26.2000 ;
	    RECT 76.6000 24.8000 77.0000 25.2000 ;
	    RECT 76.6000 22.2000 76.9000 24.8000 ;
	    RECT 76.6000 21.8000 77.0000 22.2000 ;
	    RECT 82.2000 19.2000 82.5000 25.8000 ;
	    RECT 87.0000 25.2000 87.3000 25.8000 ;
	    RECT 87.0000 24.8000 87.4000 25.2000 ;
	    RECT 83.0000 23.8000 83.4000 24.2000 ;
	    RECT 83.0000 22.2000 83.3000 23.8000 ;
	    RECT 83.0000 21.8000 83.4000 22.2000 ;
	    RECT 85.4000 21.8000 85.8000 22.2000 ;
	    RECT 85.4000 19.2000 85.7000 21.8000 ;
	    RECT 82.2000 18.8000 82.6000 19.2000 ;
	    RECT 85.4000 18.8000 85.8000 19.2000 ;
	    RECT 81.4000 16.8000 81.8000 17.2000 ;
	    RECT 83.0000 16.8000 83.4000 17.2000 ;
	    RECT 83.8000 16.8000 84.2000 17.2000 ;
	    RECT 85.4000 17.1000 85.8000 17.2000 ;
	    RECT 86.2000 17.1000 86.6000 17.2000 ;
	    RECT 85.4000 16.8000 86.6000 17.1000 ;
	    RECT 87.8000 16.8000 88.2000 17.2000 ;
	    RECT 81.4000 16.2000 81.7000 16.8000 ;
	    RECT 80.6000 15.8000 81.0000 16.2000 ;
	    RECT 81.4000 15.8000 81.8000 16.2000 ;
	    RECT 82.2000 15.8000 82.6000 16.2000 ;
	    RECT 80.6000 15.2000 80.9000 15.8000 ;
	    RECT 81.4000 15.2000 81.7000 15.8000 ;
	    RECT 82.2000 15.2000 82.5000 15.8000 ;
	    RECT 75.8000 14.8000 76.2000 15.2000 ;
	    RECT 78.2000 14.8000 78.6000 15.2000 ;
	    RECT 80.6000 14.8000 81.0000 15.2000 ;
	    RECT 81.4000 14.8000 81.8000 15.2000 ;
	    RECT 82.2000 14.8000 82.6000 15.2000 ;
	    RECT 78.2000 13.2000 78.5000 14.8000 ;
	    RECT 70.2000 12.8000 70.6000 13.2000 ;
	    RECT 74.2000 12.8000 74.6000 13.2000 ;
	    RECT 75.8000 12.8000 76.2000 13.2000 ;
	    RECT 78.2000 12.8000 78.6000 13.2000 ;
	    RECT 55.8000 8.8000 56.2000 9.2000 ;
	    RECT 57.4000 8.8000 57.8000 9.2000 ;
	    RECT 64.6000 8.8000 65.0000 9.2000 ;
	    RECT 67.0000 8.8000 67.4000 9.2000 ;
	    RECT 69.4000 8.8000 69.8000 9.2000 ;
	    RECT 70.2000 8.2000 70.5000 12.8000 ;
	    RECT 72.6000 11.8000 73.0000 12.2000 ;
	    RECT 72.6000 9.2000 72.9000 11.8000 ;
	    RECT 75.8000 9.2000 76.1000 12.8000 ;
	    RECT 83.0000 12.2000 83.3000 16.8000 ;
	    RECT 83.0000 11.8000 83.4000 12.2000 ;
	    RECT 83.8000 9.2000 84.1000 16.8000 ;
	    RECT 87.8000 16.2000 88.1000 16.8000 ;
	    RECT 85.4000 15.8000 85.8000 16.2000 ;
	    RECT 87.8000 15.8000 88.2000 16.2000 ;
	    RECT 85.4000 15.2000 85.7000 15.8000 ;
	    RECT 85.4000 14.8000 85.8000 15.2000 ;
	    RECT 89.4000 15.1000 89.7000 26.8000 ;
	    RECT 90.2000 22.1000 90.6000 22.2000 ;
	    RECT 91.0000 22.1000 91.4000 22.2000 ;
	    RECT 90.2000 21.8000 91.4000 22.1000 ;
	    RECT 91.8000 19.2000 92.1000 29.8000 ;
	    RECT 98.2000 29.2000 98.5000 30.8000 ;
	    RECT 99.8000 29.2000 100.1000 35.8000 ;
	    RECT 100.6000 35.2000 100.9000 35.8000 ;
	    RECT 100.6000 34.8000 101.0000 35.2000 ;
	    RECT 101.4000 29.2000 101.7000 45.8000 ;
	    RECT 102.2000 44.8000 102.6000 45.2000 ;
	    RECT 102.2000 44.2000 102.5000 44.8000 ;
	    RECT 102.2000 43.8000 102.6000 44.2000 ;
	    RECT 104.6000 40.2000 104.9000 45.8000 ;
	    RECT 106.2000 40.8000 106.6000 41.2000 ;
	    RECT 104.6000 39.8000 105.0000 40.2000 ;
	    RECT 104.6000 36.2000 104.9000 39.8000 ;
	    RECT 106.2000 37.2000 106.5000 40.8000 ;
	    RECT 107.0000 39.2000 107.3000 93.8000 ;
	    RECT 108.6000 93.1000 109.0000 93.2000 ;
	    RECT 109.4000 93.1000 109.8000 93.2000 ;
	    RECT 108.6000 92.8000 109.8000 93.1000 ;
	    RECT 113.4000 92.8000 113.8000 93.2000 ;
	    RECT 111.0000 92.1000 111.4000 92.2000 ;
	    RECT 111.8000 92.1000 112.2000 92.2000 ;
	    RECT 111.0000 91.8000 112.2000 92.1000 ;
	    RECT 112.6000 89.1000 113.0000 89.2000 ;
	    RECT 113.4000 89.1000 113.7000 92.8000 ;
	    RECT 107.8000 83.1000 108.2000 88.9000 ;
	    RECT 112.6000 88.8000 113.7000 89.1000 ;
	    RECT 113.4000 87.1000 113.8000 87.2000 ;
	    RECT 114.2000 87.1000 114.6000 87.2000 ;
	    RECT 113.4000 86.8000 114.6000 87.1000 ;
	    RECT 111.0000 86.1000 111.4000 86.2000 ;
	    RECT 111.8000 86.1000 112.2000 86.2000 ;
	    RECT 111.0000 85.8000 112.2000 86.1000 ;
	    RECT 111.0000 81.8000 111.4000 82.2000 ;
	    RECT 111.0000 73.2000 111.3000 81.8000 ;
	    RECT 111.0000 72.8000 111.4000 73.2000 ;
	    RECT 114.2000 73.1000 114.6000 75.9000 ;
	    RECT 110.2000 71.8000 110.6000 72.2000 ;
	    RECT 107.8000 63.1000 108.2000 68.9000 ;
	    RECT 110.2000 68.2000 110.5000 71.8000 ;
	    RECT 111.0000 69.1000 111.4000 69.2000 ;
	    RECT 111.8000 69.1000 112.2000 69.2000 ;
	    RECT 111.0000 68.8000 112.2000 69.1000 ;
	    RECT 110.2000 67.8000 110.6000 68.2000 ;
	    RECT 115.0000 67.2000 115.3000 93.8000 ;
	    RECT 115.8000 93.1000 116.2000 93.2000 ;
	    RECT 116.6000 93.1000 117.0000 93.2000 ;
	    RECT 117.4000 93.1000 117.8000 95.9000 ;
	    RECT 118.2000 93.8000 118.6000 94.2000 ;
	    RECT 115.8000 92.8000 117.0000 93.1000 ;
	    RECT 118.2000 92.1000 118.5000 93.8000 ;
	    RECT 119.0000 92.1000 119.4000 97.9000 ;
	    RECT 119.8000 95.0000 120.2000 95.1000 ;
	    RECT 120.6000 95.0000 121.0000 95.1000 ;
	    RECT 119.8000 94.7000 121.0000 95.0000 ;
	    RECT 117.4000 91.8000 118.5000 92.1000 ;
	    RECT 116.6000 90.8000 117.0000 91.2000 ;
	    RECT 116.6000 89.2000 116.9000 90.8000 ;
	    RECT 116.6000 88.8000 117.0000 89.2000 ;
	    RECT 117.4000 88.2000 117.7000 91.8000 ;
	    RECT 118.2000 88.8000 118.6000 89.2000 ;
	    RECT 119.0000 89.1000 119.4000 89.2000 ;
	    RECT 119.8000 89.1000 120.2000 89.2000 ;
	    RECT 119.0000 88.8000 120.2000 89.1000 ;
	    RECT 117.4000 87.8000 117.8000 88.2000 ;
	    RECT 118.2000 87.0000 118.5000 88.8000 ;
	    RECT 119.0000 87.1000 119.4000 87.2000 ;
	    RECT 119.8000 87.1000 120.2000 87.2000 ;
	    RECT 118.2000 86.6000 118.6000 87.0000 ;
	    RECT 119.0000 86.8000 120.2000 87.1000 ;
	    RECT 122.2000 83.1000 122.6000 88.9000 ;
	    RECT 123.0000 87.2000 123.3000 106.8000 ;
	    RECT 123.8000 102.2000 124.1000 106.8000 ;
	    RECT 124.6000 106.2000 124.9000 114.8000 ;
	    RECT 127.0000 113.8000 127.4000 114.2000 ;
	    RECT 126.2000 112.8000 126.6000 113.2000 ;
	    RECT 125.4000 111.8000 125.8000 112.2000 ;
	    RECT 125.4000 106.2000 125.7000 111.8000 ;
	    RECT 124.6000 105.8000 125.0000 106.2000 ;
	    RECT 125.4000 105.8000 125.8000 106.2000 ;
	    RECT 123.8000 101.8000 124.2000 102.2000 ;
	    RECT 124.6000 101.2000 124.9000 105.8000 ;
	    RECT 126.2000 102.2000 126.5000 112.8000 ;
	    RECT 127.0000 112.2000 127.3000 113.8000 ;
	    RECT 129.4000 112.2000 129.7000 114.8000 ;
	    RECT 132.6000 113.8000 133.0000 114.2000 ;
	    RECT 131.8000 112.8000 132.2000 113.2000 ;
	    RECT 131.8000 112.2000 132.1000 112.8000 ;
	    RECT 127.0000 111.8000 127.4000 112.2000 ;
	    RECT 129.4000 111.8000 129.8000 112.2000 ;
	    RECT 131.8000 111.8000 132.2000 112.2000 ;
	    RECT 127.8000 107.8000 128.2000 108.2000 ;
	    RECT 127.8000 106.2000 128.1000 107.8000 ;
	    RECT 129.4000 107.1000 129.7000 111.8000 ;
	    RECT 130.2000 108.1000 130.6000 108.2000 ;
	    RECT 131.0000 108.1000 131.4000 108.2000 ;
	    RECT 130.2000 107.8000 131.4000 108.1000 ;
	    RECT 130.2000 107.1000 130.6000 107.2000 ;
	    RECT 129.4000 106.8000 130.6000 107.1000 ;
	    RECT 132.6000 106.2000 132.9000 113.8000 ;
	    RECT 134.2000 109.2000 134.5000 122.8000 ;
	    RECT 137.4000 122.2000 137.7000 127.8000 ;
	    RECT 138.2000 127.2000 138.5000 128.8000 ;
	    RECT 141.4000 127.2000 141.7000 128.8000 ;
	    RECT 144.6000 128.2000 144.9000 134.8000 ;
	    RECT 147.0000 134.1000 147.3000 136.8000 ;
	    RECT 147.8000 135.2000 148.1000 139.8000 ;
	    RECT 150.2000 137.2000 150.5000 145.8000 ;
	    RECT 151.0000 144.2000 151.3000 147.8000 ;
	    RECT 154.2000 146.2000 154.5000 150.8000 ;
	    RECT 155.0000 147.2000 155.3000 152.8000 ;
	    RECT 156.6000 147.2000 156.9000 153.8000 ;
	    RECT 157.4000 149.2000 157.7000 154.8000 ;
	    RECT 159.8000 153.8000 160.2000 154.2000 ;
	    RECT 159.8000 151.2000 160.1000 153.8000 ;
	    RECT 161.4000 153.2000 161.7000 155.8000 ;
	    RECT 161.4000 152.8000 161.8000 153.2000 ;
	    RECT 162.2000 153.1000 162.6000 155.9000 ;
	    RECT 160.6000 151.8000 161.0000 152.2000 ;
	    RECT 161.4000 151.8000 161.8000 152.2000 ;
	    RECT 163.8000 152.1000 164.2000 157.9000 ;
	    RECT 164.6000 154.7000 165.0000 155.1000 ;
	    RECT 164.6000 154.2000 164.9000 154.7000 ;
	    RECT 164.6000 153.8000 165.0000 154.2000 ;
	    RECT 165.4000 153.8000 165.8000 154.2000 ;
	    RECT 159.8000 150.8000 160.2000 151.2000 ;
	    RECT 160.6000 149.2000 160.9000 151.8000 ;
	    RECT 157.4000 148.8000 157.8000 149.2000 ;
	    RECT 160.6000 148.8000 161.0000 149.2000 ;
	    RECT 161.4000 148.2000 161.7000 151.8000 ;
	    RECT 159.8000 147.8000 160.2000 148.2000 ;
	    RECT 161.4000 147.8000 161.8000 148.2000 ;
	    RECT 155.0000 146.8000 155.4000 147.2000 ;
	    RECT 156.6000 146.8000 157.0000 147.2000 ;
	    RECT 152.6000 145.8000 153.0000 146.2000 ;
	    RECT 154.2000 145.8000 154.6000 146.2000 ;
	    RECT 151.0000 143.8000 151.4000 144.2000 ;
	    RECT 151.0000 139.2000 151.3000 143.8000 ;
	    RECT 152.6000 140.2000 152.9000 145.8000 ;
	    RECT 155.0000 144.2000 155.3000 146.8000 ;
	    RECT 157.4000 145.8000 157.8000 146.2000 ;
	    RECT 155.8000 144.8000 156.2000 145.2000 ;
	    RECT 155.8000 144.2000 156.1000 144.8000 ;
	    RECT 155.0000 143.8000 155.4000 144.2000 ;
	    RECT 155.8000 143.8000 156.2000 144.2000 ;
	    RECT 157.4000 143.2000 157.7000 145.8000 ;
	    RECT 158.2000 145.1000 158.6000 145.2000 ;
	    RECT 159.0000 145.1000 159.4000 145.2000 ;
	    RECT 158.2000 144.8000 159.4000 145.1000 ;
	    RECT 157.4000 142.8000 157.8000 143.2000 ;
	    RECT 157.4000 141.8000 157.8000 142.2000 ;
	    RECT 152.6000 139.8000 153.0000 140.2000 ;
	    RECT 155.0000 139.8000 155.4000 140.2000 ;
	    RECT 155.0000 139.2000 155.3000 139.8000 ;
	    RECT 151.0000 138.8000 151.4000 139.2000 ;
	    RECT 153.4000 138.8000 153.8000 139.2000 ;
	    RECT 155.0000 138.8000 155.4000 139.2000 ;
	    RECT 153.4000 138.2000 153.7000 138.8000 ;
	    RECT 157.4000 138.2000 157.7000 141.8000 ;
	    RECT 159.0000 140.8000 159.4000 141.2000 ;
	    RECT 159.0000 139.2000 159.3000 140.8000 ;
	    RECT 159.0000 138.8000 159.4000 139.2000 ;
	    RECT 153.4000 137.8000 153.8000 138.2000 ;
	    RECT 157.4000 137.8000 157.8000 138.2000 ;
	    RECT 159.8000 137.2000 160.1000 147.8000 ;
	    RECT 161.4000 145.8000 161.8000 146.2000 ;
	    RECT 161.4000 144.2000 161.7000 145.8000 ;
	    RECT 162.2000 145.1000 162.6000 147.9000 ;
	    RECT 161.4000 143.8000 161.8000 144.2000 ;
	    RECT 161.4000 142.2000 161.7000 143.8000 ;
	    RECT 163.8000 143.1000 164.2000 148.9000 ;
	    RECT 165.4000 147.2000 165.7000 153.8000 ;
	    RECT 167.8000 152.8000 168.2000 153.2000 ;
	    RECT 165.4000 147.1000 165.8000 147.2000 ;
	    RECT 166.2000 147.1000 166.6000 147.2000 ;
	    RECT 165.4000 146.8000 166.6000 147.1000 ;
	    RECT 165.4000 146.1000 165.8000 146.2000 ;
	    RECT 166.2000 146.1000 166.6000 146.2000 ;
	    RECT 165.4000 145.8000 166.6000 146.1000 ;
	    RECT 167.0000 143.8000 167.4000 144.2000 ;
	    RECT 161.4000 141.8000 161.8000 142.2000 ;
	    RECT 167.0000 139.2000 167.3000 143.8000 ;
	    RECT 167.8000 143.2000 168.1000 152.8000 ;
	    RECT 168.6000 152.1000 169.0000 157.9000 ;
	    RECT 167.8000 142.8000 168.2000 143.2000 ;
	    RECT 168.6000 143.1000 169.0000 148.9000 ;
	    RECT 169.4000 147.8000 169.8000 148.2000 ;
	    RECT 167.0000 138.8000 167.4000 139.2000 ;
	    RECT 150.2000 136.8000 150.6000 137.2000 ;
	    RECT 157.4000 137.1000 157.8000 137.2000 ;
	    RECT 158.2000 137.1000 158.6000 137.2000 ;
	    RECT 157.4000 136.8000 158.6000 137.1000 ;
	    RECT 159.8000 136.8000 160.2000 137.2000 ;
	    RECT 163.0000 136.8000 163.4000 137.2000 ;
	    RECT 163.0000 136.2000 163.3000 136.8000 ;
	    RECT 149.4000 135.8000 149.8000 136.2000 ;
	    RECT 151.0000 136.1000 151.4000 136.2000 ;
	    RECT 151.8000 136.1000 152.2000 136.2000 ;
	    RECT 151.0000 135.8000 152.2000 136.1000 ;
	    RECT 158.2000 135.8000 158.6000 136.2000 ;
	    RECT 159.0000 135.8000 159.4000 136.2000 ;
	    RECT 163.0000 135.8000 163.4000 136.2000 ;
	    RECT 167.8000 136.1000 168.2000 136.2000 ;
	    RECT 168.6000 136.1000 169.0000 136.2000 ;
	    RECT 167.8000 135.8000 169.0000 136.1000 ;
	    RECT 147.8000 134.8000 148.2000 135.2000 ;
	    RECT 147.0000 133.8000 148.1000 134.1000 ;
	    RECT 145.4000 133.1000 145.8000 133.2000 ;
	    RECT 146.2000 133.1000 146.6000 133.2000 ;
	    RECT 145.4000 132.8000 146.6000 133.1000 ;
	    RECT 147.0000 130.8000 147.4000 131.2000 ;
	    RECT 145.4000 129.8000 145.8000 130.2000 ;
	    RECT 142.2000 128.1000 142.6000 128.2000 ;
	    RECT 143.0000 128.1000 143.4000 128.2000 ;
	    RECT 142.2000 127.8000 143.4000 128.1000 ;
	    RECT 144.6000 127.8000 145.0000 128.2000 ;
	    RECT 138.2000 126.8000 138.6000 127.2000 ;
	    RECT 141.4000 126.8000 141.8000 127.2000 ;
	    RECT 143.8000 126.8000 144.2000 127.2000 ;
	    RECT 139.8000 124.8000 140.2000 125.2000 ;
	    RECT 139.8000 123.2000 140.1000 124.8000 ;
	    RECT 139.8000 122.8000 140.2000 123.2000 ;
	    RECT 135.0000 121.8000 135.4000 122.2000 ;
	    RECT 137.4000 121.8000 137.8000 122.2000 ;
	    RECT 139.0000 121.8000 139.4000 122.2000 ;
	    RECT 135.0000 116.2000 135.3000 121.8000 ;
	    RECT 139.0000 116.2000 139.3000 121.8000 ;
	    RECT 143.8000 119.2000 144.1000 126.8000 ;
	    RECT 144.6000 124.8000 145.0000 125.2000 ;
	    RECT 144.6000 123.2000 144.9000 124.8000 ;
	    RECT 144.6000 122.8000 145.0000 123.2000 ;
	    RECT 145.4000 119.2000 145.7000 129.8000 ;
	    RECT 147.0000 128.2000 147.3000 130.8000 ;
	    RECT 147.8000 129.2000 148.1000 133.8000 ;
	    RECT 149.4000 130.2000 149.7000 135.8000 ;
	    RECT 153.4000 134.8000 153.8000 135.2000 ;
	    RECT 151.0000 133.8000 151.4000 134.2000 ;
	    RECT 149.4000 129.8000 149.8000 130.2000 ;
	    RECT 147.8000 128.8000 148.2000 129.2000 ;
	    RECT 147.0000 127.8000 147.4000 128.2000 ;
	    RECT 148.6000 127.8000 149.0000 128.2000 ;
	    RECT 148.6000 127.2000 148.9000 127.8000 ;
	    RECT 146.2000 126.8000 146.6000 127.2000 ;
	    RECT 148.6000 126.8000 149.0000 127.2000 ;
	    RECT 150.2000 127.1000 150.6000 127.2000 ;
	    RECT 151.0000 127.1000 151.3000 133.8000 ;
	    RECT 153.4000 128.1000 153.7000 134.8000 ;
	    RECT 155.8000 134.3000 156.2000 134.4000 ;
	    RECT 156.6000 134.3000 157.0000 134.4000 ;
	    RECT 154.2000 133.8000 154.6000 134.2000 ;
	    RECT 155.8000 134.0000 157.0000 134.3000 ;
	    RECT 158.2000 134.2000 158.5000 135.8000 ;
	    RECT 159.0000 135.2000 159.3000 135.8000 ;
	    RECT 159.0000 134.8000 159.4000 135.2000 ;
	    RECT 164.6000 134.8000 165.0000 135.2000 ;
	    RECT 165.4000 134.8000 165.8000 135.2000 ;
	    RECT 166.2000 135.1000 166.6000 135.2000 ;
	    RECT 167.0000 135.1000 167.4000 135.2000 ;
	    RECT 166.2000 134.8000 167.4000 135.1000 ;
	    RECT 164.6000 134.2000 164.9000 134.8000 ;
	    RECT 165.4000 134.2000 165.7000 134.8000 ;
	    RECT 169.4000 134.2000 169.7000 147.8000 ;
	    RECT 171.0000 141.8000 171.4000 142.2000 ;
	    RECT 157.4000 133.8000 157.8000 134.2000 ;
	    RECT 158.2000 133.8000 158.6000 134.2000 ;
	    RECT 159.8000 133.8000 160.2000 134.2000 ;
	    RECT 162.2000 134.1000 162.6000 134.2000 ;
	    RECT 163.0000 134.1000 163.4000 134.2000 ;
	    RECT 162.2000 133.8000 163.4000 134.1000 ;
	    RECT 164.6000 133.8000 165.0000 134.2000 ;
	    RECT 165.4000 133.8000 165.8000 134.2000 ;
	    RECT 166.2000 134.1000 166.6000 134.2000 ;
	    RECT 167.0000 134.1000 167.4000 134.2000 ;
	    RECT 166.2000 133.8000 167.4000 134.1000 ;
	    RECT 169.4000 133.8000 169.8000 134.2000 ;
	    RECT 154.2000 130.2000 154.5000 133.8000 ;
	    RECT 156.6000 131.8000 157.0000 132.2000 ;
	    RECT 154.2000 129.8000 154.6000 130.2000 ;
	    RECT 154.2000 129.1000 154.6000 129.2000 ;
	    RECT 155.0000 129.1000 155.4000 129.2000 ;
	    RECT 154.2000 128.8000 155.4000 129.1000 ;
	    RECT 153.4000 127.8000 154.5000 128.1000 ;
	    RECT 150.2000 126.8000 151.3000 127.1000 ;
	    RECT 143.8000 118.8000 144.2000 119.2000 ;
	    RECT 145.4000 118.8000 145.8000 119.2000 ;
	    RECT 135.0000 115.8000 135.4000 116.2000 ;
	    RECT 135.8000 116.1000 136.2000 116.2000 ;
	    RECT 135.8000 115.8000 136.9000 116.1000 ;
	    RECT 139.0000 115.8000 139.4000 116.2000 ;
	    RECT 140.6000 115.8000 141.0000 116.2000 ;
	    RECT 135.0000 115.1000 135.4000 115.2000 ;
	    RECT 135.8000 115.1000 136.2000 115.2000 ;
	    RECT 135.0000 114.8000 136.2000 115.1000 ;
	    RECT 135.8000 111.8000 136.2000 112.2000 ;
	    RECT 134.2000 108.8000 134.6000 109.2000 ;
	    RECT 135.8000 107.2000 136.1000 111.8000 ;
	    RECT 136.6000 107.2000 136.9000 115.8000 ;
	    RECT 140.6000 115.2000 140.9000 115.8000 ;
	    RECT 137.4000 114.8000 137.8000 115.2000 ;
	    RECT 140.6000 115.1000 141.0000 115.2000 ;
	    RECT 144.6000 115.1000 145.0000 115.2000 ;
	    RECT 140.6000 114.8000 141.7000 115.1000 ;
	    RECT 133.4000 106.8000 133.8000 107.2000 ;
	    RECT 135.8000 106.8000 136.2000 107.2000 ;
	    RECT 136.6000 106.8000 137.0000 107.2000 ;
	    RECT 127.0000 106.1000 127.4000 106.2000 ;
	    RECT 127.8000 106.1000 128.2000 106.2000 ;
	    RECT 127.0000 105.8000 128.2000 106.1000 ;
	    RECT 129.4000 106.1000 129.8000 106.2000 ;
	    RECT 130.2000 106.1000 130.6000 106.2000 ;
	    RECT 129.4000 105.8000 130.6000 106.1000 ;
	    RECT 132.6000 105.8000 133.0000 106.2000 ;
	    RECT 130.2000 104.8000 130.6000 105.2000 ;
	    RECT 126.2000 101.8000 126.6000 102.2000 ;
	    RECT 128.6000 101.8000 129.0000 102.2000 ;
	    RECT 124.6000 100.8000 125.0000 101.2000 ;
	    RECT 126.2000 99.8000 126.6000 100.2000 ;
	    RECT 127.0000 99.8000 127.4000 100.2000 ;
	    RECT 126.2000 99.2000 126.5000 99.8000 ;
	    RECT 127.0000 99.2000 127.3000 99.8000 ;
	    RECT 126.2000 98.8000 126.6000 99.2000 ;
	    RECT 127.0000 98.8000 127.4000 99.2000 ;
	    RECT 123.8000 92.1000 124.2000 97.9000 ;
	    RECT 128.6000 90.2000 128.9000 101.8000 ;
	    RECT 129.4000 92.1000 129.8000 97.9000 ;
	    RECT 130.2000 95.2000 130.5000 104.8000 ;
	    RECT 131.8000 103.8000 132.2000 104.2000 ;
	    RECT 130.2000 94.8000 130.6000 95.2000 ;
	    RECT 125.4000 89.8000 125.8000 90.2000 ;
	    RECT 128.6000 89.8000 129.0000 90.2000 ;
	    RECT 123.0000 86.8000 123.4000 87.2000 ;
	    RECT 115.8000 72.1000 116.2000 77.9000 ;
	    RECT 116.6000 74.7000 117.0000 75.1000 ;
	    RECT 116.6000 74.2000 116.9000 74.7000 ;
	    RECT 116.6000 73.8000 117.0000 74.2000 ;
	    RECT 118.2000 73.8000 118.6000 74.2000 ;
	    RECT 116.6000 71.8000 117.0000 72.2000 ;
	    RECT 110.2000 66.8000 110.6000 67.2000 ;
	    RECT 115.0000 66.8000 115.4000 67.2000 ;
	    RECT 110.2000 59.2000 110.5000 66.8000 ;
	    RECT 116.6000 59.2000 116.9000 71.8000 ;
	    RECT 118.2000 69.2000 118.5000 73.8000 ;
	    RECT 120.6000 72.1000 121.0000 77.9000 ;
	    RECT 123.0000 74.1000 123.3000 86.8000 ;
	    RECT 125.4000 86.2000 125.7000 89.8000 ;
	    RECT 131.8000 89.2000 132.1000 103.8000 ;
	    RECT 133.4000 103.2000 133.7000 106.8000 ;
	    RECT 137.4000 105.2000 137.7000 114.8000 ;
	    RECT 141.4000 114.2000 141.7000 114.8000 ;
	    RECT 143.8000 114.8000 145.0000 115.1000 ;
	    RECT 146.2000 115.1000 146.5000 126.8000 ;
	    RECT 149.4000 125.8000 149.8000 126.2000 ;
	    RECT 149.4000 117.2000 149.7000 125.8000 ;
	    RECT 147.0000 116.8000 147.4000 117.2000 ;
	    RECT 149.4000 116.8000 149.8000 117.2000 ;
	    RECT 147.0000 116.2000 147.3000 116.8000 ;
	    RECT 147.0000 115.8000 147.4000 116.2000 ;
	    RECT 147.8000 115.8000 148.2000 116.2000 ;
	    RECT 147.8000 115.2000 148.1000 115.8000 ;
	    RECT 149.4000 115.2000 149.7000 116.8000 ;
	    RECT 151.0000 116.2000 151.3000 126.8000 ;
	    RECT 153.4000 126.8000 153.8000 127.2000 ;
	    RECT 153.4000 126.2000 153.7000 126.8000 ;
	    RECT 153.4000 125.8000 153.8000 126.2000 ;
	    RECT 151.8000 124.8000 152.2000 125.2000 ;
	    RECT 151.8000 117.2000 152.1000 124.8000 ;
	    RECT 151.8000 116.8000 152.2000 117.2000 ;
	    RECT 152.6000 116.8000 153.0000 117.2000 ;
	    RECT 152.6000 116.2000 152.9000 116.8000 ;
	    RECT 151.0000 116.1000 151.4000 116.2000 ;
	    RECT 151.8000 116.1000 152.2000 116.2000 ;
	    RECT 151.0000 115.8000 152.2000 116.1000 ;
	    RECT 152.6000 115.8000 153.0000 116.2000 ;
	    RECT 154.2000 115.2000 154.5000 127.8000 ;
	    RECT 155.0000 127.8000 155.4000 128.2000 ;
	    RECT 155.0000 127.2000 155.3000 127.8000 ;
	    RECT 155.0000 126.8000 155.4000 127.2000 ;
	    RECT 155.8000 125.8000 156.2000 126.2000 ;
	    RECT 155.8000 119.2000 156.1000 125.8000 ;
	    RECT 156.6000 125.2000 156.9000 131.8000 ;
	    RECT 157.4000 130.2000 157.7000 133.8000 ;
	    RECT 157.4000 129.8000 157.8000 130.2000 ;
	    RECT 159.0000 129.8000 159.4000 130.2000 ;
	    RECT 158.2000 128.8000 158.6000 129.2000 ;
	    RECT 158.2000 127.2000 158.5000 128.8000 ;
	    RECT 158.2000 126.8000 158.6000 127.2000 ;
	    RECT 159.0000 125.2000 159.3000 129.8000 ;
	    RECT 159.8000 129.2000 160.1000 133.8000 ;
	    RECT 161.4000 132.8000 161.8000 133.2000 ;
	    RECT 163.0000 132.8000 163.4000 133.2000 ;
	    RECT 161.4000 132.2000 161.7000 132.8000 ;
	    RECT 161.4000 131.8000 161.8000 132.2000 ;
	    RECT 163.0000 131.2000 163.3000 132.8000 ;
	    RECT 166.2000 131.8000 166.6000 132.2000 ;
	    RECT 163.0000 130.8000 163.4000 131.2000 ;
	    RECT 159.8000 128.8000 160.2000 129.2000 ;
	    RECT 161.4000 127.8000 161.8000 128.2000 ;
	    RECT 161.4000 127.2000 161.7000 127.8000 ;
	    RECT 160.6000 126.8000 161.0000 127.2000 ;
	    RECT 161.4000 126.8000 161.8000 127.2000 ;
	    RECT 163.0000 127.1000 163.4000 127.2000 ;
	    RECT 162.2000 126.8000 163.4000 127.1000 ;
	    RECT 160.6000 126.2000 160.9000 126.8000 ;
	    RECT 162.2000 126.2000 162.5000 126.8000 ;
	    RECT 160.6000 125.8000 161.0000 126.2000 ;
	    RECT 162.2000 125.8000 162.6000 126.2000 ;
	    RECT 156.6000 124.8000 157.0000 125.2000 ;
	    RECT 159.0000 124.8000 159.4000 125.2000 ;
	    RECT 160.6000 125.1000 161.0000 125.2000 ;
	    RECT 161.4000 125.1000 161.8000 125.2000 ;
	    RECT 160.6000 124.8000 161.8000 125.1000 ;
	    RECT 156.6000 124.2000 156.9000 124.8000 ;
	    RECT 156.6000 123.8000 157.0000 124.2000 ;
	    RECT 161.4000 123.8000 161.8000 124.2000 ;
	    RECT 155.8000 118.8000 156.2000 119.2000 ;
	    RECT 158.2000 116.8000 158.6000 117.2000 ;
	    RECT 158.2000 116.2000 158.5000 116.8000 ;
	    RECT 156.6000 115.8000 157.0000 116.2000 ;
	    RECT 158.2000 115.8000 158.6000 116.2000 ;
	    RECT 160.6000 115.8000 161.0000 116.2000 ;
	    RECT 147.0000 115.1000 147.4000 115.2000 ;
	    RECT 146.2000 114.8000 147.4000 115.1000 ;
	    RECT 147.8000 114.8000 148.2000 115.2000 ;
	    RECT 149.4000 114.8000 149.8000 115.2000 ;
	    RECT 154.2000 114.8000 154.6000 115.2000 ;
	    RECT 138.2000 113.8000 138.6000 114.2000 ;
	    RECT 139.8000 114.1000 140.2000 114.2000 ;
	    RECT 140.6000 114.1000 141.0000 114.2000 ;
	    RECT 139.8000 113.8000 141.0000 114.1000 ;
	    RECT 141.4000 113.8000 141.8000 114.2000 ;
	    RECT 142.2000 114.0000 142.6000 114.4000 ;
	    RECT 138.2000 112.2000 138.5000 113.8000 ;
	    RECT 142.2000 113.2000 142.5000 114.0000 ;
	    RECT 140.6000 112.8000 141.0000 113.2000 ;
	    RECT 142.2000 112.8000 142.6000 113.2000 ;
	    RECT 138.2000 111.8000 138.6000 112.2000 ;
	    RECT 140.6000 109.2000 140.9000 112.8000 ;
	    RECT 142.2000 111.8000 142.6000 112.2000 ;
	    RECT 140.6000 108.8000 141.0000 109.2000 ;
	    RECT 141.4000 108.8000 141.8000 109.2000 ;
	    RECT 141.4000 108.2000 141.7000 108.8000 ;
	    RECT 142.2000 108.2000 142.5000 111.8000 ;
	    RECT 138.2000 107.8000 138.6000 108.2000 ;
	    RECT 141.4000 107.8000 141.8000 108.2000 ;
	    RECT 142.2000 107.8000 142.6000 108.2000 ;
	    RECT 138.2000 107.2000 138.5000 107.8000 ;
	    RECT 138.2000 106.8000 138.6000 107.2000 ;
	    RECT 139.0000 107.1000 139.4000 107.2000 ;
	    RECT 139.8000 107.1000 140.2000 107.2000 ;
	    RECT 139.0000 106.8000 140.2000 107.1000 ;
	    RECT 136.6000 105.1000 137.0000 105.2000 ;
	    RECT 137.4000 105.1000 137.8000 105.2000 ;
	    RECT 136.6000 104.8000 137.8000 105.1000 ;
	    RECT 139.0000 104.8000 139.4000 105.2000 ;
	    RECT 143.0000 105.1000 143.4000 107.9000 ;
	    RECT 133.4000 102.8000 133.8000 103.2000 ;
	    RECT 137.4000 102.8000 137.8000 103.2000 ;
	    RECT 136.6000 100.8000 137.0000 101.2000 ;
	    RECT 132.6000 94.8000 133.0000 95.2000 ;
	    RECT 132.6000 94.2000 132.9000 94.8000 ;
	    RECT 132.6000 93.8000 133.0000 94.2000 ;
	    RECT 134.2000 92.1000 134.6000 97.9000 ;
	    RECT 136.6000 96.2000 136.9000 100.8000 ;
	    RECT 137.4000 99.2000 137.7000 102.8000 ;
	    RECT 138.2000 101.8000 138.6000 102.2000 ;
	    RECT 138.2000 99.2000 138.5000 101.8000 ;
	    RECT 139.0000 99.2000 139.3000 104.8000 ;
	    RECT 137.4000 98.8000 137.8000 99.2000 ;
	    RECT 138.2000 98.8000 138.6000 99.2000 ;
	    RECT 139.0000 98.8000 139.4000 99.2000 ;
	    RECT 142.2000 99.1000 142.6000 99.2000 ;
	    RECT 143.0000 99.1000 143.4000 99.2000 ;
	    RECT 142.2000 98.8000 143.4000 99.1000 ;
	    RECT 135.0000 94.8000 135.4000 95.2000 ;
	    RECT 135.0000 94.2000 135.3000 94.8000 ;
	    RECT 135.0000 93.8000 135.4000 94.2000 ;
	    RECT 135.8000 93.1000 136.2000 95.9000 ;
	    RECT 136.6000 95.8000 137.0000 96.2000 ;
	    RECT 136.6000 89.2000 136.9000 95.8000 ;
	    RECT 138.2000 94.2000 138.5000 98.8000 ;
	    RECT 143.8000 98.1000 144.1000 114.8000 ;
	    RECT 144.6000 113.8000 145.0000 114.2000 ;
	    RECT 144.6000 113.2000 144.9000 113.8000 ;
	    RECT 144.6000 112.8000 145.0000 113.2000 ;
	    RECT 144.6000 103.1000 145.0000 108.9000 ;
	    RECT 146.2000 106.8000 146.6000 107.2000 ;
	    RECT 145.4000 105.9000 145.8000 106.3000 ;
	    RECT 145.4000 104.2000 145.7000 105.9000 ;
	    RECT 145.4000 103.8000 145.8000 104.2000 ;
	    RECT 143.0000 97.8000 144.1000 98.1000 ;
	    RECT 138.2000 93.8000 138.6000 94.2000 ;
	    RECT 139.8000 92.8000 140.2000 93.2000 ;
	    RECT 142.2000 92.8000 142.6000 93.2000 ;
	    RECT 125.4000 85.8000 125.8000 86.2000 ;
	    RECT 126.2000 84.8000 126.6000 85.2000 ;
	    RECT 126.2000 79.2000 126.5000 84.8000 ;
	    RECT 127.0000 83.1000 127.4000 88.9000 ;
	    RECT 131.8000 88.8000 132.2000 89.2000 ;
	    RECT 127.8000 86.8000 128.2000 87.2000 ;
	    RECT 127.8000 83.2000 128.1000 86.8000 ;
	    RECT 128.6000 85.1000 129.0000 87.9000 ;
	    RECT 129.4000 87.8000 129.8000 88.2000 ;
	    RECT 129.4000 87.2000 129.7000 87.8000 ;
	    RECT 129.4000 86.8000 129.8000 87.2000 ;
	    RECT 129.4000 86.1000 129.8000 86.2000 ;
	    RECT 130.2000 86.1000 130.6000 86.2000 ;
	    RECT 129.4000 85.8000 130.6000 86.1000 ;
	    RECT 132.6000 85.1000 133.0000 87.9000 ;
	    RECT 133.4000 86.8000 133.8000 87.2000 ;
	    RECT 133.4000 83.2000 133.7000 86.8000 ;
	    RECT 127.8000 82.8000 128.2000 83.2000 ;
	    RECT 133.4000 82.8000 133.8000 83.2000 ;
	    RECT 134.2000 83.1000 134.6000 88.9000 ;
	    RECT 136.6000 88.8000 137.0000 89.2000 ;
	    RECT 135.0000 85.9000 135.4000 86.3000 ;
	    RECT 135.0000 85.2000 135.3000 85.9000 ;
	    RECT 135.0000 84.8000 135.4000 85.2000 ;
	    RECT 139.0000 83.1000 139.4000 88.9000 ;
	    RECT 126.2000 78.8000 126.6000 79.2000 ;
	    RECT 123.8000 75.8000 124.2000 76.2000 ;
	    RECT 123.8000 75.1000 124.1000 75.8000 ;
	    RECT 124.6000 75.1000 125.0000 75.2000 ;
	    RECT 123.8000 74.8000 125.0000 75.1000 ;
	    RECT 123.8000 74.1000 124.2000 74.2000 ;
	    RECT 123.0000 73.8000 124.2000 74.1000 ;
	    RECT 127.0000 73.1000 127.4000 75.9000 ;
	    RECT 127.8000 74.2000 128.1000 82.8000 ;
	    RECT 139.8000 79.2000 140.1000 92.8000 ;
	    RECT 142.2000 92.2000 142.5000 92.8000 ;
	    RECT 142.2000 91.8000 142.6000 92.2000 ;
	    RECT 142.2000 89.8000 142.6000 90.2000 ;
	    RECT 140.6000 89.1000 141.0000 89.2000 ;
	    RECT 141.4000 89.1000 141.8000 89.2000 ;
	    RECT 140.6000 88.8000 141.8000 89.1000 ;
	    RECT 142.2000 88.2000 142.5000 89.8000 ;
	    RECT 143.0000 89.2000 143.3000 97.8000 ;
	    RECT 144.6000 95.8000 145.0000 96.2000 ;
	    RECT 143.0000 88.8000 143.4000 89.2000 ;
	    RECT 142.2000 87.8000 142.6000 88.2000 ;
	    RECT 143.8000 87.8000 144.2000 88.2000 ;
	    RECT 143.8000 87.2000 144.1000 87.8000 ;
	    RECT 143.8000 86.8000 144.2000 87.2000 ;
	    RECT 144.6000 86.2000 144.9000 95.8000 ;
	    RECT 145.4000 92.1000 145.8000 97.9000 ;
	    RECT 146.2000 95.2000 146.5000 106.8000 ;
	    RECT 146.2000 94.8000 146.6000 95.2000 ;
	    RECT 147.8000 87.2000 148.1000 114.8000 ;
	    RECT 154.2000 114.2000 154.5000 114.8000 ;
	    RECT 156.6000 114.2000 156.9000 115.8000 ;
	    RECT 160.6000 115.2000 160.9000 115.8000 ;
	    RECT 161.4000 115.2000 161.7000 123.8000 ;
	    RECT 159.8000 114.8000 160.2000 115.2000 ;
	    RECT 160.6000 114.8000 161.0000 115.2000 ;
	    RECT 161.4000 114.8000 161.8000 115.2000 ;
	    RECT 159.8000 114.2000 160.1000 114.8000 ;
	    RECT 162.2000 114.2000 162.5000 125.8000 ;
	    RECT 163.8000 125.1000 164.2000 127.9000 ;
	    RECT 165.4000 123.1000 165.8000 128.9000 ;
	    RECT 166.2000 127.2000 166.5000 131.8000 ;
	    RECT 166.2000 126.8000 166.6000 127.2000 ;
	    RECT 167.0000 126.8000 167.4000 127.2000 ;
	    RECT 150.2000 113.8000 150.6000 114.2000 ;
	    RECT 151.8000 114.1000 152.2000 114.2000 ;
	    RECT 152.6000 114.1000 153.0000 114.2000 ;
	    RECT 151.8000 113.8000 153.0000 114.1000 ;
	    RECT 154.2000 113.8000 154.6000 114.2000 ;
	    RECT 155.0000 113.8000 155.4000 114.2000 ;
	    RECT 156.6000 113.8000 157.0000 114.2000 ;
	    RECT 157.4000 113.8000 157.8000 114.2000 ;
	    RECT 159.8000 113.8000 160.2000 114.2000 ;
	    RECT 161.4000 114.1000 161.8000 114.2000 ;
	    RECT 162.2000 114.1000 162.6000 114.2000 ;
	    RECT 161.4000 113.8000 162.6000 114.1000 ;
	    RECT 150.2000 113.2000 150.5000 113.8000 ;
	    RECT 150.2000 112.8000 150.6000 113.2000 ;
	    RECT 151.0000 111.8000 151.4000 112.2000 ;
	    RECT 149.4000 103.1000 149.8000 108.9000 ;
	    RECT 148.6000 94.8000 149.0000 95.2000 ;
	    RECT 147.8000 86.8000 148.2000 87.2000 ;
	    RECT 144.6000 85.8000 145.0000 86.2000 ;
	    RECT 148.6000 85.2000 148.9000 94.8000 ;
	    RECT 150.2000 92.1000 150.6000 97.9000 ;
	    RECT 151.0000 96.2000 151.3000 111.8000 ;
	    RECT 151.8000 109.2000 152.1000 113.8000 ;
	    RECT 155.0000 113.2000 155.3000 113.8000 ;
	    RECT 157.4000 113.2000 157.7000 113.8000 ;
	    RECT 152.6000 112.8000 153.0000 113.2000 ;
	    RECT 155.0000 112.8000 155.4000 113.2000 ;
	    RECT 157.4000 112.8000 157.8000 113.2000 ;
	    RECT 163.0000 113.1000 163.4000 115.9000 ;
	    RECT 152.6000 109.2000 152.9000 112.8000 ;
	    RECT 164.6000 112.1000 165.0000 117.9000 ;
	    RECT 166.2000 114.2000 166.5000 126.8000 ;
	    RECT 167.0000 126.2000 167.3000 126.8000 ;
	    RECT 167.0000 125.8000 167.4000 126.2000 ;
	    RECT 170.2000 123.1000 170.6000 128.9000 ;
	    RECT 167.0000 115.1000 167.4000 115.2000 ;
	    RECT 167.8000 115.1000 168.2000 115.2000 ;
	    RECT 167.0000 114.8000 168.2000 115.1000 ;
	    RECT 166.2000 113.8000 166.6000 114.2000 ;
	    RECT 165.4000 112.8000 165.8000 113.2000 ;
	    RECT 151.8000 108.8000 152.2000 109.2000 ;
	    RECT 152.6000 108.8000 153.0000 109.2000 ;
	    RECT 155.0000 103.1000 155.4000 108.9000 ;
	    RECT 155.8000 105.8000 156.2000 106.2000 ;
	    RECT 159.0000 105.9000 159.4000 106.3000 ;
	    RECT 151.0000 95.8000 151.4000 96.2000 ;
	    RECT 151.0000 94.8000 151.4000 95.2000 ;
	    RECT 151.0000 94.2000 151.3000 94.8000 ;
	    RECT 151.0000 93.8000 151.4000 94.2000 ;
	    RECT 151.8000 93.1000 152.2000 95.9000 ;
	    RECT 155.8000 95.2000 156.1000 105.8000 ;
	    RECT 159.0000 104.2000 159.3000 105.9000 ;
	    RECT 159.0000 103.8000 159.4000 104.2000 ;
	    RECT 159.8000 103.1000 160.2000 108.9000 ;
	    RECT 161.4000 105.1000 161.8000 107.9000 ;
	    RECT 162.2000 105.1000 162.6000 107.9000 ;
	    RECT 163.0000 106.8000 163.4000 107.2000 ;
	    RECT 152.6000 94.8000 153.0000 95.2000 ;
	    RECT 155.8000 94.8000 156.2000 95.2000 ;
	    RECT 152.6000 94.2000 152.9000 94.8000 ;
	    RECT 152.6000 93.8000 153.0000 94.2000 ;
	    RECT 159.8000 93.1000 160.2000 95.9000 ;
	    RECT 160.6000 93.8000 161.0000 94.2000 ;
	    RECT 151.0000 91.8000 151.4000 92.2000 ;
	    RECT 151.0000 89.2000 151.3000 91.8000 ;
	    RECT 152.6000 89.8000 153.0000 90.2000 ;
	    RECT 152.6000 89.2000 152.9000 89.8000 ;
	    RECT 151.0000 88.8000 151.4000 89.2000 ;
	    RECT 152.6000 88.8000 153.0000 89.2000 ;
	    RECT 144.6000 84.8000 145.0000 85.2000 ;
	    RECT 148.6000 84.8000 149.0000 85.2000 ;
	    RECT 143.8000 79.8000 144.2000 80.2000 ;
	    RECT 135.8000 79.1000 136.2000 79.2000 ;
	    RECT 136.6000 79.1000 137.0000 79.2000 ;
	    RECT 135.8000 78.8000 137.0000 79.1000 ;
	    RECT 139.8000 78.8000 140.2000 79.2000 ;
	    RECT 127.8000 73.8000 128.2000 74.2000 ;
	    RECT 118.2000 68.8000 118.6000 69.2000 ;
	    RECT 118.2000 67.2000 118.5000 68.8000 ;
	    RECT 118.2000 66.8000 118.6000 67.2000 ;
	    RECT 119.8000 65.1000 120.2000 67.9000 ;
	    RECT 120.6000 67.8000 121.0000 68.2000 ;
	    RECT 120.6000 67.2000 120.9000 67.8000 ;
	    RECT 120.6000 66.8000 121.0000 67.2000 ;
	    RECT 121.4000 63.1000 121.8000 68.9000 ;
	    RECT 122.2000 65.9000 122.6000 66.3000 ;
	    RECT 122.2000 65.2000 122.5000 65.9000 ;
	    RECT 122.2000 64.8000 122.6000 65.2000 ;
	    RECT 126.2000 63.1000 126.6000 68.9000 ;
	    RECT 127.8000 68.2000 128.1000 73.8000 ;
	    RECT 128.6000 72.1000 129.0000 77.9000 ;
	    RECT 129.4000 74.7000 129.8000 75.1000 ;
	    RECT 129.4000 69.2000 129.7000 74.7000 ;
	    RECT 133.4000 72.1000 133.8000 77.9000 ;
	    RECT 136.6000 75.8000 137.0000 76.2000 ;
	    RECT 136.6000 75.2000 136.9000 75.8000 ;
	    RECT 143.8000 75.2000 144.1000 79.8000 ;
	    RECT 136.6000 74.8000 137.0000 75.2000 ;
	    RECT 143.8000 74.8000 144.2000 75.2000 ;
	    RECT 137.4000 73.8000 137.8000 74.2000 ;
	    RECT 142.2000 73.8000 142.6000 74.2000 ;
	    RECT 143.0000 73.8000 143.4000 74.2000 ;
	    RECT 143.8000 73.8000 144.2000 74.2000 ;
	    RECT 129.4000 68.8000 129.8000 69.2000 ;
	    RECT 127.8000 67.8000 128.2000 68.2000 ;
	    RECT 128.6000 66.8000 129.0000 67.2000 ;
	    RECT 131.8000 66.8000 132.2000 67.2000 ;
	    RECT 128.6000 66.2000 128.9000 66.8000 ;
	    RECT 131.8000 66.2000 132.1000 66.8000 ;
	    RECT 128.6000 65.8000 129.0000 66.2000 ;
	    RECT 130.2000 66.1000 130.6000 66.2000 ;
	    RECT 131.0000 66.1000 131.4000 66.2000 ;
	    RECT 130.2000 65.8000 131.4000 66.1000 ;
	    RECT 131.8000 65.8000 132.2000 66.2000 ;
	    RECT 132.6000 65.1000 133.0000 67.9000 ;
	    RECT 133.4000 67.8000 133.8000 68.2000 ;
	    RECT 133.4000 67.2000 133.7000 67.8000 ;
	    RECT 133.4000 66.8000 133.8000 67.2000 ;
	    RECT 134.2000 63.1000 134.6000 68.9000 ;
	    RECT 135.8000 66.1000 136.2000 66.2000 ;
	    RECT 136.6000 66.1000 137.0000 66.2000 ;
	    RECT 135.8000 65.8000 137.0000 66.1000 ;
	    RECT 137.4000 59.2000 137.7000 73.8000 ;
	    RECT 139.0000 73.1000 139.4000 73.2000 ;
	    RECT 139.8000 73.1000 140.2000 73.2000 ;
	    RECT 139.0000 72.8000 140.2000 73.1000 ;
	    RECT 138.2000 71.8000 138.6000 72.2000 ;
	    RECT 138.2000 66.2000 138.5000 71.8000 ;
	    RECT 142.2000 69.2000 142.5000 73.8000 ;
	    RECT 143.0000 73.2000 143.3000 73.8000 ;
	    RECT 143.0000 72.8000 143.4000 73.2000 ;
	    RECT 138.2000 65.8000 138.6000 66.2000 ;
	    RECT 139.0000 63.1000 139.4000 68.9000 ;
	    RECT 142.2000 68.8000 142.6000 69.2000 ;
	    RECT 142.2000 67.2000 142.5000 68.8000 ;
	    RECT 142.2000 66.8000 142.6000 67.2000 ;
	    RECT 143.0000 66.1000 143.4000 66.2000 ;
	    RECT 142.2000 65.8000 143.4000 66.1000 ;
	    RECT 142.2000 65.2000 142.5000 65.8000 ;
	    RECT 142.2000 64.8000 142.6000 65.2000 ;
	    RECT 110.2000 58.8000 110.6000 59.2000 ;
	    RECT 116.6000 58.8000 117.0000 59.2000 ;
	    RECT 133.4000 59.1000 133.8000 59.2000 ;
	    RECT 134.2000 59.1000 134.6000 59.2000 ;
	    RECT 133.4000 58.8000 134.6000 59.1000 ;
	    RECT 137.4000 58.8000 137.8000 59.2000 ;
	    RECT 135.8000 57.8000 136.2000 58.2000 ;
	    RECT 142.2000 57.8000 142.6000 58.2000 ;
	    RECT 143.0000 57.8000 143.4000 58.2000 ;
	    RECT 108.6000 57.1000 109.0000 57.2000 ;
	    RECT 109.4000 57.1000 109.8000 57.2000 ;
	    RECT 108.6000 56.8000 109.8000 57.1000 ;
	    RECT 117.4000 57.1000 117.8000 57.2000 ;
	    RECT 118.2000 57.1000 118.6000 57.2000 ;
	    RECT 117.4000 56.8000 118.6000 57.1000 ;
	    RECT 135.8000 55.2000 136.1000 57.8000 ;
	    RECT 142.2000 57.2000 142.5000 57.8000 ;
	    RECT 143.0000 57.2000 143.3000 57.8000 ;
	    RECT 136.6000 56.8000 137.0000 57.2000 ;
	    RECT 142.2000 56.8000 142.6000 57.2000 ;
	    RECT 143.0000 56.8000 143.4000 57.2000 ;
	    RECT 136.6000 56.2000 136.9000 56.8000 ;
	    RECT 136.6000 55.8000 137.0000 56.2000 ;
	    RECT 140.6000 55.8000 141.0000 56.2000 ;
	    RECT 142.2000 56.1000 142.6000 56.2000 ;
	    RECT 143.0000 56.1000 143.4000 56.2000 ;
	    RECT 142.2000 55.8000 143.4000 56.1000 ;
	    RECT 140.6000 55.2000 140.9000 55.8000 ;
	    RECT 109.4000 54.8000 109.8000 55.2000 ;
	    RECT 116.6000 54.8000 117.0000 55.2000 ;
	    RECT 135.8000 54.8000 136.2000 55.2000 ;
	    RECT 140.6000 54.8000 141.0000 55.2000 ;
	    RECT 142.2000 54.8000 142.6000 55.2000 ;
	    RECT 108.6000 53.8000 109.0000 54.2000 ;
	    RECT 108.6000 46.2000 108.9000 53.8000 ;
	    RECT 108.6000 45.8000 109.0000 46.2000 ;
	    RECT 108.6000 44.8000 109.0000 45.2000 ;
	    RECT 108.6000 44.2000 108.9000 44.8000 ;
	    RECT 108.6000 43.8000 109.0000 44.2000 ;
	    RECT 109.4000 39.2000 109.7000 54.8000 ;
	    RECT 111.8000 54.1000 112.2000 54.2000 ;
	    RECT 112.6000 54.1000 113.0000 54.2000 ;
	    RECT 111.8000 53.8000 113.0000 54.1000 ;
	    RECT 116.6000 51.2000 116.9000 54.8000 ;
	    RECT 121.4000 53.8000 121.8000 54.2000 ;
	    RECT 122.2000 54.1000 122.6000 54.2000 ;
	    RECT 123.0000 54.1000 123.4000 54.2000 ;
	    RECT 122.2000 53.8000 123.4000 54.1000 ;
	    RECT 124.6000 54.1000 125.0000 54.2000 ;
	    RECT 125.4000 54.1000 125.8000 54.2000 ;
	    RECT 124.6000 53.8000 125.8000 54.1000 ;
	    RECT 128.6000 54.1000 129.0000 54.2000 ;
	    RECT 129.4000 54.1000 129.8000 54.2000 ;
	    RECT 128.6000 53.8000 129.8000 54.1000 ;
	    RECT 135.0000 53.8000 135.4000 54.2000 ;
	    RECT 120.6000 51.8000 121.0000 52.2000 ;
	    RECT 116.6000 50.8000 117.0000 51.2000 ;
	    RECT 120.6000 50.2000 120.9000 51.8000 ;
	    RECT 118.2000 49.8000 118.6000 50.2000 ;
	    RECT 120.6000 49.8000 121.0000 50.2000 ;
	    RECT 112.6000 45.8000 113.0000 46.2000 ;
	    RECT 116.6000 46.1000 117.0000 46.2000 ;
	    RECT 117.4000 46.1000 117.8000 46.2000 ;
	    RECT 116.6000 45.8000 117.8000 46.1000 ;
	    RECT 110.2000 39.8000 110.6000 40.2000 ;
	    RECT 107.0000 38.8000 107.4000 39.2000 ;
	    RECT 109.4000 38.8000 109.8000 39.2000 ;
	    RECT 109.4000 37.8000 109.8000 38.2000 ;
	    RECT 106.2000 36.8000 106.6000 37.2000 ;
	    RECT 109.4000 36.2000 109.7000 37.8000 ;
	    RECT 110.2000 37.2000 110.5000 39.8000 ;
	    RECT 110.2000 36.8000 110.6000 37.2000 ;
	    RECT 102.2000 35.8000 102.6000 36.2000 ;
	    RECT 104.6000 35.8000 105.0000 36.2000 ;
	    RECT 109.4000 35.8000 109.8000 36.2000 ;
	    RECT 102.2000 34.2000 102.5000 35.8000 ;
	    RECT 103.8000 35.1000 104.2000 35.2000 ;
	    RECT 104.6000 35.1000 105.0000 35.2000 ;
	    RECT 103.8000 34.8000 105.0000 35.1000 ;
	    RECT 107.0000 35.1000 107.4000 35.2000 ;
	    RECT 107.0000 34.8000 108.1000 35.1000 ;
	    RECT 102.2000 33.8000 102.6000 34.2000 ;
	    RECT 105.4000 29.8000 105.8000 30.2000 ;
	    RECT 105.4000 29.2000 105.7000 29.8000 ;
	    RECT 107.8000 29.2000 108.1000 34.8000 ;
	    RECT 109.4000 34.8000 109.8000 35.2000 ;
	    RECT 109.4000 34.2000 109.7000 34.8000 ;
	    RECT 109.4000 33.8000 109.8000 34.2000 ;
	    RECT 112.6000 33.2000 112.9000 45.8000 ;
	    RECT 117.4000 44.1000 117.8000 44.2000 ;
	    RECT 118.2000 44.1000 118.5000 49.8000 ;
	    RECT 121.4000 48.2000 121.7000 53.8000 ;
	    RECT 127.0000 51.8000 127.4000 52.2000 ;
	    RECT 131.0000 51.8000 131.4000 52.2000 ;
	    RECT 123.0000 50.8000 123.4000 51.2000 ;
	    RECT 126.2000 51.1000 126.6000 51.2000 ;
	    RECT 127.0000 51.1000 127.3000 51.8000 ;
	    RECT 126.2000 50.8000 127.3000 51.1000 ;
	    RECT 123.0000 49.2000 123.3000 50.8000 ;
	    RECT 123.0000 48.8000 123.4000 49.2000 ;
	    RECT 121.4000 47.8000 121.8000 48.2000 ;
	    RECT 119.0000 46.8000 119.4000 47.2000 ;
	    RECT 119.0000 46.2000 119.3000 46.8000 ;
	    RECT 119.0000 45.8000 119.4000 46.2000 ;
	    RECT 123.0000 46.1000 123.4000 46.2000 ;
	    RECT 123.8000 46.1000 124.2000 46.2000 ;
	    RECT 123.0000 45.8000 124.2000 46.1000 ;
	    RECT 126.2000 46.1000 126.6000 46.2000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 126.2000 45.8000 127.4000 46.1000 ;
	    RECT 129.4000 46.1000 129.8000 46.2000 ;
	    RECT 130.2000 46.1000 130.6000 46.2000 ;
	    RECT 129.4000 45.8000 130.6000 46.1000 ;
	    RECT 127.0000 44.8000 127.4000 45.2000 ;
	    RECT 128.6000 45.1000 129.0000 45.2000 ;
	    RECT 127.8000 44.8000 129.0000 45.1000 ;
	    RECT 127.0000 44.2000 127.3000 44.8000 ;
	    RECT 117.4000 43.8000 118.5000 44.1000 ;
	    RECT 123.8000 44.1000 124.2000 44.2000 ;
	    RECT 124.6000 44.1000 125.0000 44.2000 ;
	    RECT 123.8000 43.8000 125.0000 44.1000 ;
	    RECT 126.2000 43.8000 126.6000 44.2000 ;
	    RECT 127.0000 43.8000 127.4000 44.2000 ;
	    RECT 126.2000 43.2000 126.5000 43.8000 ;
	    RECT 126.2000 42.8000 126.6000 43.2000 ;
	    RECT 114.2000 41.8000 114.6000 42.2000 ;
	    RECT 116.6000 41.8000 117.0000 42.2000 ;
	    RECT 125.4000 41.8000 125.8000 42.2000 ;
	    RECT 114.2000 36.2000 114.5000 41.8000 ;
	    RECT 116.6000 40.2000 116.9000 41.8000 ;
	    RECT 120.6000 40.8000 121.0000 41.2000 ;
	    RECT 116.6000 39.8000 117.0000 40.2000 ;
	    RECT 120.6000 39.2000 120.9000 40.8000 ;
	    RECT 125.4000 39.2000 125.7000 41.8000 ;
	    RECT 120.6000 38.8000 121.0000 39.2000 ;
	    RECT 125.4000 38.8000 125.8000 39.2000 ;
	    RECT 119.8000 37.8000 120.2000 38.2000 ;
	    RECT 123.8000 38.1000 124.2000 38.2000 ;
	    RECT 124.6000 38.1000 125.0000 38.2000 ;
	    RECT 123.8000 37.8000 125.0000 38.1000 ;
	    RECT 117.4000 36.8000 117.8000 37.2000 ;
	    RECT 114.2000 35.8000 114.6000 36.2000 ;
	    RECT 112.6000 32.8000 113.0000 33.2000 ;
	    RECT 114.2000 29.2000 114.5000 35.8000 ;
	    RECT 115.8000 34.1000 116.2000 34.2000 ;
	    RECT 116.6000 34.1000 117.0000 34.2000 ;
	    RECT 115.8000 33.8000 117.0000 34.1000 ;
	    RECT 117.4000 31.2000 117.7000 36.8000 ;
	    RECT 119.8000 36.2000 120.1000 37.8000 ;
	    RECT 121.4000 36.8000 121.8000 37.2000 ;
	    RECT 126.2000 36.8000 126.6000 37.2000 ;
	    RECT 118.2000 36.1000 118.6000 36.2000 ;
	    RECT 119.0000 36.1000 119.4000 36.2000 ;
	    RECT 118.2000 35.8000 119.4000 36.1000 ;
	    RECT 119.8000 35.8000 120.2000 36.2000 ;
	    RECT 118.2000 34.8000 118.6000 35.2000 ;
	    RECT 120.6000 34.8000 121.0000 35.2000 ;
	    RECT 118.2000 34.2000 118.5000 34.8000 ;
	    RECT 120.6000 34.2000 120.9000 34.8000 ;
	    RECT 118.2000 33.8000 118.6000 34.2000 ;
	    RECT 119.0000 33.8000 119.4000 34.2000 ;
	    RECT 120.6000 33.8000 121.0000 34.2000 ;
	    RECT 118.2000 33.1000 118.6000 33.2000 ;
	    RECT 119.0000 33.1000 119.3000 33.8000 ;
	    RECT 118.2000 32.8000 119.3000 33.1000 ;
	    RECT 117.4000 30.8000 117.8000 31.2000 ;
	    RECT 121.4000 30.2000 121.7000 36.8000 ;
	    RECT 125.4000 34.8000 125.8000 35.2000 ;
	    RECT 125.4000 34.2000 125.7000 34.8000 ;
	    RECT 125.4000 33.8000 125.8000 34.2000 ;
	    RECT 117.4000 29.8000 117.8000 30.2000 ;
	    RECT 121.4000 29.8000 121.8000 30.2000 ;
	    RECT 117.4000 29.2000 117.7000 29.8000 ;
	    RECT 126.2000 29.2000 126.5000 36.8000 ;
	    RECT 127.8000 36.2000 128.1000 44.8000 ;
	    RECT 130.2000 44.1000 130.6000 44.2000 ;
	    RECT 131.0000 44.1000 131.3000 51.8000 ;
	    RECT 135.0000 48.2000 135.3000 53.8000 ;
	    RECT 138.2000 53.1000 138.6000 53.2000 ;
	    RECT 138.2000 52.8000 139.3000 53.1000 ;
	    RECT 139.0000 48.2000 139.3000 52.8000 ;
	    RECT 142.2000 49.2000 142.5000 54.8000 ;
	    RECT 143.8000 53.2000 144.1000 73.8000 ;
	    RECT 144.6000 69.2000 144.9000 84.8000 ;
	    RECT 155.0000 83.1000 155.4000 88.9000 ;
	    RECT 159.0000 86.8000 159.4000 87.2000 ;
	    RECT 157.4000 85.8000 157.8000 86.2000 ;
	    RECT 147.0000 80.8000 147.4000 81.2000 ;
	    RECT 146.2000 76.8000 146.6000 77.2000 ;
	    RECT 146.2000 76.2000 146.5000 76.8000 ;
	    RECT 146.2000 75.8000 146.6000 76.2000 ;
	    RECT 147.0000 75.2000 147.3000 80.8000 ;
	    RECT 147.0000 74.8000 147.4000 75.2000 ;
	    RECT 151.8000 75.1000 152.2000 75.2000 ;
	    RECT 152.6000 75.1000 153.0000 75.2000 ;
	    RECT 151.8000 74.8000 153.0000 75.1000 ;
	    RECT 147.8000 73.8000 148.2000 74.2000 ;
	    RECT 149.4000 73.8000 149.8000 74.2000 ;
	    RECT 151.8000 74.1000 152.2000 74.2000 ;
	    RECT 152.6000 74.1000 153.0000 74.2000 ;
	    RECT 151.8000 73.8000 153.0000 74.1000 ;
	    RECT 147.8000 73.2000 148.1000 73.8000 ;
	    RECT 149.4000 73.2000 149.7000 73.8000 ;
	    RECT 145.4000 73.1000 145.8000 73.2000 ;
	    RECT 146.2000 73.1000 146.6000 73.2000 ;
	    RECT 145.4000 72.8000 146.6000 73.1000 ;
	    RECT 147.8000 72.8000 148.2000 73.2000 ;
	    RECT 149.4000 72.8000 149.8000 73.2000 ;
	    RECT 153.4000 73.1000 153.8000 75.9000 ;
	    RECT 148.6000 71.8000 149.0000 72.2000 ;
	    RECT 151.0000 71.8000 151.4000 72.2000 ;
	    RECT 155.0000 72.1000 155.4000 77.9000 ;
	    RECT 155.8000 75.8000 156.2000 76.2000 ;
	    RECT 155.8000 75.1000 156.1000 75.8000 ;
	    RECT 155.8000 74.7000 156.2000 75.1000 ;
	    RECT 144.6000 68.8000 145.0000 69.2000 ;
	    RECT 147.0000 66.8000 147.4000 67.2000 ;
	    RECT 147.0000 66.2000 147.3000 66.8000 ;
	    RECT 147.0000 65.8000 147.4000 66.2000 ;
	    RECT 147.8000 63.1000 148.2000 68.9000 ;
	    RECT 148.6000 65.2000 148.9000 71.8000 ;
	    RECT 151.0000 66.2000 151.3000 71.8000 ;
	    RECT 157.4000 69.2000 157.7000 85.8000 ;
	    RECT 159.0000 75.2000 159.3000 86.8000 ;
	    RECT 159.8000 83.1000 160.2000 88.9000 ;
	    RECT 160.6000 87.2000 160.9000 93.8000 ;
	    RECT 161.4000 92.1000 161.8000 97.9000 ;
	    RECT 163.0000 92.2000 163.3000 106.8000 ;
	    RECT 163.8000 103.1000 164.2000 108.9000 ;
	    RECT 165.4000 107.2000 165.7000 112.8000 ;
	    RECT 169.4000 112.1000 169.8000 117.9000 ;
	    RECT 171.0000 111.2000 171.3000 141.8000 ;
	    RECT 171.8000 135.8000 172.2000 136.2000 ;
	    RECT 171.8000 135.2000 172.1000 135.8000 ;
	    RECT 171.8000 134.8000 172.2000 135.2000 ;
	    RECT 171.8000 131.8000 172.2000 132.2000 ;
	    RECT 171.8000 115.2000 172.1000 131.8000 ;
	    RECT 172.6000 121.8000 173.0000 122.2000 ;
	    RECT 171.8000 114.8000 172.2000 115.2000 ;
	    RECT 171.8000 111.8000 172.2000 112.2000 ;
	    RECT 169.4000 110.8000 169.8000 111.2000 ;
	    RECT 171.0000 110.8000 171.4000 111.2000 ;
	    RECT 165.4000 106.8000 165.8000 107.2000 ;
	    RECT 164.6000 105.9000 165.0000 106.3000 ;
	    RECT 164.6000 105.2000 164.9000 105.9000 ;
	    RECT 164.6000 104.8000 165.0000 105.2000 ;
	    RECT 165.4000 103.8000 165.8000 104.2000 ;
	    RECT 164.6000 94.8000 165.0000 95.2000 ;
	    RECT 163.0000 91.8000 163.4000 92.2000 ;
	    RECT 164.6000 89.2000 164.9000 94.8000 ;
	    RECT 165.4000 89.2000 165.7000 103.8000 ;
	    RECT 168.6000 103.1000 169.0000 108.9000 ;
	    RECT 167.8000 98.1000 168.2000 98.2000 ;
	    RECT 168.6000 98.1000 169.0000 98.2000 ;
	    RECT 166.2000 92.1000 166.6000 97.9000 ;
	    RECT 167.8000 97.8000 169.0000 98.1000 ;
	    RECT 169.4000 97.1000 169.7000 110.8000 ;
	    RECT 171.0000 102.1000 171.4000 102.2000 ;
	    RECT 168.6000 96.8000 169.7000 97.1000 ;
	    RECT 170.2000 101.8000 171.4000 102.1000 ;
	    RECT 164.6000 88.8000 165.0000 89.2000 ;
	    RECT 165.4000 88.8000 165.8000 89.2000 ;
	    RECT 160.6000 86.8000 161.0000 87.2000 ;
	    RECT 161.4000 85.1000 161.8000 87.9000 ;
	    RECT 162.2000 87.1000 162.6000 87.2000 ;
	    RECT 163.0000 87.1000 163.4000 87.2000 ;
	    RECT 162.2000 86.8000 163.4000 87.1000 ;
	    RECT 167.0000 87.1000 167.4000 87.2000 ;
	    RECT 167.8000 87.1000 168.2000 87.2000 ;
	    RECT 167.0000 86.8000 168.2000 87.1000 ;
	    RECT 168.6000 86.2000 168.9000 96.8000 ;
	    RECT 169.4000 91.8000 169.8000 92.2000 ;
	    RECT 163.0000 86.1000 163.4000 86.2000 ;
	    RECT 162.2000 85.8000 163.4000 86.1000 ;
	    RECT 167.0000 85.8000 167.4000 86.2000 ;
	    RECT 167.8000 85.8000 168.2000 86.2000 ;
	    RECT 168.6000 85.8000 169.0000 86.2000 ;
	    RECT 162.2000 79.2000 162.5000 85.8000 ;
	    RECT 165.4000 84.8000 165.8000 85.2000 ;
	    RECT 162.2000 78.8000 162.6000 79.2000 ;
	    RECT 159.0000 74.8000 159.4000 75.2000 ;
	    RECT 151.0000 65.8000 151.4000 66.2000 ;
	    RECT 148.6000 64.8000 149.0000 65.2000 ;
	    RECT 152.6000 63.1000 153.0000 68.9000 ;
	    RECT 155.0000 68.8000 155.4000 69.2000 ;
	    RECT 157.4000 68.8000 157.8000 69.2000 ;
	    RECT 153.4000 67.8000 153.8000 68.2000 ;
	    RECT 153.4000 67.2000 153.7000 67.8000 ;
	    RECT 153.4000 66.8000 153.8000 67.2000 ;
	    RECT 154.2000 65.1000 154.6000 67.9000 ;
	    RECT 155.0000 67.2000 155.3000 68.8000 ;
	    RECT 155.0000 66.8000 155.4000 67.2000 ;
	    RECT 155.0000 66.1000 155.4000 66.2000 ;
	    RECT 155.8000 66.1000 156.2000 66.2000 ;
	    RECT 155.0000 65.8000 156.2000 66.1000 ;
	    RECT 158.2000 65.1000 158.6000 67.9000 ;
	    RECT 159.0000 67.2000 159.3000 74.8000 ;
	    RECT 159.8000 72.1000 160.2000 77.9000 ;
	    RECT 163.0000 73.1000 163.4000 75.9000 ;
	    RECT 163.8000 73.8000 164.2000 74.2000 ;
	    RECT 159.0000 66.8000 159.4000 67.2000 ;
	    RECT 159.0000 66.2000 159.3000 66.8000 ;
	    RECT 159.0000 65.8000 159.4000 66.2000 ;
	    RECT 159.8000 63.1000 160.2000 68.9000 ;
	    RECT 163.8000 67.2000 164.1000 73.8000 ;
	    RECT 164.6000 72.1000 165.0000 77.9000 ;
	    RECT 163.8000 66.8000 164.2000 67.2000 ;
	    RECT 160.6000 65.9000 161.0000 66.3000 ;
	    RECT 160.6000 65.2000 160.9000 65.9000 ;
	    RECT 160.6000 64.8000 161.0000 65.2000 ;
	    RECT 164.6000 63.1000 165.0000 68.9000 ;
	    RECT 165.4000 59.2000 165.7000 84.8000 ;
	    RECT 166.2000 78.8000 166.6000 79.2000 ;
	    RECT 166.2000 75.2000 166.5000 78.8000 ;
	    RECT 166.2000 74.8000 166.6000 75.2000 ;
	    RECT 167.0000 69.2000 167.3000 85.8000 ;
	    RECT 167.0000 68.8000 167.4000 69.2000 ;
	    RECT 167.8000 66.2000 168.1000 85.8000 ;
	    RECT 169.4000 79.2000 169.7000 91.8000 ;
	    RECT 170.2000 86.2000 170.5000 101.8000 ;
	    RECT 171.0000 95.1000 171.4000 95.2000 ;
	    RECT 171.8000 95.1000 172.1000 111.8000 ;
	    RECT 171.0000 94.8000 172.1000 95.1000 ;
	    RECT 171.0000 94.1000 171.4000 94.2000 ;
	    RECT 171.8000 94.1000 172.2000 94.2000 ;
	    RECT 171.0000 93.8000 172.2000 94.1000 ;
	    RECT 171.8000 91.8000 172.2000 92.2000 ;
	    RECT 171.0000 89.8000 171.4000 90.2000 ;
	    RECT 170.2000 85.8000 170.6000 86.2000 ;
	    RECT 171.0000 85.2000 171.3000 89.8000 ;
	    RECT 171.8000 89.2000 172.1000 91.8000 ;
	    RECT 172.6000 89.2000 172.9000 121.8000 ;
	    RECT 171.8000 88.8000 172.2000 89.2000 ;
	    RECT 172.6000 88.8000 173.0000 89.2000 ;
	    RECT 172.6000 87.8000 173.0000 88.2000 ;
	    RECT 172.6000 87.2000 172.9000 87.8000 ;
	    RECT 172.6000 86.8000 173.0000 87.2000 ;
	    RECT 171.0000 84.8000 171.4000 85.2000 ;
	    RECT 169.4000 78.8000 169.8000 79.2000 ;
	    RECT 169.4000 72.1000 169.8000 77.9000 ;
	    RECT 170.2000 71.8000 170.6000 72.2000 ;
	    RECT 171.0000 72.1000 171.4000 72.2000 ;
	    RECT 171.8000 72.1000 172.2000 72.2000 ;
	    RECT 171.0000 71.8000 172.2000 72.1000 ;
	    RECT 170.2000 66.2000 170.5000 71.8000 ;
	    RECT 167.8000 65.8000 168.2000 66.2000 ;
	    RECT 170.2000 65.8000 170.6000 66.2000 ;
	    RECT 148.6000 58.8000 149.0000 59.2000 ;
	    RECT 165.4000 58.8000 165.8000 59.2000 ;
	    RECT 148.6000 58.2000 148.9000 58.8000 ;
	    RECT 145.4000 57.8000 145.8000 58.2000 ;
	    RECT 146.2000 57.8000 146.6000 58.2000 ;
	    RECT 148.6000 57.8000 149.0000 58.2000 ;
	    RECT 145.4000 57.2000 145.7000 57.8000 ;
	    RECT 146.2000 57.2000 146.5000 57.8000 ;
	    RECT 145.4000 56.8000 145.8000 57.2000 ;
	    RECT 146.2000 56.8000 146.6000 57.2000 ;
	    RECT 149.4000 55.8000 149.8000 56.2000 ;
	    RECT 154.2000 56.1000 154.6000 56.2000 ;
	    RECT 155.0000 56.1000 155.4000 56.2000 ;
	    RECT 154.2000 55.8000 155.4000 56.1000 ;
	    RECT 159.8000 56.1000 160.2000 56.2000 ;
	    RECT 160.6000 56.1000 161.0000 56.2000 ;
	    RECT 162.2000 56.1000 162.6000 56.2000 ;
	    RECT 159.8000 55.8000 161.0000 56.1000 ;
	    RECT 161.4000 55.8000 162.6000 56.1000 ;
	    RECT 145.4000 55.1000 145.8000 55.2000 ;
	    RECT 146.2000 55.1000 146.6000 55.2000 ;
	    RECT 145.4000 54.8000 146.6000 55.1000 ;
	    RECT 147.8000 53.8000 148.2000 54.2000 ;
	    RECT 143.8000 52.8000 144.2000 53.2000 ;
	    RECT 142.2000 48.8000 142.6000 49.2000 ;
	    RECT 135.0000 47.8000 135.4000 48.2000 ;
	    RECT 139.0000 47.8000 139.4000 48.2000 ;
	    RECT 146.2000 47.8000 146.6000 48.2000 ;
	    RECT 139.0000 47.2000 139.3000 47.8000 ;
	    RECT 146.2000 47.2000 146.5000 47.8000 ;
	    RECT 147.8000 47.2000 148.1000 53.8000 ;
	    RECT 148.6000 52.8000 149.0000 53.2000 ;
	    RECT 148.6000 49.2000 148.9000 52.8000 ;
	    RECT 148.6000 48.8000 149.0000 49.2000 ;
	    RECT 139.0000 46.8000 139.4000 47.2000 ;
	    RECT 140.6000 46.8000 141.0000 47.2000 ;
	    RECT 142.2000 46.8000 142.6000 47.2000 ;
	    RECT 146.2000 47.1000 146.6000 47.2000 ;
	    RECT 147.0000 47.1000 147.4000 47.2000 ;
	    RECT 146.2000 46.8000 147.4000 47.1000 ;
	    RECT 147.8000 46.8000 148.2000 47.2000 ;
	    RECT 136.6000 46.1000 137.0000 46.2000 ;
	    RECT 137.4000 46.1000 137.8000 46.2000 ;
	    RECT 136.6000 45.8000 137.8000 46.1000 ;
	    RECT 130.2000 43.8000 131.3000 44.1000 ;
	    RECT 131.8000 44.8000 132.2000 45.2000 ;
	    RECT 137.4000 44.8000 137.8000 45.2000 ;
	    RECT 131.8000 44.2000 132.1000 44.8000 ;
	    RECT 131.8000 43.8000 132.2000 44.2000 ;
	    RECT 129.4000 42.1000 129.8000 42.2000 ;
	    RECT 130.2000 42.1000 130.6000 42.2000 ;
	    RECT 129.4000 41.8000 130.6000 42.1000 ;
	    RECT 128.6000 40.8000 129.0000 41.2000 ;
	    RECT 128.6000 39.2000 128.9000 40.8000 ;
	    RECT 137.4000 39.2000 137.7000 44.8000 ;
	    RECT 128.6000 38.8000 129.0000 39.2000 ;
	    RECT 137.4000 38.8000 137.8000 39.2000 ;
	    RECT 132.6000 37.1000 133.0000 37.2000 ;
	    RECT 133.4000 37.1000 133.8000 37.2000 ;
	    RECT 132.6000 36.8000 133.8000 37.1000 ;
	    RECT 138.2000 36.8000 138.6000 37.2000 ;
	    RECT 127.8000 35.8000 128.2000 36.2000 ;
	    RECT 134.2000 35.8000 134.6000 36.2000 ;
	    RECT 134.2000 35.2000 134.5000 35.8000 ;
	    RECT 132.6000 34.8000 133.0000 35.2000 ;
	    RECT 134.2000 34.8000 134.6000 35.2000 ;
	    RECT 137.4000 34.8000 137.8000 35.2000 ;
	    RECT 132.6000 34.2000 132.9000 34.8000 ;
	    RECT 132.6000 33.8000 133.0000 34.2000 ;
	    RECT 135.8000 33.8000 136.2000 34.2000 ;
	    RECT 129.4000 32.8000 129.8000 33.2000 ;
	    RECT 129.4000 30.2000 129.7000 32.8000 ;
	    RECT 135.0000 31.8000 135.4000 32.2000 ;
	    RECT 127.8000 29.8000 128.2000 30.2000 ;
	    RECT 129.4000 29.8000 129.8000 30.2000 ;
	    RECT 95.8000 28.8000 96.2000 29.2000 ;
	    RECT 98.2000 28.8000 98.6000 29.2000 ;
	    RECT 99.8000 28.8000 100.2000 29.2000 ;
	    RECT 101.4000 28.8000 101.8000 29.2000 ;
	    RECT 105.4000 28.8000 105.8000 29.2000 ;
	    RECT 107.8000 28.8000 108.2000 29.2000 ;
	    RECT 111.0000 28.8000 111.4000 29.2000 ;
	    RECT 114.2000 28.8000 114.6000 29.2000 ;
	    RECT 117.4000 28.8000 117.8000 29.2000 ;
	    RECT 126.2000 28.8000 126.6000 29.2000 ;
	    RECT 95.0000 27.8000 95.4000 28.2000 ;
	    RECT 95.0000 27.2000 95.3000 27.8000 ;
	    RECT 95.0000 26.8000 95.4000 27.2000 ;
	    RECT 95.0000 25.8000 95.4000 26.2000 ;
	    RECT 95.0000 25.2000 95.3000 25.8000 ;
	    RECT 95.8000 25.2000 96.1000 28.8000 ;
	    RECT 110.2000 27.8000 110.6000 28.2000 ;
	    RECT 110.2000 27.2000 110.5000 27.8000 ;
	    RECT 98.2000 26.8000 98.6000 27.2000 ;
	    RECT 100.6000 26.8000 101.0000 27.2000 ;
	    RECT 106.2000 27.1000 106.6000 27.2000 ;
	    RECT 107.0000 27.1000 107.4000 27.2000 ;
	    RECT 106.2000 26.8000 107.4000 27.1000 ;
	    RECT 110.2000 26.8000 110.6000 27.2000 ;
	    RECT 98.2000 26.2000 98.5000 26.8000 ;
	    RECT 100.6000 26.2000 100.9000 26.8000 ;
	    RECT 98.2000 25.8000 98.6000 26.2000 ;
	    RECT 100.6000 25.8000 101.0000 26.2000 ;
	    RECT 108.6000 26.1000 109.0000 26.2000 ;
	    RECT 108.6000 25.8000 109.7000 26.1000 ;
	    RECT 95.0000 24.8000 95.4000 25.2000 ;
	    RECT 95.8000 24.8000 96.2000 25.2000 ;
	    RECT 94.2000 23.8000 94.6000 24.2000 ;
	    RECT 99.8000 23.8000 100.2000 24.2000 ;
	    RECT 101.4000 23.8000 101.8000 24.2000 ;
	    RECT 108.6000 23.8000 109.0000 24.2000 ;
	    RECT 94.2000 22.2000 94.5000 23.8000 ;
	    RECT 94.2000 21.8000 94.6000 22.2000 ;
	    RECT 91.8000 18.8000 92.2000 19.2000 ;
	    RECT 92.6000 17.1000 93.0000 17.2000 ;
	    RECT 93.4000 17.1000 93.8000 17.2000 ;
	    RECT 92.6000 16.8000 93.8000 17.1000 ;
	    RECT 97.4000 16.8000 97.8000 17.2000 ;
	    RECT 97.4000 16.2000 97.7000 16.8000 ;
	    RECT 88.6000 14.8000 89.7000 15.1000 ;
	    RECT 91.0000 15.8000 91.4000 16.2000 ;
	    RECT 94.2000 15.8000 94.6000 16.2000 ;
	    RECT 97.4000 15.8000 97.8000 16.2000 ;
	    RECT 91.0000 15.2000 91.3000 15.8000 ;
	    RECT 94.2000 15.2000 94.5000 15.8000 ;
	    RECT 91.0000 14.8000 91.4000 15.2000 ;
	    RECT 91.8000 15.1000 92.2000 15.2000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 91.8000 14.8000 93.0000 15.1000 ;
	    RECT 94.2000 14.8000 94.6000 15.2000 ;
	    RECT 87.8000 11.8000 88.2000 12.2000 ;
	    RECT 84.6000 10.8000 85.0000 11.2000 ;
	    RECT 72.6000 8.8000 73.0000 9.2000 ;
	    RECT 75.8000 8.8000 76.2000 9.2000 ;
	    RECT 80.6000 8.8000 81.0000 9.2000 ;
	    RECT 83.8000 8.8000 84.2000 9.2000 ;
	    RECT 80.6000 8.2000 80.9000 8.8000 ;
	    RECT 84.6000 8.2000 84.9000 10.8000 ;
	    RECT 87.8000 9.2000 88.1000 11.8000 ;
	    RECT 87.8000 8.8000 88.2000 9.2000 ;
	    RECT 54.2000 7.8000 54.6000 8.2000 ;
	    RECT 55.0000 7.8000 55.4000 8.2000 ;
	    RECT 58.2000 7.8000 58.6000 8.2000 ;
	    RECT 60.6000 8.1000 61.0000 8.2000 ;
	    RECT 61.4000 8.1000 61.8000 8.2000 ;
	    RECT 60.6000 7.8000 61.8000 8.1000 ;
	    RECT 70.2000 7.8000 70.6000 8.2000 ;
	    RECT 71.0000 7.8000 71.4000 8.2000 ;
	    RECT 75.0000 7.8000 75.4000 8.2000 ;
	    RECT 80.6000 7.8000 81.0000 8.2000 ;
	    RECT 84.6000 7.8000 85.0000 8.2000 ;
	    RECT 54.2000 7.2000 54.5000 7.8000 ;
	    RECT 58.2000 7.2000 58.5000 7.8000 ;
	    RECT 71.0000 7.2000 71.3000 7.8000 ;
	    RECT 75.0000 7.2000 75.3000 7.8000 ;
	    RECT 84.6000 7.2000 84.9000 7.8000 ;
	    RECT 88.6000 7.2000 88.9000 14.8000 ;
	    RECT 90.2000 12.8000 90.6000 13.2000 ;
	    RECT 91.0000 12.8000 91.4000 13.2000 ;
	    RECT 96.6000 12.8000 97.0000 13.2000 ;
	    RECT 90.2000 11.2000 90.5000 12.8000 ;
	    RECT 90.2000 10.8000 90.6000 11.2000 ;
	    RECT 91.0000 9.2000 91.3000 12.8000 ;
	    RECT 96.6000 11.2000 96.9000 12.8000 ;
	    RECT 99.8000 12.1000 100.1000 23.8000 ;
	    RECT 101.4000 19.2000 101.7000 23.8000 ;
	    RECT 108.6000 22.2000 108.9000 23.8000 ;
	    RECT 107.8000 21.8000 108.2000 22.2000 ;
	    RECT 108.6000 21.8000 109.0000 22.2000 ;
	    RECT 107.8000 19.2000 108.1000 21.8000 ;
	    RECT 109.4000 19.2000 109.7000 25.8000 ;
	    RECT 111.0000 21.2000 111.3000 28.8000 ;
	    RECT 127.8000 28.2000 128.1000 29.8000 ;
	    RECT 115.8000 27.8000 116.2000 28.2000 ;
	    RECT 119.0000 28.1000 119.4000 28.2000 ;
	    RECT 119.8000 28.1000 120.2000 28.2000 ;
	    RECT 119.0000 27.8000 120.2000 28.1000 ;
	    RECT 127.8000 27.8000 128.2000 28.2000 ;
	    RECT 115.8000 27.2000 116.1000 27.8000 ;
	    RECT 115.8000 26.8000 116.2000 27.2000 ;
	    RECT 130.2000 26.8000 130.6000 27.2000 ;
	    RECT 135.0000 27.1000 135.3000 31.8000 ;
	    RECT 135.8000 30.2000 136.1000 33.8000 ;
	    RECT 137.4000 33.2000 137.7000 34.8000 ;
	    RECT 137.4000 32.8000 137.8000 33.2000 ;
	    RECT 136.6000 31.8000 137.0000 32.2000 ;
	    RECT 135.8000 29.8000 136.2000 30.2000 ;
	    RECT 136.6000 29.2000 136.9000 31.8000 ;
	    RECT 138.2000 29.2000 138.5000 36.8000 ;
	    RECT 139.0000 35.2000 139.3000 46.8000 ;
	    RECT 140.6000 46.2000 140.9000 46.8000 ;
	    RECT 142.2000 46.2000 142.5000 46.8000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 142.2000 45.8000 142.6000 46.2000 ;
	    RECT 147.8000 45.8000 148.2000 46.2000 ;
	    RECT 141.4000 44.8000 141.8000 45.2000 ;
	    RECT 143.8000 45.1000 144.2000 45.2000 ;
	    RECT 144.6000 45.1000 145.0000 45.2000 ;
	    RECT 143.8000 44.8000 145.0000 45.1000 ;
	    RECT 141.4000 42.2000 141.7000 44.8000 ;
	    RECT 143.0000 44.1000 143.4000 44.2000 ;
	    RECT 145.4000 44.1000 145.8000 44.2000 ;
	    RECT 143.0000 43.8000 145.8000 44.1000 ;
	    RECT 141.4000 41.8000 141.8000 42.2000 ;
	    RECT 144.6000 41.8000 145.0000 42.2000 ;
	    RECT 139.8000 36.8000 140.2000 37.2000 ;
	    RECT 141.4000 36.8000 141.8000 37.2000 ;
	    RECT 142.2000 37.1000 142.6000 37.2000 ;
	    RECT 143.0000 37.1000 143.4000 37.2000 ;
	    RECT 142.2000 36.8000 143.4000 37.1000 ;
	    RECT 139.8000 36.2000 140.1000 36.8000 ;
	    RECT 141.4000 36.2000 141.7000 36.8000 ;
	    RECT 144.6000 36.2000 144.9000 41.8000 ;
	    RECT 147.8000 40.2000 148.1000 45.8000 ;
	    RECT 149.4000 45.2000 149.7000 55.8000 ;
	    RECT 159.8000 54.8000 160.2000 55.2000 ;
	    RECT 154.2000 53.8000 154.6000 54.2000 ;
	    RECT 152.6000 51.8000 153.0000 52.2000 ;
	    RECT 151.0000 45.8000 151.4000 46.2000 ;
	    RECT 151.0000 45.2000 151.3000 45.8000 ;
	    RECT 149.4000 45.1000 149.8000 45.2000 ;
	    RECT 150.2000 45.1000 150.6000 45.2000 ;
	    RECT 149.4000 44.8000 150.6000 45.1000 ;
	    RECT 151.0000 44.8000 151.4000 45.2000 ;
	    RECT 148.6000 43.8000 149.0000 44.2000 ;
	    RECT 150.2000 43.8000 150.6000 44.2000 ;
	    RECT 151.8000 44.1000 152.2000 44.2000 ;
	    RECT 152.6000 44.1000 152.9000 51.8000 ;
	    RECT 153.4000 48.1000 153.8000 48.2000 ;
	    RECT 154.2000 48.1000 154.5000 53.8000 ;
	    RECT 159.8000 53.2000 160.1000 54.8000 ;
	    RECT 159.8000 52.8000 160.2000 53.2000 ;
	    RECT 153.4000 47.8000 154.5000 48.1000 ;
	    RECT 155.8000 51.8000 156.2000 52.2000 ;
	    RECT 155.8000 48.1000 156.1000 51.8000 ;
	    RECT 155.8000 47.8000 156.9000 48.1000 ;
	    RECT 151.8000 43.8000 152.9000 44.1000 ;
	    RECT 154.2000 47.2000 154.5000 47.8000 ;
	    RECT 154.2000 46.8000 154.6000 47.2000 ;
	    RECT 155.8000 46.8000 156.2000 47.2000 ;
	    RECT 148.6000 42.2000 148.9000 43.8000 ;
	    RECT 150.2000 42.2000 150.5000 43.8000 ;
	    RECT 154.2000 42.2000 154.5000 46.8000 ;
	    RECT 155.8000 46.2000 156.1000 46.8000 ;
	    RECT 155.8000 45.8000 156.2000 46.2000 ;
	    RECT 156.6000 44.1000 156.9000 47.8000 ;
	    RECT 158.2000 47.8000 158.6000 48.2000 ;
	    RECT 158.2000 47.2000 158.5000 47.8000 ;
	    RECT 159.8000 47.2000 160.1000 52.8000 ;
	    RECT 161.4000 49.2000 161.7000 55.8000 ;
	    RECT 163.0000 54.8000 163.4000 55.2000 ;
	    RECT 163.8000 55.1000 164.2000 55.2000 ;
	    RECT 164.6000 55.1000 165.0000 55.2000 ;
	    RECT 163.8000 54.8000 165.0000 55.1000 ;
	    RECT 170.2000 54.8000 170.6000 55.2000 ;
	    RECT 163.0000 54.2000 163.3000 54.8000 ;
	    RECT 170.2000 54.2000 170.5000 54.8000 ;
	    RECT 163.0000 53.8000 163.4000 54.2000 ;
	    RECT 169.4000 53.8000 169.8000 54.2000 ;
	    RECT 170.2000 53.8000 170.6000 54.2000 ;
	    RECT 169.4000 53.2000 169.7000 53.8000 ;
	    RECT 169.4000 52.8000 169.8000 53.2000 ;
	    RECT 167.8000 51.8000 168.2000 52.2000 ;
	    RECT 161.4000 48.8000 161.8000 49.2000 ;
	    RECT 158.2000 46.8000 158.6000 47.2000 ;
	    RECT 159.8000 46.8000 160.2000 47.2000 ;
	    RECT 163.0000 46.8000 163.4000 47.2000 ;
	    RECT 157.4000 46.1000 157.8000 46.2000 ;
	    RECT 158.2000 46.1000 158.6000 46.2000 ;
	    RECT 157.4000 45.8000 158.6000 46.1000 ;
	    RECT 159.0000 44.8000 159.4000 45.2000 ;
	    RECT 157.4000 44.1000 157.8000 44.2000 ;
	    RECT 156.6000 43.8000 157.8000 44.1000 ;
	    RECT 159.0000 43.2000 159.3000 44.8000 ;
	    RECT 159.0000 42.8000 159.4000 43.2000 ;
	    RECT 148.6000 41.8000 149.0000 42.2000 ;
	    RECT 150.2000 41.8000 150.6000 42.2000 ;
	    RECT 154.2000 41.8000 154.6000 42.2000 ;
	    RECT 156.6000 41.8000 157.0000 42.2000 ;
	    RECT 148.6000 40.8000 149.0000 41.2000 ;
	    RECT 147.8000 39.8000 148.2000 40.2000 ;
	    RECT 148.6000 39.2000 148.9000 40.8000 ;
	    RECT 156.6000 39.2000 156.9000 41.8000 ;
	    RECT 148.6000 38.8000 149.0000 39.2000 ;
	    RECT 156.6000 38.8000 157.0000 39.2000 ;
	    RECT 146.2000 36.8000 146.6000 37.2000 ;
	    RECT 147.0000 36.8000 147.4000 37.2000 ;
	    RECT 147.8000 37.1000 148.2000 37.2000 ;
	    RECT 148.6000 37.1000 149.0000 37.2000 ;
	    RECT 149.4000 37.1000 149.8000 37.2000 ;
	    RECT 147.8000 36.8000 149.8000 37.1000 ;
	    RECT 155.0000 36.8000 155.4000 37.2000 ;
	    RECT 155.8000 37.1000 156.2000 37.2000 ;
	    RECT 156.6000 37.1000 157.0000 37.2000 ;
	    RECT 155.8000 36.8000 157.0000 37.1000 ;
	    RECT 139.8000 35.8000 140.2000 36.2000 ;
	    RECT 141.4000 35.8000 141.8000 36.2000 ;
	    RECT 144.6000 35.8000 145.0000 36.2000 ;
	    RECT 145.4000 35.8000 145.8000 36.2000 ;
	    RECT 139.0000 34.8000 139.4000 35.2000 ;
	    RECT 141.4000 34.8000 141.8000 35.2000 ;
	    RECT 143.0000 34.8000 143.4000 35.2000 ;
	    RECT 141.4000 34.2000 141.7000 34.8000 ;
	    RECT 143.0000 34.2000 143.3000 34.8000 ;
	    RECT 141.4000 33.8000 141.8000 34.2000 ;
	    RECT 143.0000 33.8000 143.4000 34.2000 ;
	    RECT 143.8000 33.8000 144.2000 34.2000 ;
	    RECT 139.8000 29.8000 140.2000 30.2000 ;
	    RECT 136.6000 28.8000 137.0000 29.2000 ;
	    RECT 138.2000 28.8000 138.6000 29.2000 ;
	    RECT 139.8000 28.2000 140.1000 29.8000 ;
	    RECT 143.8000 29.2000 144.1000 33.8000 ;
	    RECT 144.6000 32.2000 144.9000 35.8000 ;
	    RECT 145.4000 35.2000 145.7000 35.8000 ;
	    RECT 146.2000 35.2000 146.5000 36.8000 ;
	    RECT 147.0000 36.1000 147.3000 36.8000 ;
	    RECT 147.0000 35.8000 148.1000 36.1000 ;
	    RECT 145.4000 34.8000 145.8000 35.2000 ;
	    RECT 146.2000 34.8000 146.6000 35.2000 ;
	    RECT 146.2000 32.8000 146.6000 33.2000 ;
	    RECT 144.6000 31.8000 145.0000 32.2000 ;
	    RECT 143.8000 28.8000 144.2000 29.2000 ;
	    RECT 139.8000 27.8000 140.2000 28.2000 ;
	    RECT 135.0000 26.8000 136.1000 27.1000 ;
	    RECT 130.2000 26.2000 130.5000 26.8000 ;
	    RECT 115.8000 25.8000 116.2000 26.2000 ;
	    RECT 121.4000 26.1000 121.8000 26.2000 ;
	    RECT 122.2000 26.1000 122.6000 26.2000 ;
	    RECT 121.4000 25.8000 122.6000 26.1000 ;
	    RECT 123.0000 26.1000 123.4000 26.2000 ;
	    RECT 123.8000 26.1000 124.2000 26.2000 ;
	    RECT 123.0000 25.8000 124.2000 26.1000 ;
	    RECT 130.2000 25.8000 130.6000 26.2000 ;
	    RECT 131.8000 26.1000 132.2000 26.2000 ;
	    RECT 132.6000 26.1000 133.0000 26.2000 ;
	    RECT 131.8000 25.8000 133.0000 26.1000 ;
	    RECT 135.0000 25.8000 135.4000 26.2000 ;
	    RECT 115.8000 25.2000 116.1000 25.8000 ;
	    RECT 135.0000 25.2000 135.3000 25.8000 ;
	    RECT 135.8000 25.2000 136.1000 26.8000 ;
	    RECT 142.2000 26.8000 142.6000 27.2000 ;
	    RECT 142.2000 26.2000 142.5000 26.8000 ;
	    RECT 142.2000 25.8000 142.6000 26.2000 ;
	    RECT 143.8000 26.1000 144.2000 26.2000 ;
	    RECT 144.6000 26.1000 145.0000 26.2000 ;
	    RECT 143.8000 25.8000 145.0000 26.1000 ;
	    RECT 114.2000 25.1000 114.6000 25.2000 ;
	    RECT 115.0000 25.1000 115.4000 25.2000 ;
	    RECT 114.2000 24.8000 115.4000 25.1000 ;
	    RECT 115.8000 24.8000 116.2000 25.2000 ;
	    RECT 116.6000 24.8000 117.0000 25.2000 ;
	    RECT 123.0000 24.8000 123.4000 25.2000 ;
	    RECT 125.4000 24.8000 125.8000 25.2000 ;
	    RECT 127.0000 24.8000 127.4000 25.2000 ;
	    RECT 132.6000 24.8000 133.0000 25.2000 ;
	    RECT 133.4000 24.8000 133.8000 25.2000 ;
	    RECT 135.0000 24.8000 135.4000 25.2000 ;
	    RECT 135.8000 24.8000 136.2000 25.2000 ;
	    RECT 139.0000 24.8000 139.4000 25.2000 ;
	    RECT 116.6000 22.2000 116.9000 24.8000 ;
	    RECT 123.0000 24.2000 123.3000 24.8000 ;
	    RECT 123.0000 23.8000 123.4000 24.2000 ;
	    RECT 123.8000 23.8000 124.2000 24.2000 ;
	    RECT 123.8000 23.2000 124.1000 23.8000 ;
	    RECT 123.8000 22.8000 124.2000 23.2000 ;
	    RECT 111.8000 21.8000 112.2000 22.2000 ;
	    RECT 116.6000 21.8000 117.0000 22.2000 ;
	    RECT 111.0000 20.8000 111.4000 21.2000 ;
	    RECT 101.4000 18.8000 101.8000 19.2000 ;
	    RECT 107.8000 18.8000 108.2000 19.2000 ;
	    RECT 109.4000 18.8000 109.8000 19.2000 ;
	    RECT 106.2000 17.8000 106.6000 18.2000 ;
	    RECT 101.4000 17.1000 101.8000 17.2000 ;
	    RECT 102.2000 17.1000 102.6000 17.2000 ;
	    RECT 101.4000 16.8000 102.6000 17.1000 ;
	    RECT 103.0000 15.1000 103.4000 15.2000 ;
	    RECT 103.8000 15.1000 104.2000 15.2000 ;
	    RECT 103.0000 14.8000 104.2000 15.1000 ;
	    RECT 104.6000 12.8000 105.0000 13.2000 ;
	    RECT 99.8000 11.8000 100.9000 12.1000 ;
	    RECT 96.6000 10.8000 97.0000 11.2000 ;
	    RECT 100.6000 9.2000 100.9000 11.8000 ;
	    RECT 103.8000 11.8000 104.2000 12.2000 ;
	    RECT 103.8000 9.2000 104.1000 11.8000 ;
	    RECT 104.6000 9.2000 104.9000 12.8000 ;
	    RECT 106.2000 12.2000 106.5000 17.8000 ;
	    RECT 108.6000 16.8000 109.0000 17.2000 ;
	    RECT 107.0000 15.1000 107.4000 15.2000 ;
	    RECT 107.8000 15.1000 108.2000 15.2000 ;
	    RECT 107.0000 14.8000 108.2000 15.1000 ;
	    RECT 108.6000 13.2000 108.9000 16.8000 ;
	    RECT 111.0000 16.2000 111.3000 20.8000 ;
	    RECT 111.8000 19.2000 112.1000 21.8000 ;
	    RECT 124.6000 20.8000 125.0000 21.2000 ;
	    RECT 111.8000 18.8000 112.2000 19.2000 ;
	    RECT 122.2000 19.1000 122.6000 19.2000 ;
	    RECT 123.0000 19.1000 123.4000 19.2000 ;
	    RECT 122.2000 18.8000 123.4000 19.1000 ;
	    RECT 113.4000 17.8000 113.8000 18.2000 ;
	    RECT 123.8000 17.8000 124.2000 18.2000 ;
	    RECT 113.4000 17.2000 113.7000 17.8000 ;
	    RECT 112.6000 16.8000 113.0000 17.2000 ;
	    RECT 113.4000 16.8000 113.8000 17.2000 ;
	    RECT 122.2000 17.1000 122.6000 17.2000 ;
	    RECT 123.0000 17.1000 123.4000 17.2000 ;
	    RECT 122.2000 16.8000 123.4000 17.1000 ;
	    RECT 111.0000 15.8000 111.4000 16.2000 ;
	    RECT 109.4000 15.1000 109.8000 15.2000 ;
	    RECT 110.2000 15.1000 110.6000 15.2000 ;
	    RECT 109.4000 14.8000 110.6000 15.1000 ;
	    RECT 112.6000 13.2000 112.9000 16.8000 ;
	    RECT 115.8000 15.8000 116.2000 16.2000 ;
	    RECT 116.6000 15.8000 117.0000 16.2000 ;
	    RECT 119.0000 15.8000 119.4000 16.2000 ;
	    RECT 115.8000 15.2000 116.1000 15.8000 ;
	    RECT 114.2000 15.1000 114.6000 15.2000 ;
	    RECT 114.2000 14.8000 115.3000 15.1000 ;
	    RECT 115.8000 14.8000 116.2000 15.2000 ;
	    RECT 115.0000 14.1000 115.3000 14.8000 ;
	    RECT 116.6000 14.1000 116.9000 15.8000 ;
	    RECT 119.0000 15.2000 119.3000 15.8000 ;
	    RECT 123.8000 15.2000 124.1000 17.8000 ;
	    RECT 124.6000 16.2000 124.9000 20.8000 ;
	    RECT 125.4000 19.2000 125.7000 24.8000 ;
	    RECT 125.4000 18.8000 125.8000 19.2000 ;
	    RECT 127.0000 17.2000 127.3000 24.8000 ;
	    RECT 131.8000 23.8000 132.2000 24.2000 ;
	    RECT 131.0000 18.8000 131.4000 19.2000 ;
	    RECT 131.0000 18.2000 131.3000 18.8000 ;
	    RECT 131.0000 17.8000 131.4000 18.2000 ;
	    RECT 126.2000 16.8000 126.6000 17.2000 ;
	    RECT 127.0000 16.8000 127.4000 17.2000 ;
	    RECT 124.6000 15.8000 125.0000 16.2000 ;
	    RECT 119.0000 14.8000 119.4000 15.2000 ;
	    RECT 123.8000 14.8000 124.2000 15.2000 ;
	    RECT 115.0000 13.8000 116.9000 14.1000 ;
	    RECT 108.6000 12.8000 109.0000 13.2000 ;
	    RECT 109.4000 12.8000 109.8000 13.2000 ;
	    RECT 112.6000 12.8000 113.0000 13.2000 ;
	    RECT 115.0000 12.8000 115.4000 13.2000 ;
	    RECT 118.2000 12.8000 118.6000 13.2000 ;
	    RECT 121.4000 12.8000 121.8000 13.2000 ;
	    RECT 106.2000 11.8000 106.6000 12.2000 ;
	    RECT 109.4000 9.2000 109.7000 12.8000 ;
	    RECT 115.0000 9.2000 115.3000 12.8000 ;
	    RECT 118.2000 11.2000 118.5000 12.8000 ;
	    RECT 121.4000 11.2000 121.7000 12.8000 ;
	    RECT 124.6000 11.8000 125.0000 12.2000 ;
	    RECT 118.2000 10.8000 118.6000 11.2000 ;
	    RECT 119.8000 10.8000 120.2000 11.2000 ;
	    RECT 121.4000 10.8000 121.8000 11.2000 ;
	    RECT 123.8000 10.8000 124.2000 11.2000 ;
	    RECT 119.8000 9.2000 120.1000 10.8000 ;
	    RECT 123.8000 9.2000 124.1000 10.8000 ;
	    RECT 91.0000 8.8000 91.4000 9.2000 ;
	    RECT 99.0000 8.8000 99.4000 9.2000 ;
	    RECT 100.6000 8.8000 101.0000 9.2000 ;
	    RECT 103.0000 8.8000 103.4000 9.2000 ;
	    RECT 103.8000 8.8000 104.2000 9.2000 ;
	    RECT 104.6000 8.8000 105.0000 9.2000 ;
	    RECT 109.4000 8.8000 109.8000 9.2000 ;
	    RECT 110.2000 8.8000 110.6000 9.2000 ;
	    RECT 115.0000 8.8000 115.4000 9.2000 ;
	    RECT 119.8000 8.8000 120.2000 9.2000 ;
	    RECT 123.8000 8.8000 124.2000 9.2000 ;
	    RECT 42.2000 7.1000 42.6000 7.2000 ;
	    RECT 43.0000 7.1000 43.4000 7.2000 ;
	    RECT 42.2000 6.8000 43.4000 7.1000 ;
	    RECT 46.2000 6.8000 46.6000 7.2000 ;
	    RECT 47.8000 6.8000 48.2000 7.2000 ;
	    RECT 54.2000 6.8000 54.6000 7.2000 ;
	    RECT 58.2000 6.8000 58.6000 7.2000 ;
	    RECT 71.0000 6.8000 71.4000 7.2000 ;
	    RECT 75.0000 6.8000 75.4000 7.2000 ;
	    RECT 84.6000 6.8000 85.0000 7.2000 ;
	    RECT 88.6000 6.8000 89.0000 7.2000 ;
	    RECT 92.6000 7.1000 93.0000 7.2000 ;
	    RECT 93.4000 7.1000 93.8000 7.2000 ;
	    RECT 92.6000 6.8000 93.8000 7.1000 ;
	    RECT 95.8000 7.1000 96.2000 7.2000 ;
	    RECT 96.6000 7.1000 97.0000 7.2000 ;
	    RECT 95.8000 6.8000 97.0000 7.1000 ;
	    RECT 47.8000 6.2000 48.1000 6.8000 ;
	    RECT 99.0000 6.2000 99.3000 8.8000 ;
	    RECT 99.8000 7.8000 100.2000 8.2000 ;
	    RECT 99.8000 7.2000 100.1000 7.8000 ;
	    RECT 103.0000 7.2000 103.3000 8.8000 ;
	    RECT 110.2000 7.2000 110.5000 8.8000 ;
	    RECT 124.6000 7.2000 124.9000 11.8000 ;
	    RECT 126.2000 9.2000 126.5000 16.8000 ;
	    RECT 127.0000 16.1000 127.4000 16.2000 ;
	    RECT 127.8000 16.1000 128.2000 16.2000 ;
	    RECT 127.0000 15.8000 128.2000 16.1000 ;
	    RECT 127.0000 14.8000 127.4000 15.2000 ;
	    RECT 129.4000 14.8000 129.8000 15.2000 ;
	    RECT 127.0000 14.1000 127.3000 14.8000 ;
	    RECT 129.4000 14.1000 129.7000 14.8000 ;
	    RECT 127.0000 13.8000 129.7000 14.1000 ;
	    RECT 130.2000 12.8000 130.6000 13.2000 ;
	    RECT 130.2000 12.2000 130.5000 12.8000 ;
	    RECT 130.2000 11.8000 130.6000 12.2000 ;
	    RECT 131.8000 9.2000 132.1000 23.8000 ;
	    RECT 132.6000 23.2000 132.9000 24.8000 ;
	    RECT 132.6000 22.8000 133.0000 23.2000 ;
	    RECT 133.4000 21.2000 133.7000 24.8000 ;
	    RECT 139.0000 24.2000 139.3000 24.8000 ;
	    RECT 135.0000 24.1000 135.4000 24.2000 ;
	    RECT 135.8000 24.1000 136.2000 24.2000 ;
	    RECT 135.0000 23.8000 136.2000 24.1000 ;
	    RECT 139.0000 23.8000 139.4000 24.2000 ;
	    RECT 140.6000 23.8000 141.0000 24.2000 ;
	    RECT 144.6000 23.8000 145.0000 24.2000 ;
	    RECT 133.4000 20.8000 133.8000 21.2000 ;
	    RECT 140.6000 19.2000 140.9000 23.8000 ;
	    RECT 140.6000 18.8000 141.0000 19.2000 ;
	    RECT 143.8000 17.8000 144.2000 18.2000 ;
	    RECT 143.8000 17.2000 144.1000 17.8000 ;
	    RECT 143.8000 16.8000 144.2000 17.2000 ;
	    RECT 134.2000 15.8000 134.6000 16.2000 ;
	    RECT 139.0000 15.8000 139.4000 16.2000 ;
	    RECT 141.4000 16.1000 141.8000 16.2000 ;
	    RECT 142.2000 16.1000 142.6000 16.2000 ;
	    RECT 141.4000 15.8000 142.6000 16.1000 ;
	    RECT 134.2000 15.2000 134.5000 15.8000 ;
	    RECT 134.2000 14.8000 134.6000 15.2000 ;
	    RECT 137.4000 14.1000 137.8000 14.2000 ;
	    RECT 138.2000 14.1000 138.6000 14.2000 ;
	    RECT 137.4000 13.8000 138.6000 14.1000 ;
	    RECT 133.4000 12.8000 133.8000 13.2000 ;
	    RECT 136.6000 12.8000 137.0000 13.2000 ;
	    RECT 133.4000 12.2000 133.7000 12.8000 ;
	    RECT 136.6000 12.2000 136.9000 12.8000 ;
	    RECT 133.4000 11.8000 133.8000 12.2000 ;
	    RECT 136.6000 11.8000 137.0000 12.2000 ;
	    RECT 136.6000 10.8000 137.0000 11.2000 ;
	    RECT 136.6000 9.2000 136.9000 10.8000 ;
	    RECT 138.2000 9.8000 138.6000 10.2000 ;
	    RECT 138.2000 9.2000 138.5000 9.8000 ;
	    RECT 139.0000 9.2000 139.3000 15.8000 ;
	    RECT 142.2000 14.8000 142.6000 15.2000 ;
	    RECT 143.8000 14.8000 144.2000 15.2000 ;
	    RECT 140.6000 14.1000 141.0000 14.2000 ;
	    RECT 141.4000 14.1000 141.8000 14.2000 ;
	    RECT 140.6000 13.8000 141.8000 14.1000 ;
	    RECT 141.4000 10.8000 141.8000 11.2000 ;
	    RECT 139.8000 9.8000 140.2000 10.2000 ;
	    RECT 126.2000 8.8000 126.6000 9.2000 ;
	    RECT 131.8000 8.8000 132.2000 9.2000 ;
	    RECT 133.4000 8.8000 133.8000 9.2000 ;
	    RECT 136.6000 8.8000 137.0000 9.2000 ;
	    RECT 138.2000 8.8000 138.6000 9.2000 ;
	    RECT 139.0000 8.8000 139.4000 9.2000 ;
	    RECT 133.4000 7.2000 133.7000 8.8000 ;
	    RECT 138.2000 7.2000 138.5000 8.8000 ;
	    RECT 139.8000 7.2000 140.1000 9.8000 ;
	    RECT 141.4000 9.2000 141.7000 10.8000 ;
	    RECT 142.2000 10.2000 142.5000 14.8000 ;
	    RECT 143.8000 12.2000 144.1000 14.8000 ;
	    RECT 143.8000 11.8000 144.2000 12.2000 ;
	    RECT 142.2000 9.8000 142.6000 10.2000 ;
	    RECT 141.4000 8.8000 141.8000 9.2000 ;
	    RECT 142.2000 7.2000 142.5000 9.8000 ;
	    RECT 144.6000 9.2000 144.9000 23.8000 ;
	    RECT 146.2000 20.1000 146.5000 32.8000 ;
	    RECT 147.8000 32.2000 148.1000 35.8000 ;
	    RECT 150.2000 34.8000 150.6000 35.2000 ;
	    RECT 151.0000 35.1000 151.4000 35.2000 ;
	    RECT 151.8000 35.1000 152.2000 35.2000 ;
	    RECT 151.0000 34.8000 152.2000 35.1000 ;
	    RECT 154.2000 34.8000 154.6000 35.2000 ;
	    RECT 150.2000 32.2000 150.5000 34.8000 ;
	    RECT 154.2000 34.2000 154.5000 34.8000 ;
	    RECT 154.2000 33.8000 154.6000 34.2000 ;
	    RECT 147.0000 31.8000 147.4000 32.2000 ;
	    RECT 147.8000 31.8000 148.2000 32.2000 ;
	    RECT 149.4000 31.8000 149.8000 32.2000 ;
	    RECT 150.2000 31.8000 150.6000 32.2000 ;
	    RECT 151.8000 31.8000 152.2000 32.2000 ;
	    RECT 147.0000 29.2000 147.3000 31.8000 ;
	    RECT 149.4000 29.2000 149.7000 31.8000 ;
	    RECT 151.8000 29.2000 152.1000 31.8000 ;
	    RECT 155.0000 29.2000 155.3000 36.8000 ;
	    RECT 159.0000 31.8000 159.4000 32.2000 ;
	    RECT 159.0000 30.2000 159.3000 31.8000 ;
	    RECT 159.0000 29.8000 159.4000 30.2000 ;
	    RECT 147.0000 28.8000 147.4000 29.2000 ;
	    RECT 149.4000 28.8000 149.8000 29.2000 ;
	    RECT 151.8000 28.8000 152.2000 29.2000 ;
	    RECT 155.0000 28.8000 155.4000 29.2000 ;
	    RECT 156.6000 28.8000 157.0000 29.2000 ;
	    RECT 156.6000 28.2000 156.9000 28.8000 ;
	    RECT 159.8000 28.2000 160.1000 46.8000 ;
	    RECT 163.0000 46.2000 163.3000 46.8000 ;
	    RECT 167.8000 46.2000 168.1000 51.8000 ;
	    RECT 169.4000 48.2000 169.7000 52.8000 ;
	    RECT 171.0000 48.8000 171.4000 49.2000 ;
	    RECT 171.0000 48.2000 171.3000 48.8000 ;
	    RECT 169.4000 47.8000 169.8000 48.2000 ;
	    RECT 171.0000 47.8000 171.4000 48.2000 ;
	    RECT 163.0000 45.8000 163.4000 46.2000 ;
	    RECT 166.2000 45.8000 166.6000 46.2000 ;
	    RECT 167.0000 45.8000 167.4000 46.2000 ;
	    RECT 167.8000 45.8000 168.2000 46.2000 ;
	    RECT 168.6000 45.8000 169.0000 46.2000 ;
	    RECT 163.8000 44.8000 164.2000 45.2000 ;
	    RECT 165.4000 44.8000 165.8000 45.2000 ;
	    RECT 163.8000 44.2000 164.1000 44.8000 ;
	    RECT 165.4000 44.2000 165.7000 44.8000 ;
	    RECT 166.2000 44.2000 166.5000 45.8000 ;
	    RECT 167.0000 45.2000 167.3000 45.8000 ;
	    RECT 168.6000 45.2000 168.9000 45.8000 ;
	    RECT 167.0000 44.8000 167.4000 45.2000 ;
	    RECT 168.6000 44.8000 169.0000 45.2000 ;
	    RECT 163.8000 43.8000 164.2000 44.2000 ;
	    RECT 165.4000 43.8000 165.8000 44.2000 ;
	    RECT 166.2000 43.8000 166.6000 44.2000 ;
	    RECT 164.6000 42.8000 165.0000 43.2000 ;
	    RECT 163.0000 41.8000 163.4000 42.2000 ;
	    RECT 163.0000 39.2000 163.3000 41.8000 ;
	    RECT 163.8000 40.8000 164.2000 41.2000 ;
	    RECT 163.8000 39.2000 164.1000 40.8000 ;
	    RECT 163.0000 38.8000 163.4000 39.2000 ;
	    RECT 163.8000 38.8000 164.2000 39.2000 ;
	    RECT 163.0000 36.8000 163.4000 37.2000 ;
	    RECT 163.0000 36.2000 163.3000 36.8000 ;
	    RECT 164.6000 36.2000 164.9000 42.8000 ;
	    RECT 165.4000 39.8000 165.8000 40.2000 ;
	    RECT 165.4000 39.2000 165.7000 39.8000 ;
	    RECT 165.4000 38.8000 165.8000 39.2000 ;
	    RECT 166.2000 36.8000 166.6000 37.2000 ;
	    RECT 166.2000 36.2000 166.5000 36.8000 ;
	    RECT 163.0000 35.8000 163.4000 36.2000 ;
	    RECT 164.6000 35.8000 165.0000 36.2000 ;
	    RECT 166.2000 35.8000 166.6000 36.2000 ;
	    RECT 170.2000 36.1000 170.6000 36.2000 ;
	    RECT 171.0000 36.1000 171.4000 36.2000 ;
	    RECT 170.2000 35.8000 171.4000 36.1000 ;
	    RECT 162.2000 35.1000 162.6000 35.2000 ;
	    RECT 163.0000 35.1000 163.4000 35.2000 ;
	    RECT 162.2000 34.8000 163.4000 35.1000 ;
	    RECT 161.4000 33.8000 161.8000 34.2000 ;
	    RECT 156.6000 27.8000 157.0000 28.2000 ;
	    RECT 151.8000 25.8000 152.2000 26.2000 ;
	    RECT 151.8000 25.2000 152.1000 25.8000 ;
	    RECT 147.8000 24.8000 148.2000 25.2000 ;
	    RECT 150.2000 24.8000 150.6000 25.2000 ;
	    RECT 151.8000 24.8000 152.2000 25.2000 ;
	    RECT 155.8000 24.8000 156.2000 25.2000 ;
	    RECT 159.0000 25.1000 159.4000 27.9000 ;
	    RECT 159.8000 27.8000 160.2000 28.2000 ;
	    RECT 147.0000 21.8000 147.4000 22.2000 ;
	    RECT 147.0000 21.2000 147.3000 21.8000 ;
	    RECT 147.0000 20.8000 147.4000 21.2000 ;
	    RECT 146.2000 19.8000 147.3000 20.1000 ;
	    RECT 147.0000 19.2000 147.3000 19.8000 ;
	    RECT 147.0000 18.8000 147.4000 19.2000 ;
	    RECT 147.8000 17.2000 148.1000 24.8000 ;
	    RECT 150.2000 24.2000 150.5000 24.8000 ;
	    RECT 150.2000 23.8000 150.6000 24.2000 ;
	    RECT 152.6000 24.1000 153.0000 24.2000 ;
	    RECT 153.4000 24.1000 153.8000 24.2000 ;
	    RECT 152.6000 23.8000 153.8000 24.1000 ;
	    RECT 149.4000 20.8000 149.8000 21.2000 ;
	    RECT 147.8000 16.8000 148.2000 17.2000 ;
	    RECT 149.4000 16.2000 149.7000 20.8000 ;
	    RECT 155.8000 20.2000 156.1000 24.8000 ;
	    RECT 159.0000 23.8000 159.4000 24.2000 ;
	    RECT 155.8000 19.8000 156.2000 20.2000 ;
	    RECT 159.0000 19.2000 159.3000 23.8000 ;
	    RECT 160.6000 23.1000 161.0000 28.9000 ;
	    RECT 161.4000 27.2000 161.7000 33.8000 ;
	    RECT 161.4000 26.8000 161.8000 27.2000 ;
	    RECT 161.4000 22.1000 161.7000 26.8000 ;
	    RECT 162.2000 26.1000 162.6000 26.2000 ;
	    RECT 163.0000 26.1000 163.4000 26.2000 ;
	    RECT 162.2000 25.8000 163.4000 26.1000 ;
	    RECT 160.6000 21.8000 161.7000 22.1000 ;
	    RECT 162.2000 24.8000 162.6000 25.2000 ;
	    RECT 159.0000 18.8000 159.4000 19.2000 ;
	    RECT 151.0000 16.8000 151.4000 17.2000 ;
	    RECT 159.0000 17.1000 159.4000 17.2000 ;
	    RECT 159.8000 17.1000 160.2000 17.2000 ;
	    RECT 159.0000 16.8000 160.2000 17.1000 ;
	    RECT 149.4000 15.8000 149.8000 16.2000 ;
	    RECT 150.2000 15.8000 150.6000 16.2000 ;
	    RECT 150.2000 15.2000 150.5000 15.8000 ;
	    RECT 148.6000 15.1000 149.0000 15.2000 ;
	    RECT 149.4000 15.1000 149.8000 15.2000 ;
	    RECT 148.6000 14.8000 149.8000 15.1000 ;
	    RECT 150.2000 14.8000 150.6000 15.2000 ;
	    RECT 147.8000 13.8000 148.2000 14.2000 ;
	    RECT 151.0000 14.1000 151.3000 16.8000 ;
	    RECT 152.6000 16.1000 153.0000 16.2000 ;
	    RECT 153.4000 16.1000 153.8000 16.2000 ;
	    RECT 152.6000 15.8000 153.8000 16.1000 ;
	    RECT 159.8000 15.8000 160.2000 16.2000 ;
	    RECT 153.4000 15.1000 153.8000 15.2000 ;
	    RECT 154.2000 15.1000 154.6000 15.2000 ;
	    RECT 153.4000 14.8000 154.6000 15.1000 ;
	    RECT 155.0000 14.8000 155.4000 15.2000 ;
	    RECT 157.4000 14.8000 157.8000 15.2000 ;
	    RECT 158.2000 15.1000 158.6000 15.2000 ;
	    RECT 159.0000 15.1000 159.4000 15.2000 ;
	    RECT 158.2000 14.8000 159.4000 15.1000 ;
	    RECT 150.2000 13.8000 151.3000 14.1000 ;
	    RECT 147.8000 9.2000 148.1000 13.8000 ;
	    RECT 150.2000 9.2000 150.5000 13.8000 ;
	    RECT 152.6000 12.8000 153.0000 13.2000 ;
	    RECT 152.6000 10.2000 152.9000 12.8000 ;
	    RECT 154.2000 10.8000 154.6000 11.2000 ;
	    RECT 152.6000 9.8000 153.0000 10.2000 ;
	    RECT 154.2000 9.2000 154.5000 10.8000 ;
	    RECT 155.0000 10.2000 155.3000 14.8000 ;
	    RECT 155.0000 9.8000 155.4000 10.2000 ;
	    RECT 157.4000 9.2000 157.7000 14.8000 ;
	    RECT 159.8000 14.2000 160.1000 15.8000 ;
	    RECT 159.8000 13.8000 160.2000 14.2000 ;
	    RECT 159.0000 11.8000 159.4000 12.2000 ;
	    RECT 144.6000 8.8000 145.0000 9.2000 ;
	    RECT 146.2000 8.8000 146.6000 9.2000 ;
	    RECT 147.8000 8.8000 148.2000 9.2000 ;
	    RECT 148.6000 8.8000 149.0000 9.2000 ;
	    RECT 150.2000 8.8000 150.6000 9.2000 ;
	    RECT 151.8000 8.8000 152.2000 9.2000 ;
	    RECT 154.2000 8.8000 154.6000 9.2000 ;
	    RECT 155.0000 8.8000 155.4000 9.2000 ;
	    RECT 157.4000 8.8000 157.8000 9.2000 ;
	    RECT 146.2000 7.2000 146.5000 8.8000 ;
	    RECT 148.6000 7.2000 148.9000 8.8000 ;
	    RECT 151.8000 8.2000 152.1000 8.8000 ;
	    RECT 155.0000 8.2000 155.3000 8.8000 ;
	    RECT 151.8000 7.8000 152.2000 8.2000 ;
	    RECT 155.0000 7.8000 155.4000 8.2000 ;
	    RECT 157.4000 8.1000 157.8000 8.2000 ;
	    RECT 158.2000 8.1000 158.6000 8.2000 ;
	    RECT 157.4000 7.8000 158.6000 8.1000 ;
	    RECT 159.0000 7.2000 159.3000 11.8000 ;
	    RECT 160.6000 9.2000 160.9000 21.8000 ;
	    RECT 161.4000 20.8000 161.8000 21.2000 ;
	    RECT 161.4000 16.2000 161.7000 20.8000 ;
	    RECT 162.2000 19.2000 162.5000 24.8000 ;
	    RECT 164.6000 21.2000 164.9000 35.8000 ;
	    RECT 165.4000 35.1000 165.8000 35.2000 ;
	    RECT 166.2000 35.1000 166.6000 35.2000 ;
	    RECT 165.4000 34.8000 166.6000 35.1000 ;
	    RECT 171.8000 34.8000 172.2000 35.2000 ;
	    RECT 171.0000 33.8000 171.4000 34.2000 ;
	    RECT 167.8000 29.1000 168.2000 29.2000 ;
	    RECT 168.6000 29.1000 169.0000 29.2000 ;
	    RECT 165.4000 23.1000 165.8000 28.9000 ;
	    RECT 167.8000 28.8000 169.0000 29.1000 ;
	    RECT 171.0000 28.2000 171.3000 33.8000 ;
	    RECT 171.8000 29.2000 172.1000 34.8000 ;
	    RECT 171.8000 28.8000 172.2000 29.2000 ;
	    RECT 167.8000 28.1000 168.2000 28.2000 ;
	    RECT 168.6000 28.1000 169.0000 28.2000 ;
	    RECT 167.8000 27.8000 169.0000 28.1000 ;
	    RECT 171.0000 27.8000 171.4000 28.2000 ;
	    RECT 171.8000 25.8000 172.2000 26.2000 ;
	    RECT 164.6000 20.8000 165.0000 21.2000 ;
	    RECT 165.4000 19.8000 165.8000 20.2000 ;
	    RECT 162.2000 18.8000 162.6000 19.2000 ;
	    RECT 163.0000 16.8000 163.4000 17.2000 ;
	    RECT 161.4000 15.8000 161.8000 16.2000 ;
	    RECT 163.0000 15.2000 163.3000 16.8000 ;
	    RECT 163.8000 16.1000 164.2000 16.2000 ;
	    RECT 164.6000 16.1000 165.0000 16.2000 ;
	    RECT 163.8000 15.8000 165.0000 16.1000 ;
	    RECT 165.4000 15.2000 165.7000 19.8000 ;
	    RECT 162.2000 14.8000 162.6000 15.2000 ;
	    RECT 163.0000 14.8000 163.4000 15.2000 ;
	    RECT 165.4000 14.8000 165.8000 15.2000 ;
	    RECT 166.2000 14.8000 166.6000 15.2000 ;
	    RECT 162.2000 11.2000 162.5000 14.8000 ;
	    RECT 166.2000 14.2000 166.5000 14.8000 ;
	    RECT 166.2000 13.8000 166.6000 14.2000 ;
	    RECT 169.4000 13.8000 169.8000 14.2000 ;
	    RECT 162.2000 10.8000 162.6000 11.2000 ;
	    RECT 166.2000 9.2000 166.5000 13.8000 ;
	    RECT 169.4000 13.2000 169.7000 13.8000 ;
	    RECT 169.4000 12.8000 169.8000 13.2000 ;
	    RECT 167.0000 9.8000 167.4000 10.2000 ;
	    RECT 167.0000 9.2000 167.3000 9.8000 ;
	    RECT 171.8000 9.2000 172.1000 25.8000 ;
	    RECT 160.6000 8.8000 161.0000 9.2000 ;
	    RECT 166.2000 8.8000 166.6000 9.2000 ;
	    RECT 167.0000 8.8000 167.4000 9.2000 ;
	    RECT 171.8000 8.8000 172.2000 9.2000 ;
	    RECT 99.8000 6.8000 100.2000 7.2000 ;
	    RECT 103.0000 6.8000 103.4000 7.2000 ;
	    RECT 110.2000 6.8000 110.6000 7.2000 ;
	    RECT 111.8000 7.1000 112.2000 7.2000 ;
	    RECT 112.6000 7.1000 113.0000 7.2000 ;
	    RECT 111.8000 6.8000 113.0000 7.1000 ;
	    RECT 116.6000 6.8000 117.0000 7.2000 ;
	    RECT 122.2000 7.1000 122.6000 7.2000 ;
	    RECT 123.0000 7.1000 123.4000 7.2000 ;
	    RECT 122.2000 6.8000 123.4000 7.1000 ;
	    RECT 124.6000 6.8000 125.0000 7.2000 ;
	    RECT 133.4000 6.8000 133.8000 7.2000 ;
	    RECT 135.0000 7.1000 135.4000 7.2000 ;
	    RECT 135.8000 7.1000 136.2000 7.2000 ;
	    RECT 135.0000 6.8000 136.2000 7.1000 ;
	    RECT 138.2000 6.8000 138.6000 7.2000 ;
	    RECT 139.8000 6.8000 140.2000 7.2000 ;
	    RECT 142.2000 6.8000 142.6000 7.2000 ;
	    RECT 146.2000 6.8000 146.6000 7.2000 ;
	    RECT 148.6000 6.8000 149.0000 7.2000 ;
	    RECT 149.4000 6.8000 149.8000 7.2000 ;
	    RECT 159.0000 6.8000 159.4000 7.2000 ;
	    RECT 168.6000 7.1000 169.0000 7.2000 ;
	    RECT 169.4000 7.1000 169.8000 7.2000 ;
	    RECT 168.6000 6.8000 169.8000 7.1000 ;
	    RECT 170.2000 6.9000 170.6000 7.0000 ;
	    RECT 171.0000 6.9000 171.4000 7.0000 ;
	    RECT 116.6000 6.2000 116.9000 6.8000 ;
	    RECT 41.4000 5.8000 41.8000 6.2000 ;
	    RECT 42.2000 5.8000 42.6000 6.2000 ;
	    RECT 47.8000 5.8000 48.2000 6.2000 ;
	    RECT 95.8000 5.8000 96.2000 6.2000 ;
	    RECT 97.4000 6.1000 97.8000 6.2000 ;
	    RECT 98.2000 6.1000 98.6000 6.2000 ;
	    RECT 97.4000 5.8000 98.6000 6.1000 ;
	    RECT 99.0000 5.8000 99.4000 6.2000 ;
	    RECT 100.6000 5.8000 101.0000 6.2000 ;
	    RECT 116.6000 5.8000 117.0000 6.2000 ;
	    RECT 128.6000 6.1000 129.0000 6.2000 ;
	    RECT 129.4000 6.1000 129.8000 6.2000 ;
	    RECT 128.6000 5.8000 129.8000 6.1000 ;
	    RECT 135.8000 5.8000 136.2000 6.2000 ;
	    RECT 42.2000 5.2000 42.5000 5.8000 ;
	    RECT 2.2000 4.8000 2.6000 5.2000 ;
	    RECT 3.0000 5.1000 3.4000 5.2000 ;
	    RECT 3.8000 5.1000 4.2000 5.2000 ;
	    RECT 3.0000 4.8000 4.2000 5.1000 ;
	    RECT 7.0000 5.1000 7.4000 5.2000 ;
	    RECT 7.8000 5.1000 8.2000 5.2000 ;
	    RECT 7.0000 4.8000 8.2000 5.1000 ;
	    RECT 17.4000 4.8000 17.8000 5.2000 ;
	    RECT 27.8000 4.8000 28.2000 5.2000 ;
	    RECT 34.2000 5.1000 34.6000 5.2000 ;
	    RECT 35.0000 5.1000 35.4000 5.2000 ;
	    RECT 34.2000 4.8000 35.4000 5.1000 ;
	    RECT 37.4000 4.8000 37.8000 5.2000 ;
	    RECT 41.4000 4.8000 41.8000 5.2000 ;
	    RECT 42.2000 4.8000 42.6000 5.2000 ;
	    RECT 95.8000 5.1000 96.1000 5.8000 ;
	    RECT 100.6000 5.2000 100.9000 5.8000 ;
	    RECT 135.8000 5.2000 136.1000 5.8000 ;
	    RECT 149.4000 5.2000 149.7000 6.8000 ;
	    RECT 170.2000 6.6000 171.4000 6.9000 ;
	    RECT 97.4000 5.1000 97.8000 5.2000 ;
	    RECT 95.8000 4.8000 97.8000 5.1000 ;
	    RECT 100.6000 4.8000 101.0000 5.2000 ;
	    RECT 135.8000 4.8000 136.2000 5.2000 ;
	    RECT 149.4000 4.8000 149.8000 5.2000 ;
	    RECT 17.4000 4.2000 17.7000 4.8000 ;
	    RECT 17.4000 3.8000 17.8000 4.2000 ;
	    RECT 27.8000 2.2000 28.1000 4.8000 ;
	    RECT 41.4000 4.2000 41.7000 4.8000 ;
	    RECT 41.4000 3.8000 41.8000 4.2000 ;
	    RECT 27.8000 1.8000 28.2000 2.2000 ;
	    RECT 44.6000 2.1000 45.0000 2.2000 ;
	    RECT 45.4000 2.1000 45.8000 2.2000 ;
	    RECT 44.6000 1.8000 45.8000 2.1000 ;
         LAYER metal3 ;
	    RECT 90.2000 156.8000 90.6000 157.2000 ;
	    RECT 139.8000 157.1000 140.2000 157.2000 ;
	    RECT 147.8000 157.1000 148.2000 157.2000 ;
	    RECT 151.0000 157.1000 151.4000 157.2000 ;
	    RECT 159.0000 157.1000 159.4000 157.2000 ;
	    RECT 139.8000 156.8000 148.2000 157.1000 ;
	    RECT 150.2000 156.8000 159.4000 157.1000 ;
	    RECT 62.2000 156.1000 62.6000 156.2000 ;
	    RECT 70.2000 156.1000 70.6000 156.2000 ;
	    RECT 62.2000 155.8000 70.6000 156.1000 ;
	    RECT 75.8000 156.1000 76.2000 156.2000 ;
	    RECT 79.0000 156.1000 79.4000 156.2000 ;
	    RECT 90.2000 156.1000 90.5000 156.8000 ;
	    RECT 75.8000 155.8000 90.5000 156.1000 ;
	    RECT 97.4000 156.1000 97.8000 156.2000 ;
	    RECT 99.8000 156.1000 100.2000 156.2000 ;
	    RECT 97.4000 155.8000 100.2000 156.1000 ;
	    RECT 100.6000 156.1000 101.0000 156.2000 ;
	    RECT 107.0000 156.1000 107.4000 156.2000 ;
	    RECT 100.6000 155.8000 107.4000 156.1000 ;
	    RECT 115.8000 156.1000 116.2000 156.2000 ;
	    RECT 116.6000 156.1000 117.0000 156.2000 ;
	    RECT 129.4000 156.1000 129.8000 156.2000 ;
	    RECT 115.8000 155.8000 117.0000 156.1000 ;
	    RECT 122.2000 155.8000 129.8000 156.1000 ;
	    RECT 143.0000 156.1000 143.4000 156.2000 ;
	    RECT 155.0000 156.1000 155.4000 156.2000 ;
	    RECT 143.0000 155.8000 155.4000 156.1000 ;
	    RECT 39.8000 155.1000 40.2000 155.2000 ;
	    RECT 51.8000 155.1000 52.2000 155.2000 ;
	    RECT 39.8000 154.8000 52.2000 155.1000 ;
	    RECT 55.8000 155.1000 56.2000 155.2000 ;
	    RECT 58.2000 155.1000 58.6000 155.2000 ;
	    RECT 60.6000 155.1000 61.0000 155.2000 ;
	    RECT 64.6000 155.1000 65.0000 155.2000 ;
	    RECT 71.8000 155.1000 72.2000 155.2000 ;
	    RECT 55.8000 154.8000 72.2000 155.1000 ;
	    RECT 77.4000 155.1000 77.8000 155.2000 ;
	    RECT 80.6000 155.1000 81.0000 155.2000 ;
	    RECT 93.4000 155.1000 93.8000 155.2000 ;
	    RECT 109.4000 155.1000 109.8000 155.2000 ;
	    RECT 77.4000 154.8000 109.8000 155.1000 ;
	    RECT 116.6000 155.1000 117.0000 155.2000 ;
	    RECT 122.2000 155.1000 122.5000 155.8000 ;
	    RECT 116.6000 154.8000 122.5000 155.1000 ;
	    RECT 123.0000 155.1000 123.4000 155.2000 ;
	    RECT 123.8000 155.1000 124.2000 155.2000 ;
	    RECT 123.0000 154.8000 124.2000 155.1000 ;
	    RECT 129.4000 155.1000 129.8000 155.2000 ;
	    RECT 131.0000 155.1000 131.4000 155.2000 ;
	    RECT 129.4000 154.8000 131.4000 155.1000 ;
	    RECT 131.8000 155.1000 132.2000 155.2000 ;
	    RECT 132.6000 155.1000 133.0000 155.2000 ;
	    RECT 131.8000 154.8000 133.0000 155.1000 ;
	    RECT 138.2000 155.1000 138.6000 155.2000 ;
	    RECT 141.4000 155.1000 141.8000 155.2000 ;
	    RECT 138.2000 154.8000 141.8000 155.1000 ;
	    RECT 147.0000 155.1000 147.4000 155.2000 ;
	    RECT 147.8000 155.1000 148.2000 155.2000 ;
	    RECT 147.0000 154.8000 148.2000 155.1000 ;
	    RECT 149.4000 155.1000 149.8000 155.2000 ;
	    RECT 151.8000 155.1000 152.2000 155.2000 ;
	    RECT 149.4000 154.8000 152.2000 155.1000 ;
	    RECT 159.8000 155.1000 160.2000 155.2000 ;
	    RECT 159.8000 154.8000 164.9000 155.1000 ;
	    RECT 164.6000 154.2000 164.9000 154.8000 ;
	    RECT 9.4000 154.1000 9.8000 154.2000 ;
	    RECT 12.6000 154.1000 13.0000 154.2000 ;
	    RECT 16.6000 154.1000 17.0000 154.2000 ;
	    RECT 18.2000 154.1000 18.6000 154.2000 ;
	    RECT 9.4000 153.8000 18.6000 154.1000 ;
	    RECT 22.2000 154.1000 22.6000 154.2000 ;
	    RECT 25.4000 154.1000 25.8000 154.2000 ;
	    RECT 22.2000 153.8000 25.8000 154.1000 ;
	    RECT 28.6000 154.1000 29.0000 154.2000 ;
	    RECT 31.8000 154.1000 32.2000 154.2000 ;
	    RECT 28.6000 153.8000 32.2000 154.1000 ;
	    RECT 35.0000 154.1000 35.4000 154.2000 ;
	    RECT 36.6000 154.1000 37.0000 154.2000 ;
	    RECT 35.0000 153.8000 37.0000 154.1000 ;
	    RECT 38.2000 154.1000 38.6000 154.2000 ;
	    RECT 42.2000 154.1000 42.6000 154.2000 ;
	    RECT 44.6000 154.1000 45.0000 154.2000 ;
	    RECT 38.2000 153.8000 45.0000 154.1000 ;
	    RECT 47.8000 154.1000 48.2000 154.2000 ;
	    RECT 49.4000 154.1000 49.8000 154.2000 ;
	    RECT 47.8000 153.8000 49.8000 154.1000 ;
	    RECT 85.4000 154.1000 85.8000 154.2000 ;
	    RECT 94.2000 154.1000 94.6000 154.2000 ;
	    RECT 85.4000 153.8000 94.6000 154.1000 ;
	    RECT 96.6000 154.1000 97.0000 154.2000 ;
	    RECT 109.4000 154.1000 109.8000 154.2000 ;
	    RECT 111.8000 154.1000 112.2000 154.2000 ;
	    RECT 96.6000 153.8000 112.2000 154.1000 ;
	    RECT 114.2000 154.1000 114.6000 154.2000 ;
	    RECT 115.0000 154.1000 115.4000 154.2000 ;
	    RECT 118.2000 154.1000 118.6000 154.2000 ;
	    RECT 114.2000 153.8000 118.6000 154.1000 ;
	    RECT 123.0000 154.1000 123.4000 154.2000 ;
	    RECT 139.0000 154.1000 139.4000 154.2000 ;
	    RECT 123.0000 153.8000 139.4000 154.1000 ;
	    RECT 141.4000 154.1000 141.8000 154.2000 ;
	    RECT 142.2000 154.1000 142.6000 154.2000 ;
	    RECT 141.4000 153.8000 142.6000 154.1000 ;
	    RECT 151.0000 154.1000 151.4000 154.2000 ;
	    RECT 155.0000 154.1000 155.4000 154.2000 ;
	    RECT 151.0000 153.8000 155.4000 154.1000 ;
	    RECT 164.6000 153.8000 165.0000 154.2000 ;
	    RECT 40.6000 153.2000 40.9000 153.8000 ;
	    RECT 33.4000 153.1000 33.8000 153.2000 ;
	    RECT 40.6000 153.1000 41.0000 153.2000 ;
	    RECT 33.4000 152.8000 41.0000 153.1000 ;
	    RECT 87.0000 152.8000 87.4000 153.2000 ;
	    RECT 91.0000 153.1000 91.4000 153.2000 ;
	    RECT 96.6000 153.1000 96.9000 153.8000 ;
	    RECT 91.0000 152.8000 96.9000 153.1000 ;
	    RECT 98.2000 153.1000 98.6000 153.2000 ;
	    RECT 99.8000 153.1000 100.2000 153.2000 ;
	    RECT 109.4000 153.1000 109.8000 153.2000 ;
	    RECT 98.2000 152.8000 109.8000 153.1000 ;
	    RECT 122.2000 153.1000 122.6000 153.2000 ;
	    RECT 125.4000 153.1000 125.8000 153.2000 ;
	    RECT 122.2000 152.8000 125.8000 153.1000 ;
	    RECT 130.2000 153.1000 130.6000 153.2000 ;
	    RECT 131.0000 153.1000 131.4000 153.2000 ;
	    RECT 130.2000 152.8000 131.4000 153.1000 ;
	    RECT 131.8000 153.1000 132.2000 153.2000 ;
	    RECT 132.6000 153.1000 133.0000 153.2000 ;
	    RECT 143.8000 153.1000 144.2000 153.2000 ;
	    RECT 147.0000 153.1000 147.4000 153.2000 ;
	    RECT 152.6000 153.1000 153.0000 153.2000 ;
	    RECT 131.8000 152.8000 133.0000 153.1000 ;
	    RECT 134.2000 152.8000 153.0000 153.1000 ;
	    RECT 155.0000 153.1000 155.4000 153.2000 ;
	    RECT 161.4000 153.1000 161.8000 153.2000 ;
	    RECT 155.0000 152.8000 161.8000 153.1000 ;
	    RECT 87.0000 152.2000 87.3000 152.8000 ;
	    RECT 134.2000 152.2000 134.5000 152.8000 ;
	    RECT 46.2000 152.1000 46.6000 152.2000 ;
	    RECT 51.8000 152.1000 52.2000 152.2000 ;
	    RECT 46.2000 151.8000 52.2000 152.1000 ;
	    RECT 52.6000 152.1000 53.0000 152.2000 ;
	    RECT 55.0000 152.1000 55.4000 152.2000 ;
	    RECT 52.6000 151.8000 55.4000 152.1000 ;
	    RECT 87.0000 151.8000 87.4000 152.2000 ;
	    RECT 93.4000 152.1000 93.8000 152.2000 ;
	    RECT 96.6000 152.1000 97.0000 152.2000 ;
	    RECT 93.4000 151.8000 97.0000 152.1000 ;
	    RECT 98.2000 152.1000 98.6000 152.2000 ;
	    RECT 100.6000 152.1000 101.0000 152.2000 ;
	    RECT 98.2000 151.8000 101.0000 152.1000 ;
	    RECT 103.8000 152.1000 104.2000 152.2000 ;
	    RECT 104.6000 152.1000 105.0000 152.2000 ;
	    RECT 103.8000 151.8000 105.0000 152.1000 ;
	    RECT 106.2000 151.8000 106.6000 152.2000 ;
	    RECT 122.2000 152.1000 122.6000 152.2000 ;
	    RECT 123.8000 152.1000 124.2000 152.2000 ;
	    RECT 122.2000 151.8000 124.2000 152.1000 ;
	    RECT 134.2000 151.8000 134.6000 152.2000 ;
	    RECT 137.4000 152.1000 137.8000 152.2000 ;
	    RECT 144.6000 152.1000 145.0000 152.2000 ;
	    RECT 137.4000 151.8000 145.0000 152.1000 ;
	    RECT 153.4000 152.1000 153.8000 152.2000 ;
	    RECT 160.6000 152.1000 161.0000 152.2000 ;
	    RECT 153.4000 151.8000 161.0000 152.1000 ;
	    RECT 106.2000 151.2000 106.5000 151.8000 ;
	    RECT 50.2000 151.1000 50.6000 151.2000 ;
	    RECT 57.4000 151.1000 57.8000 151.2000 ;
	    RECT 50.2000 150.8000 57.8000 151.1000 ;
	    RECT 87.0000 151.1000 87.4000 151.2000 ;
	    RECT 95.8000 151.1000 96.2000 151.2000 ;
	    RECT 87.0000 150.8000 96.2000 151.1000 ;
	    RECT 99.0000 151.1000 99.4000 151.2000 ;
	    RECT 101.4000 151.1000 101.8000 151.2000 ;
	    RECT 99.0000 150.8000 101.8000 151.1000 ;
	    RECT 106.2000 150.8000 106.6000 151.2000 ;
	    RECT 127.0000 151.1000 127.4000 151.2000 ;
	    RECT 137.4000 151.1000 137.8000 151.2000 ;
	    RECT 127.0000 150.8000 137.8000 151.1000 ;
	    RECT 148.6000 151.1000 149.0000 151.2000 ;
	    RECT 154.2000 151.1000 154.6000 151.2000 ;
	    RECT 159.8000 151.1000 160.2000 151.2000 ;
	    RECT 148.6000 150.8000 160.2000 151.1000 ;
	    RECT 87.8000 150.1000 88.2000 150.2000 ;
	    RECT 91.0000 150.1000 91.4000 150.2000 ;
	    RECT 87.8000 149.8000 91.4000 150.1000 ;
	    RECT 117.4000 150.1000 117.8000 150.2000 ;
	    RECT 119.0000 150.1000 119.4000 150.2000 ;
	    RECT 117.4000 149.8000 119.4000 150.1000 ;
	    RECT 119.8000 150.1000 120.2000 150.2000 ;
	    RECT 146.2000 150.1000 146.6000 150.2000 ;
	    RECT 119.8000 149.8000 146.6000 150.1000 ;
	    RECT 6.2000 149.1000 6.6000 149.2000 ;
	    RECT 7.0000 149.1000 7.4000 149.2000 ;
	    RECT 6.2000 148.8000 7.4000 149.1000 ;
	    RECT 73.4000 149.1000 73.8000 149.2000 ;
	    RECT 76.6000 149.1000 77.0000 149.2000 ;
	    RECT 73.4000 148.8000 77.0000 149.1000 ;
	    RECT 77.4000 149.1000 77.8000 149.2000 ;
	    RECT 79.8000 149.1000 80.2000 149.2000 ;
	    RECT 91.0000 149.1000 91.4000 149.2000 ;
	    RECT 77.4000 148.8000 91.4000 149.1000 ;
	    RECT 102.2000 149.1000 102.6000 149.2000 ;
	    RECT 123.8000 149.1000 124.2000 149.2000 ;
	    RECT 136.6000 149.1000 137.0000 149.2000 ;
	    RECT 157.4000 149.1000 157.8000 149.2000 ;
	    RECT 102.2000 148.8000 157.8000 149.1000 ;
	    RECT 11.8000 148.1000 12.2000 148.2000 ;
	    RECT 19.0000 148.1000 19.4000 148.2000 ;
	    RECT 11.8000 147.8000 19.4000 148.1000 ;
	    RECT 44.6000 148.1000 45.0000 148.2000 ;
	    RECT 46.2000 148.1000 46.6000 148.2000 ;
	    RECT 44.6000 147.8000 46.6000 148.1000 ;
	    RECT 67.0000 147.8000 67.4000 148.2000 ;
	    RECT 72.6000 148.1000 73.0000 148.2000 ;
	    RECT 79.0000 148.1000 79.4000 148.2000 ;
	    RECT 82.2000 148.1000 82.6000 148.2000 ;
	    RECT 72.6000 147.8000 82.6000 148.1000 ;
	    RECT 86.2000 147.8000 86.6000 148.2000 ;
	    RECT 89.4000 147.8000 89.8000 148.2000 ;
	    RECT 91.0000 148.1000 91.3000 148.8000 ;
	    RECT 95.0000 148.1000 95.4000 148.2000 ;
	    RECT 95.8000 148.1000 96.2000 148.2000 ;
	    RECT 91.0000 147.8000 96.2000 148.1000 ;
	    RECT 96.6000 148.1000 97.0000 148.2000 ;
	    RECT 103.0000 148.1000 103.4000 148.2000 ;
	    RECT 96.6000 147.8000 103.4000 148.1000 ;
	    RECT 110.2000 148.1000 110.6000 148.2000 ;
	    RECT 116.6000 148.1000 117.0000 148.2000 ;
	    RECT 121.4000 148.1000 121.8000 148.2000 ;
	    RECT 128.6000 148.1000 129.0000 148.2000 ;
	    RECT 110.2000 147.8000 129.0000 148.1000 ;
	    RECT 161.4000 148.1000 161.8000 148.2000 ;
	    RECT 169.4000 148.1000 169.8000 148.2000 ;
	    RECT 161.4000 147.8000 169.8000 148.1000 ;
	    RECT 3.8000 146.8000 4.2000 147.2000 ;
	    RECT 5.4000 147.1000 5.8000 147.2000 ;
	    RECT 7.0000 147.1000 7.4000 147.2000 ;
	    RECT 5.4000 146.8000 7.4000 147.1000 ;
	    RECT 15.8000 146.8000 16.2000 147.2000 ;
	    RECT 17.4000 147.1000 17.8000 147.2000 ;
	    RECT 18.2000 147.1000 18.6000 147.2000 ;
	    RECT 17.4000 146.8000 18.6000 147.1000 ;
	    RECT 21.4000 147.1000 21.8000 147.2000 ;
	    RECT 24.6000 147.1000 25.0000 147.2000 ;
	    RECT 21.4000 146.8000 25.0000 147.1000 ;
	    RECT 31.8000 147.1000 32.2000 147.2000 ;
	    RECT 35.0000 147.1000 35.4000 147.2000 ;
	    RECT 31.8000 146.8000 35.4000 147.1000 ;
	    RECT 53.4000 147.1000 53.8000 147.2000 ;
	    RECT 58.2000 147.1000 58.6000 147.2000 ;
	    RECT 64.6000 147.1000 65.0000 147.2000 ;
	    RECT 65.4000 147.1000 65.8000 147.2000 ;
	    RECT 53.4000 146.8000 58.6000 147.1000 ;
	    RECT 63.8000 146.8000 65.8000 147.1000 ;
	    RECT 67.0000 147.1000 67.3000 147.8000 ;
	    RECT 68.6000 147.1000 69.0000 147.2000 ;
	    RECT 67.0000 146.8000 69.0000 147.1000 ;
	    RECT 74.2000 147.1000 74.6000 147.2000 ;
	    RECT 75.8000 147.1000 76.2000 147.2000 ;
	    RECT 79.0000 147.1000 79.4000 147.2000 ;
	    RECT 85.4000 147.1000 85.8000 147.2000 ;
	    RECT 74.2000 146.8000 75.3000 147.1000 ;
	    RECT 75.8000 146.8000 85.8000 147.1000 ;
	    RECT 86.2000 147.1000 86.5000 147.8000 ;
	    RECT 89.4000 147.1000 89.7000 147.8000 ;
	    RECT 86.2000 146.8000 89.7000 147.1000 ;
	    RECT 90.2000 147.1000 90.6000 147.2000 ;
	    RECT 92.6000 147.1000 93.0000 147.2000 ;
	    RECT 99.8000 147.1000 100.2000 147.2000 ;
	    RECT 90.2000 146.8000 100.2000 147.1000 ;
	    RECT 109.4000 147.1000 109.8000 147.2000 ;
	    RECT 112.6000 147.1000 113.0000 147.2000 ;
	    RECT 114.2000 147.1000 114.6000 147.2000 ;
	    RECT 109.4000 146.8000 114.6000 147.1000 ;
	    RECT 115.8000 147.1000 116.2000 147.2000 ;
	    RECT 120.6000 147.1000 121.0000 147.2000 ;
	    RECT 115.8000 146.8000 121.0000 147.1000 ;
	    RECT 125.4000 147.1000 125.8000 147.2000 ;
	    RECT 131.8000 147.1000 132.2000 147.2000 ;
	    RECT 125.4000 146.8000 132.2000 147.1000 ;
	    RECT 142.2000 147.1000 142.6000 147.2000 ;
	    RECT 144.6000 147.1000 145.0000 147.2000 ;
	    RECT 142.2000 146.8000 145.0000 147.1000 ;
	    RECT 146.2000 147.1000 146.6000 147.2000 ;
	    RECT 155.0000 147.1000 155.4000 147.2000 ;
	    RECT 146.2000 146.8000 155.4000 147.1000 ;
	    RECT 165.4000 147.1000 165.8000 147.2000 ;
	    RECT 166.2000 147.1000 166.6000 147.2000 ;
	    RECT 165.4000 146.8000 166.6000 147.1000 ;
	    RECT 3.0000 146.1000 3.4000 146.2000 ;
	    RECT 3.8000 146.1000 4.1000 146.8000 ;
	    RECT 3.0000 145.8000 4.1000 146.1000 ;
	    RECT 4.6000 146.1000 5.0000 146.2000 ;
	    RECT 6.2000 146.1000 6.6000 146.2000 ;
	    RECT 7.8000 146.1000 8.2000 146.2000 ;
	    RECT 4.6000 145.8000 8.2000 146.1000 ;
	    RECT 13.4000 146.1000 13.8000 146.2000 ;
	    RECT 14.2000 146.1000 14.6000 146.2000 ;
	    RECT 15.8000 146.1000 16.1000 146.8000 ;
	    RECT 75.0000 146.2000 75.3000 146.8000 ;
	    RECT 26.2000 146.1000 26.6000 146.2000 ;
	    RECT 27.8000 146.1000 28.2000 146.2000 ;
	    RECT 13.4000 145.8000 28.2000 146.1000 ;
	    RECT 38.2000 146.1000 38.6000 146.2000 ;
	    RECT 39.8000 146.1000 40.2000 146.2000 ;
	    RECT 38.2000 145.8000 40.2000 146.1000 ;
	    RECT 46.2000 145.8000 46.6000 146.2000 ;
	    RECT 50.2000 146.1000 50.6000 146.2000 ;
	    RECT 52.6000 146.1000 53.0000 146.2000 ;
	    RECT 50.2000 145.8000 53.0000 146.1000 ;
	    RECT 75.0000 145.8000 75.4000 146.2000 ;
	    RECT 84.6000 146.1000 85.0000 146.2000 ;
	    RECT 86.2000 146.1000 86.6000 146.2000 ;
	    RECT 84.6000 145.8000 86.6000 146.1000 ;
	    RECT 92.6000 146.1000 93.0000 146.2000 ;
	    RECT 93.4000 146.1000 93.8000 146.2000 ;
	    RECT 92.6000 145.8000 93.8000 146.1000 ;
	    RECT 95.0000 146.1000 95.4000 146.2000 ;
	    RECT 97.4000 146.1000 97.8000 146.2000 ;
	    RECT 95.0000 145.8000 97.8000 146.1000 ;
	    RECT 99.0000 146.1000 99.4000 146.2000 ;
	    RECT 101.4000 146.1000 101.8000 146.2000 ;
	    RECT 99.0000 145.8000 101.8000 146.1000 ;
	    RECT 106.2000 146.1000 106.6000 146.2000 ;
	    RECT 107.0000 146.1000 107.4000 146.2000 ;
	    RECT 111.0000 146.1000 111.4000 146.2000 ;
	    RECT 106.2000 145.8000 111.4000 146.1000 ;
	    RECT 115.0000 146.1000 115.4000 146.2000 ;
	    RECT 125.4000 146.1000 125.8000 146.2000 ;
	    RECT 115.0000 145.8000 125.8000 146.1000 ;
	    RECT 127.0000 145.8000 127.4000 146.2000 ;
	    RECT 132.6000 146.1000 133.0000 146.2000 ;
	    RECT 139.8000 146.1000 140.2000 146.2000 ;
	    RECT 152.6000 146.1000 153.0000 146.2000 ;
	    RECT 132.6000 145.8000 153.0000 146.1000 ;
	    RECT 166.2000 145.8000 166.6000 146.2000 ;
	    RECT 20.6000 145.1000 21.0000 145.2000 ;
	    RECT 31.0000 145.1000 31.4000 145.2000 ;
	    RECT 20.6000 144.8000 31.4000 145.1000 ;
	    RECT 43.8000 145.1000 44.2000 145.2000 ;
	    RECT 46.2000 145.1000 46.5000 145.8000 ;
	    RECT 43.8000 144.8000 46.5000 145.1000 ;
	    RECT 47.8000 145.1000 48.2000 145.2000 ;
	    RECT 55.8000 145.1000 56.2000 145.2000 ;
	    RECT 64.6000 145.1000 65.0000 145.2000 ;
	    RECT 47.8000 144.8000 65.0000 145.1000 ;
	    RECT 89.4000 145.1000 89.8000 145.2000 ;
	    RECT 94.2000 145.1000 94.6000 145.2000 ;
	    RECT 89.4000 144.8000 94.6000 145.1000 ;
	    RECT 107.0000 145.1000 107.4000 145.2000 ;
	    RECT 113.4000 145.1000 113.8000 145.2000 ;
	    RECT 107.0000 144.8000 113.8000 145.1000 ;
	    RECT 115.8000 145.1000 116.2000 145.2000 ;
	    RECT 118.2000 145.1000 118.6000 145.2000 ;
	    RECT 115.8000 144.8000 118.6000 145.1000 ;
	    RECT 119.0000 145.1000 119.4000 145.2000 ;
	    RECT 127.0000 145.1000 127.3000 145.8000 ;
	    RECT 166.2000 145.2000 166.5000 145.8000 ;
	    RECT 119.0000 144.8000 127.3000 145.1000 ;
	    RECT 135.8000 145.1000 136.2000 145.2000 ;
	    RECT 143.0000 145.1000 143.4000 145.2000 ;
	    RECT 158.2000 145.1000 158.6000 145.2000 ;
	    RECT 135.8000 144.8000 143.4000 145.1000 ;
	    RECT 155.8000 144.8000 158.6000 145.1000 ;
	    RECT 166.2000 144.8000 166.6000 145.2000 ;
	    RECT 155.8000 144.2000 156.1000 144.8000 ;
	    RECT 6.2000 144.1000 6.6000 144.2000 ;
	    RECT 7.0000 144.1000 7.4000 144.2000 ;
	    RECT 6.2000 143.8000 7.4000 144.1000 ;
	    RECT 64.6000 144.1000 65.0000 144.2000 ;
	    RECT 78.2000 144.1000 78.6000 144.2000 ;
	    RECT 64.6000 143.8000 78.6000 144.1000 ;
	    RECT 94.2000 144.1000 94.6000 144.2000 ;
	    RECT 94.2000 143.8000 101.7000 144.1000 ;
	    RECT 101.4000 143.2000 101.7000 143.8000 ;
	    RECT 106.2000 143.8000 106.6000 144.2000 ;
	    RECT 109.4000 144.1000 109.8000 144.2000 ;
	    RECT 107.8000 143.8000 109.8000 144.1000 ;
	    RECT 112.6000 144.1000 113.0000 144.2000 ;
	    RECT 120.6000 144.1000 121.0000 144.2000 ;
	    RECT 123.0000 144.1000 123.4000 144.2000 ;
	    RECT 112.6000 143.8000 123.4000 144.1000 ;
	    RECT 131.8000 144.1000 132.2000 144.2000 ;
	    RECT 140.6000 144.1000 141.0000 144.2000 ;
	    RECT 151.0000 144.1000 151.4000 144.2000 ;
	    RECT 131.8000 143.8000 151.4000 144.1000 ;
	    RECT 155.8000 143.8000 156.2000 144.2000 ;
	    RECT 161.4000 144.1000 161.8000 144.2000 ;
	    RECT 167.0000 144.1000 167.4000 144.2000 ;
	    RECT 161.4000 143.8000 167.4000 144.1000 ;
	    RECT 106.2000 143.2000 106.5000 143.8000 ;
	    RECT 107.8000 143.2000 108.1000 143.8000 ;
	    RECT 29.4000 143.1000 29.8000 143.2000 ;
	    RECT 33.4000 143.1000 33.8000 143.2000 ;
	    RECT 29.4000 142.8000 33.8000 143.1000 ;
	    RECT 44.6000 142.8000 45.0000 143.2000 ;
	    RECT 101.4000 142.8000 101.8000 143.2000 ;
	    RECT 106.2000 142.8000 106.6000 143.2000 ;
	    RECT 107.8000 142.8000 108.2000 143.2000 ;
	    RECT 142.2000 143.1000 142.6000 143.2000 ;
	    RECT 157.4000 143.1000 157.8000 143.2000 ;
	    RECT 121.4000 142.8000 157.8000 143.1000 ;
	    RECT 164.6000 143.1000 165.0000 143.2000 ;
	    RECT 167.8000 143.1000 168.2000 143.2000 ;
	    RECT 164.6000 142.8000 168.2000 143.1000 ;
	    RECT 44.6000 142.1000 44.9000 142.8000 ;
	    RECT 79.0000 142.1000 79.4000 142.2000 ;
	    RECT 44.6000 141.8000 79.4000 142.1000 ;
	    RECT 91.0000 142.1000 91.4000 142.2000 ;
	    RECT 100.6000 142.1000 101.0000 142.2000 ;
	    RECT 91.0000 141.8000 101.0000 142.1000 ;
	    RECT 103.0000 142.1000 103.4000 142.2000 ;
	    RECT 121.4000 142.1000 121.7000 142.8000 ;
	    RECT 103.0000 141.8000 121.7000 142.1000 ;
	    RECT 122.2000 142.1000 122.6000 142.2000 ;
	    RECT 128.6000 142.1000 129.0000 142.2000 ;
	    RECT 122.2000 141.8000 129.0000 142.1000 ;
	    RECT 132.6000 142.1000 133.0000 142.2000 ;
	    RECT 139.0000 142.1000 139.4000 142.2000 ;
	    RECT 132.6000 141.8000 139.4000 142.1000 ;
	    RECT 149.4000 142.1000 149.8000 142.2000 ;
	    RECT 161.4000 142.1000 161.8000 142.2000 ;
	    RECT 149.4000 141.8000 161.8000 142.1000 ;
	    RECT 3.0000 141.1000 3.4000 141.2000 ;
	    RECT 8.6000 141.1000 9.0000 141.2000 ;
	    RECT 19.8000 141.1000 20.2000 141.2000 ;
	    RECT 3.0000 140.8000 20.2000 141.1000 ;
	    RECT 88.6000 141.1000 89.0000 141.2000 ;
	    RECT 105.4000 141.1000 105.8000 141.2000 ;
	    RECT 88.6000 140.8000 105.8000 141.1000 ;
	    RECT 128.6000 141.1000 129.0000 141.2000 ;
	    RECT 138.2000 141.1000 138.6000 141.2000 ;
	    RECT 128.6000 140.8000 138.6000 141.1000 ;
	    RECT 143.8000 141.1000 144.2000 141.2000 ;
	    RECT 159.0000 141.1000 159.4000 141.2000 ;
	    RECT 143.8000 140.8000 159.4000 141.1000 ;
	    RECT 2.2000 140.1000 2.6000 140.2000 ;
	    RECT 3.8000 140.1000 4.2000 140.2000 ;
	    RECT 2.2000 139.8000 4.2000 140.1000 ;
	    RECT 37.4000 140.1000 37.8000 140.2000 ;
	    RECT 57.4000 140.1000 57.8000 140.2000 ;
	    RECT 37.4000 139.8000 57.8000 140.1000 ;
	    RECT 99.8000 140.1000 100.2000 140.2000 ;
	    RECT 101.4000 140.1000 101.8000 140.2000 ;
	    RECT 99.8000 139.8000 101.8000 140.1000 ;
	    RECT 113.4000 140.1000 113.8000 140.2000 ;
	    RECT 130.2000 140.1000 130.6000 140.2000 ;
	    RECT 136.6000 140.1000 137.0000 140.2000 ;
	    RECT 147.8000 140.1000 148.2000 140.2000 ;
	    RECT 113.4000 139.8000 148.2000 140.1000 ;
	    RECT 152.6000 140.1000 153.0000 140.2000 ;
	    RECT 155.0000 140.1000 155.4000 140.2000 ;
	    RECT 152.6000 139.8000 155.4000 140.1000 ;
	    RECT 2.2000 138.8000 2.6000 139.2000 ;
	    RECT 23.0000 139.1000 23.4000 139.2000 ;
	    RECT 28.6000 139.1000 29.0000 139.2000 ;
	    RECT 23.0000 138.8000 29.0000 139.1000 ;
	    RECT 99.0000 139.1000 99.4000 139.2000 ;
	    RECT 102.2000 139.1000 102.6000 139.2000 ;
	    RECT 127.8000 139.1000 128.2000 139.2000 ;
	    RECT 135.0000 139.1000 135.4000 139.2000 ;
	    RECT 99.0000 138.8000 102.6000 139.1000 ;
	    RECT 127.0000 138.8000 135.4000 139.1000 ;
	    RECT 139.0000 138.8000 139.4000 139.2000 ;
	    RECT 151.0000 139.1000 151.4000 139.2000 ;
	    RECT 151.0000 138.8000 153.7000 139.1000 ;
	    RECT 2.2000 138.1000 2.5000 138.8000 ;
	    RECT 5.4000 138.1000 5.8000 138.2000 ;
	    RECT 2.2000 137.8000 5.8000 138.1000 ;
	    RECT 13.4000 138.1000 13.8000 138.2000 ;
	    RECT 13.4000 137.8000 26.5000 138.1000 ;
	    RECT 26.2000 137.2000 26.5000 137.8000 ;
	    RECT 56.6000 137.8000 57.0000 138.2000 ;
	    RECT 58.2000 138.1000 58.6000 138.2000 ;
	    RECT 81.4000 138.1000 81.8000 138.2000 ;
	    RECT 95.8000 138.1000 96.2000 138.2000 ;
	    RECT 99.8000 138.1000 100.2000 138.2000 ;
	    RECT 58.2000 137.8000 81.8000 138.1000 ;
	    RECT 92.6000 137.8000 100.2000 138.1000 ;
	    RECT 129.4000 138.1000 129.8000 138.2000 ;
	    RECT 139.0000 138.1000 139.3000 138.8000 ;
	    RECT 129.4000 137.8000 139.3000 138.1000 ;
	    RECT 153.4000 138.2000 153.7000 138.8000 ;
	    RECT 153.4000 137.8000 153.8000 138.2000 ;
	    RECT 157.4000 138.1000 157.8000 138.2000 ;
	    RECT 166.2000 138.1000 166.6000 138.2000 ;
	    RECT 157.4000 137.8000 166.6000 138.1000 ;
	    RECT 4.6000 137.1000 5.0000 137.2000 ;
	    RECT 5.4000 137.1000 5.8000 137.2000 ;
	    RECT 4.6000 136.8000 5.8000 137.1000 ;
	    RECT 11.0000 137.1000 11.4000 137.2000 ;
	    RECT 11.8000 137.1000 12.2000 137.2000 ;
	    RECT 11.0000 136.8000 12.2000 137.1000 ;
	    RECT 12.6000 137.1000 13.0000 137.2000 ;
	    RECT 21.4000 137.1000 21.8000 137.2000 ;
	    RECT 12.6000 136.8000 21.8000 137.1000 ;
	    RECT 26.2000 136.8000 26.6000 137.2000 ;
	    RECT 40.6000 136.8000 41.0000 137.2000 ;
	    RECT 55.0000 136.8000 55.4000 137.2000 ;
	    RECT 56.6000 137.1000 56.9000 137.8000 ;
	    RECT 92.6000 137.2000 92.9000 137.8000 ;
	    RECT 67.8000 137.1000 68.2000 137.2000 ;
	    RECT 56.6000 136.8000 68.2000 137.1000 ;
	    RECT 81.4000 137.1000 81.8000 137.2000 ;
	    RECT 92.6000 137.1000 93.0000 137.2000 ;
	    RECT 81.4000 136.8000 93.0000 137.1000 ;
	    RECT 94.2000 137.1000 94.6000 137.2000 ;
	    RECT 96.6000 137.1000 97.0000 137.2000 ;
	    RECT 126.2000 137.1000 126.6000 137.2000 ;
	    RECT 127.0000 137.1000 127.4000 137.2000 ;
	    RECT 94.2000 136.8000 99.3000 137.1000 ;
	    RECT 126.2000 136.8000 127.4000 137.1000 ;
	    RECT 130.2000 137.1000 130.6000 137.2000 ;
	    RECT 137.4000 137.1000 137.8000 137.2000 ;
	    RECT 150.2000 137.1000 150.6000 137.2000 ;
	    RECT 157.4000 137.1000 157.8000 137.2000 ;
	    RECT 158.2000 137.1000 158.6000 137.2000 ;
	    RECT 130.2000 136.8000 158.6000 137.1000 ;
	    RECT 163.0000 136.8000 163.4000 137.2000 ;
	    RECT 15.0000 136.1000 15.4000 136.2000 ;
	    RECT 15.8000 136.1000 16.2000 136.2000 ;
	    RECT 15.0000 135.8000 16.2000 136.1000 ;
	    RECT 28.6000 136.1000 29.0000 136.2000 ;
	    RECT 30.2000 136.1000 30.6000 136.2000 ;
	    RECT 28.6000 135.8000 30.6000 136.1000 ;
	    RECT 32.6000 136.1000 33.0000 136.2000 ;
	    RECT 33.4000 136.1000 33.8000 136.2000 ;
	    RECT 32.6000 135.8000 33.8000 136.1000 ;
	    RECT 38.2000 136.1000 38.6000 136.2000 ;
	    RECT 40.6000 136.1000 40.9000 136.8000 ;
	    RECT 55.0000 136.2000 55.3000 136.8000 ;
	    RECT 38.2000 135.8000 40.9000 136.1000 ;
	    RECT 49.4000 136.1000 49.8000 136.2000 ;
	    RECT 53.4000 136.1000 53.8000 136.2000 ;
	    RECT 49.4000 135.8000 53.8000 136.1000 ;
	    RECT 55.0000 135.8000 55.4000 136.2000 ;
	    RECT 57.4000 136.1000 57.8000 136.2000 ;
	    RECT 61.4000 136.1000 61.8000 136.2000 ;
	    RECT 57.4000 135.8000 61.8000 136.1000 ;
	    RECT 75.0000 136.1000 75.4000 136.2000 ;
	    RECT 81.4000 136.1000 81.7000 136.8000 ;
	    RECT 99.0000 136.2000 99.3000 136.8000 ;
	    RECT 75.0000 135.8000 81.7000 136.1000 ;
	    RECT 85.4000 136.1000 85.8000 136.2000 ;
	    RECT 94.2000 136.1000 94.6000 136.2000 ;
	    RECT 85.4000 135.8000 94.6000 136.1000 ;
	    RECT 97.4000 135.8000 97.8000 136.2000 ;
	    RECT 99.0000 135.8000 99.4000 136.2000 ;
	    RECT 131.0000 136.1000 131.4000 136.2000 ;
	    RECT 141.4000 136.1000 141.8000 136.2000 ;
	    RECT 151.0000 136.1000 151.4000 136.2000 ;
	    RECT 151.8000 136.1000 152.2000 136.2000 ;
	    RECT 131.0000 135.8000 152.2000 136.1000 ;
	    RECT 159.0000 136.1000 159.4000 136.2000 ;
	    RECT 163.0000 136.1000 163.3000 136.8000 ;
	    RECT 167.8000 136.1000 168.2000 136.2000 ;
	    RECT 159.0000 135.8000 168.2000 136.1000 ;
	    RECT 171.8000 135.8000 172.2000 136.2000 ;
	    RECT 5.4000 135.1000 5.8000 135.2000 ;
	    RECT 11.8000 135.1000 12.2000 135.2000 ;
	    RECT 5.4000 134.8000 12.2000 135.1000 ;
	    RECT 18.2000 135.1000 18.6000 135.2000 ;
	    RECT 29.4000 135.1000 29.8000 135.2000 ;
	    RECT 18.2000 134.8000 29.8000 135.1000 ;
	    RECT 39.8000 135.1000 40.2000 135.2000 ;
	    RECT 43.8000 135.1000 44.2000 135.2000 ;
	    RECT 47.0000 135.1000 47.4000 135.2000 ;
	    RECT 50.2000 135.1000 50.6000 135.2000 ;
	    RECT 39.8000 134.8000 50.6000 135.1000 ;
	    RECT 55.8000 135.1000 56.2000 135.2000 ;
	    RECT 57.4000 135.1000 57.8000 135.2000 ;
	    RECT 55.8000 134.8000 57.8000 135.1000 ;
	    RECT 70.2000 135.1000 70.6000 135.2000 ;
	    RECT 76.6000 135.1000 77.0000 135.2000 ;
	    RECT 70.2000 134.8000 77.0000 135.1000 ;
	    RECT 83.8000 135.1000 84.2000 135.2000 ;
	    RECT 88.6000 135.1000 89.0000 135.2000 ;
	    RECT 95.8000 135.1000 96.2000 135.2000 ;
	    RECT 83.8000 134.8000 89.0000 135.1000 ;
	    RECT 94.2000 134.8000 96.2000 135.1000 ;
	    RECT 97.4000 135.1000 97.7000 135.8000 ;
	    RECT 171.8000 135.2000 172.1000 135.8000 ;
	    RECT 109.4000 135.1000 109.8000 135.2000 ;
	    RECT 97.4000 134.8000 109.8000 135.1000 ;
	    RECT 114.2000 135.1000 114.6000 135.2000 ;
	    RECT 115.0000 135.1000 115.4000 135.2000 ;
	    RECT 114.2000 134.8000 115.4000 135.1000 ;
	    RECT 115.8000 135.1000 116.2000 135.2000 ;
	    RECT 116.6000 135.1000 117.0000 135.2000 ;
	    RECT 115.8000 134.8000 117.0000 135.1000 ;
	    RECT 120.6000 135.1000 121.0000 135.2000 ;
	    RECT 124.6000 135.1000 125.0000 135.2000 ;
	    RECT 120.6000 134.8000 125.0000 135.1000 ;
	    RECT 133.4000 135.1000 133.8000 135.2000 ;
	    RECT 143.8000 135.1000 144.2000 135.2000 ;
	    RECT 164.6000 135.1000 165.0000 135.2000 ;
	    RECT 166.2000 135.1000 166.6000 135.2000 ;
	    RECT 133.4000 134.8000 166.6000 135.1000 ;
	    RECT 171.8000 134.8000 172.2000 135.2000 ;
	    RECT 18.2000 134.2000 18.5000 134.8000 ;
	    RECT 94.2000 134.2000 94.5000 134.8000 ;
	    RECT 9.4000 134.1000 9.8000 134.2000 ;
	    RECT 7.8000 133.8000 9.8000 134.1000 ;
	    RECT 18.2000 133.8000 18.6000 134.2000 ;
	    RECT 52.6000 134.1000 53.0000 134.2000 ;
	    RECT 55.0000 134.1000 55.4000 134.2000 ;
	    RECT 56.6000 134.1000 57.0000 134.2000 ;
	    RECT 77.4000 134.1000 77.8000 134.2000 ;
	    RECT 52.6000 133.8000 57.0000 134.1000 ;
	    RECT 75.0000 133.8000 77.8000 134.1000 ;
	    RECT 84.6000 134.1000 85.0000 134.2000 ;
	    RECT 90.2000 134.1000 90.6000 134.2000 ;
	    RECT 91.8000 134.1000 92.2000 134.2000 ;
	    RECT 84.6000 133.8000 92.2000 134.1000 ;
	    RECT 94.2000 133.8000 94.6000 134.2000 ;
	    RECT 97.4000 134.1000 97.8000 134.2000 ;
	    RECT 102.2000 134.1000 102.6000 134.2000 ;
	    RECT 97.4000 133.8000 102.6000 134.1000 ;
	    RECT 103.0000 134.1000 103.4000 134.2000 ;
	    RECT 108.6000 134.1000 109.0000 134.2000 ;
	    RECT 103.0000 133.8000 109.0000 134.1000 ;
	    RECT 111.0000 134.1000 111.4000 134.2000 ;
	    RECT 130.2000 134.1000 130.6000 134.2000 ;
	    RECT 111.0000 133.8000 130.6000 134.1000 ;
	    RECT 133.4000 133.8000 133.8000 134.2000 ;
	    RECT 137.4000 134.1000 137.8000 134.2000 ;
	    RECT 140.6000 134.1000 141.0000 134.2000 ;
	    RECT 143.8000 134.1000 144.2000 134.2000 ;
	    RECT 137.4000 133.8000 144.2000 134.1000 ;
	    RECT 151.0000 134.1000 151.4000 134.2000 ;
	    RECT 155.8000 134.1000 156.2000 134.4000 ;
	    RECT 151.0000 134.0000 156.2000 134.1000 ;
	    RECT 158.2000 134.1000 158.6000 134.2000 ;
	    RECT 159.8000 134.1000 160.2000 134.2000 ;
	    RECT 151.0000 133.8000 156.1000 134.0000 ;
	    RECT 158.2000 133.8000 160.2000 134.1000 ;
	    RECT 161.4000 134.1000 161.8000 134.2000 ;
	    RECT 162.2000 134.1000 162.6000 134.2000 ;
	    RECT 165.4000 134.1000 165.8000 134.2000 ;
	    RECT 161.4000 133.8000 165.8000 134.1000 ;
	    RECT 167.0000 133.8000 167.4000 134.2000 ;
	    RECT 7.8000 133.2000 8.1000 133.8000 ;
	    RECT 75.0000 133.2000 75.3000 133.8000 ;
	    RECT 133.4000 133.2000 133.7000 133.8000 ;
	    RECT 167.0000 133.2000 167.3000 133.8000 ;
	    RECT 7.8000 132.8000 8.2000 133.2000 ;
	    RECT 56.6000 133.1000 57.0000 133.2000 ;
	    RECT 63.8000 133.1000 64.2000 133.2000 ;
	    RECT 70.2000 133.1000 70.6000 133.2000 ;
	    RECT 56.6000 132.8000 70.6000 133.1000 ;
	    RECT 75.0000 132.8000 75.4000 133.2000 ;
	    RECT 81.4000 132.8000 81.8000 133.2000 ;
	    RECT 87.8000 133.1000 88.2000 133.2000 ;
	    RECT 99.0000 133.1000 99.4000 133.2000 ;
	    RECT 87.8000 132.8000 99.4000 133.1000 ;
	    RECT 107.8000 133.1000 108.2000 133.2000 ;
	    RECT 115.8000 133.1000 116.2000 133.2000 ;
	    RECT 117.4000 133.1000 117.8000 133.2000 ;
	    RECT 107.8000 132.8000 117.8000 133.1000 ;
	    RECT 118.2000 133.1000 118.6000 133.2000 ;
	    RECT 121.4000 133.1000 121.8000 133.2000 ;
	    RECT 118.2000 132.8000 121.8000 133.1000 ;
	    RECT 122.2000 133.1000 122.6000 133.2000 ;
	    RECT 131.0000 133.1000 131.4000 133.2000 ;
	    RECT 122.2000 132.8000 131.4000 133.1000 ;
	    RECT 133.4000 132.8000 133.8000 133.2000 ;
	    RECT 146.2000 133.1000 146.6000 133.2000 ;
	    RECT 155.8000 133.1000 156.2000 133.2000 ;
	    RECT 146.2000 132.8000 156.2000 133.1000 ;
	    RECT 167.0000 132.8000 167.4000 133.2000 ;
	    RECT 25.4000 132.1000 25.8000 132.2000 ;
	    RECT 32.6000 132.1000 33.0000 132.2000 ;
	    RECT 39.0000 132.1000 39.4000 132.2000 ;
	    RECT 40.6000 132.1000 41.0000 132.2000 ;
	    RECT 43.0000 132.1000 43.4000 132.2000 ;
	    RECT 25.4000 131.8000 43.4000 132.1000 ;
	    RECT 81.4000 132.1000 81.7000 132.8000 ;
	    RECT 98.2000 132.1000 98.6000 132.2000 ;
	    RECT 116.6000 132.1000 117.0000 132.2000 ;
	    RECT 119.8000 132.1000 120.2000 132.2000 ;
	    RECT 127.0000 132.1000 127.4000 132.2000 ;
	    RECT 134.2000 132.1000 134.6000 132.2000 ;
	    RECT 81.4000 131.8000 127.4000 132.1000 ;
	    RECT 129.4000 131.8000 134.6000 132.1000 ;
	    RECT 142.2000 132.1000 142.6000 132.2000 ;
	    RECT 156.6000 132.1000 157.0000 132.2000 ;
	    RECT 161.4000 132.1000 161.8000 132.2000 ;
	    RECT 142.2000 131.8000 161.8000 132.1000 ;
	    RECT 165.4000 132.1000 165.8000 132.2000 ;
	    RECT 166.2000 132.1000 166.6000 132.2000 ;
	    RECT 165.4000 131.8000 166.6000 132.1000 ;
	    RECT 129.4000 131.2000 129.7000 131.8000 ;
	    RECT 77.4000 131.1000 77.8000 131.2000 ;
	    RECT 78.2000 131.1000 78.6000 131.2000 ;
	    RECT 81.4000 131.1000 81.8000 131.2000 ;
	    RECT 77.4000 130.8000 81.8000 131.1000 ;
	    RECT 115.8000 130.8000 116.2000 131.2000 ;
	    RECT 124.6000 131.1000 125.0000 131.2000 ;
	    RECT 129.4000 131.1000 129.8000 131.2000 ;
	    RECT 124.6000 130.8000 129.8000 131.1000 ;
	    RECT 131.0000 131.1000 131.4000 131.2000 ;
	    RECT 147.0000 131.1000 147.4000 131.2000 ;
	    RECT 163.0000 131.1000 163.4000 131.2000 ;
	    RECT 131.0000 130.8000 163.4000 131.1000 ;
	    RECT 115.8000 130.2000 116.1000 130.8000 ;
	    RECT 1.4000 130.1000 1.8000 130.2000 ;
	    RECT 8.6000 130.1000 9.0000 130.2000 ;
	    RECT 1.4000 129.8000 9.0000 130.1000 ;
	    RECT 103.8000 130.1000 104.2000 130.2000 ;
	    RECT 104.6000 130.1000 105.0000 130.2000 ;
	    RECT 103.8000 129.8000 105.0000 130.1000 ;
	    RECT 115.8000 129.8000 116.2000 130.2000 ;
	    RECT 123.8000 130.1000 124.2000 130.2000 ;
	    RECT 127.8000 130.1000 128.2000 130.2000 ;
	    RECT 143.0000 130.1000 143.4000 130.2000 ;
	    RECT 145.4000 130.1000 145.8000 130.2000 ;
	    RECT 149.4000 130.1000 149.8000 130.2000 ;
	    RECT 154.2000 130.1000 154.6000 130.2000 ;
	    RECT 157.4000 130.1000 157.8000 130.2000 ;
	    RECT 159.0000 130.1000 159.4000 130.2000 ;
	    RECT 123.8000 129.8000 159.4000 130.1000 ;
	    RECT 101.4000 129.1000 101.8000 129.2000 ;
	    RECT 101.4000 128.8000 104.1000 129.1000 ;
	    RECT 103.8000 128.2000 104.1000 128.8000 ;
	    RECT 118.2000 128.8000 118.6000 129.2000 ;
	    RECT 130.2000 129.1000 130.6000 129.2000 ;
	    RECT 129.4000 128.8000 130.6000 129.1000 ;
	    RECT 138.2000 129.1000 138.6000 129.2000 ;
	    RECT 141.4000 129.1000 141.8000 129.2000 ;
	    RECT 155.0000 129.1000 155.4000 129.2000 ;
	    RECT 138.2000 128.8000 155.4000 129.1000 ;
	    RECT 155.8000 129.1000 156.2000 129.2000 ;
	    RECT 158.2000 129.1000 158.6000 129.2000 ;
	    RECT 167.0000 129.1000 167.4000 129.2000 ;
	    RECT 155.8000 128.8000 167.4000 129.1000 ;
	    RECT 10.2000 128.1000 10.6000 128.2000 ;
	    RECT 22.2000 128.1000 22.6000 128.2000 ;
	    RECT 10.2000 127.8000 22.6000 128.1000 ;
	    RECT 66.2000 127.8000 66.6000 128.2000 ;
	    RECT 68.6000 128.1000 69.0000 128.2000 ;
	    RECT 69.4000 128.1000 69.8000 128.2000 ;
	    RECT 68.6000 127.8000 69.8000 128.1000 ;
	    RECT 70.2000 128.1000 70.6000 128.2000 ;
	    RECT 73.4000 128.1000 73.8000 128.2000 ;
	    RECT 70.2000 127.8000 73.8000 128.1000 ;
	    RECT 95.8000 128.1000 96.2000 128.2000 ;
	    RECT 98.2000 128.1000 98.6000 128.2000 ;
	    RECT 95.8000 127.8000 98.6000 128.1000 ;
	    RECT 100.6000 127.8000 101.0000 128.2000 ;
	    RECT 103.8000 127.8000 104.2000 128.2000 ;
	    RECT 111.8000 127.8000 112.2000 128.2000 ;
	    RECT 112.6000 128.1000 113.0000 128.2000 ;
	    RECT 118.2000 128.1000 118.5000 128.8000 ;
	    RECT 129.4000 128.2000 129.7000 128.8000 ;
	    RECT 127.8000 128.1000 128.2000 128.2000 ;
	    RECT 112.6000 127.8000 128.2000 128.1000 ;
	    RECT 129.4000 127.8000 129.8000 128.2000 ;
	    RECT 131.8000 128.1000 132.2000 128.2000 ;
	    RECT 135.8000 128.1000 136.2000 128.2000 ;
	    RECT 136.6000 128.1000 137.0000 128.2000 ;
	    RECT 131.8000 127.8000 137.0000 128.1000 ;
	    RECT 142.2000 128.1000 142.6000 128.2000 ;
	    RECT 144.6000 128.1000 145.0000 128.2000 ;
	    RECT 148.6000 128.1000 149.0000 128.2000 ;
	    RECT 142.2000 127.8000 149.0000 128.1000 ;
	    RECT 155.0000 128.1000 155.4000 128.2000 ;
	    RECT 161.4000 128.1000 161.8000 128.2000 ;
	    RECT 155.0000 127.8000 161.8000 128.1000 ;
	    RECT 21.4000 126.8000 21.8000 127.2000 ;
	    RECT 27.0000 126.8000 27.4000 127.2000 ;
	    RECT 27.8000 127.1000 28.2000 127.2000 ;
	    RECT 28.6000 127.1000 29.0000 127.2000 ;
	    RECT 27.8000 126.8000 29.0000 127.1000 ;
	    RECT 29.4000 127.1000 29.8000 127.2000 ;
	    RECT 32.6000 127.1000 33.0000 127.2000 ;
	    RECT 29.4000 126.8000 33.0000 127.1000 ;
	    RECT 46.2000 126.8000 46.6000 127.2000 ;
	    RECT 52.6000 126.8000 53.0000 127.2000 ;
	    RECT 66.2000 127.1000 66.5000 127.8000 ;
	    RECT 71.0000 127.1000 71.4000 127.2000 ;
	    RECT 66.2000 126.8000 71.4000 127.1000 ;
	    RECT 100.6000 127.1000 100.9000 127.8000 ;
	    RECT 104.6000 127.1000 105.0000 127.2000 ;
	    RECT 100.6000 126.8000 105.0000 127.1000 ;
	    RECT 110.2000 127.1000 110.6000 127.2000 ;
	    RECT 111.0000 127.1000 111.4000 127.2000 ;
	    RECT 110.2000 126.8000 111.4000 127.1000 ;
	    RECT 111.8000 127.1000 112.1000 127.8000 ;
	    RECT 166.2000 127.1000 166.6000 127.2000 ;
	    RECT 111.8000 126.8000 166.6000 127.1000 ;
	    RECT 167.0000 126.8000 167.4000 127.2000 ;
	    RECT 17.4000 126.1000 17.8000 126.2000 ;
	    RECT 21.4000 126.1000 21.7000 126.8000 ;
	    RECT 17.4000 125.8000 21.7000 126.1000 ;
	    RECT 27.0000 126.1000 27.3000 126.8000 ;
	    RECT 28.6000 126.1000 29.0000 126.2000 ;
	    RECT 27.0000 125.8000 29.0000 126.1000 ;
	    RECT 46.2000 126.1000 46.5000 126.8000 ;
	    RECT 47.8000 126.1000 48.2000 126.2000 ;
	    RECT 46.2000 125.8000 48.2000 126.1000 ;
	    RECT 52.6000 126.1000 52.9000 126.8000 ;
	    RECT 54.2000 126.1000 54.6000 126.2000 ;
	    RECT 52.6000 125.8000 54.6000 126.1000 ;
	    RECT 63.0000 126.1000 63.4000 126.2000 ;
	    RECT 66.2000 126.1000 66.6000 126.2000 ;
	    RECT 63.0000 125.8000 66.6000 126.1000 ;
	    RECT 68.6000 126.1000 69.0000 126.2000 ;
	    RECT 73.4000 126.1000 73.8000 126.2000 ;
	    RECT 68.6000 125.8000 73.8000 126.1000 ;
	    RECT 91.0000 126.1000 91.4000 126.3000 ;
	    RECT 91.8000 126.1000 92.2000 126.2000 ;
	    RECT 91.0000 125.8000 92.2000 126.1000 ;
	    RECT 99.0000 126.1000 99.4000 126.2000 ;
	    RECT 112.6000 126.1000 113.0000 126.2000 ;
	    RECT 99.0000 125.8000 113.0000 126.1000 ;
	    RECT 113.4000 126.1000 113.8000 126.2000 ;
	    RECT 119.8000 126.1000 120.2000 126.2000 ;
	    RECT 121.4000 126.1000 121.8000 126.2000 ;
	    RECT 122.2000 126.1000 122.6000 126.2000 ;
	    RECT 113.4000 125.8000 120.2000 126.1000 ;
	    RECT 120.6000 125.8000 122.6000 126.1000 ;
	    RECT 126.2000 126.1000 126.6000 126.2000 ;
	    RECT 131.0000 126.1000 131.4000 126.2000 ;
	    RECT 126.2000 125.8000 131.4000 126.1000 ;
	    RECT 135.0000 126.1000 135.4000 126.2000 ;
	    RECT 135.8000 126.1000 136.2000 126.2000 ;
	    RECT 135.0000 125.8000 136.2000 126.1000 ;
	    RECT 153.4000 126.1000 153.8000 126.2000 ;
	    RECT 155.8000 126.1000 156.2000 126.2000 ;
	    RECT 153.4000 125.8000 156.2000 126.1000 ;
	    RECT 160.6000 126.1000 161.0000 126.2000 ;
	    RECT 162.2000 126.1000 162.6000 126.2000 ;
	    RECT 160.6000 125.8000 162.6000 126.1000 ;
	    RECT 166.2000 126.1000 166.6000 126.2000 ;
	    RECT 167.0000 126.1000 167.3000 126.8000 ;
	    RECT 166.2000 125.8000 167.3000 126.1000 ;
	    RECT 38.2000 125.1000 38.6000 125.2000 ;
	    RECT 39.0000 125.1000 39.4000 125.2000 ;
	    RECT 38.2000 124.8000 39.4000 125.1000 ;
	    RECT 50.2000 125.1000 50.6000 125.2000 ;
	    RECT 56.6000 125.1000 57.0000 125.2000 ;
	    RECT 67.8000 125.1000 68.2000 125.2000 ;
	    RECT 72.6000 125.1000 73.0000 125.2000 ;
	    RECT 50.2000 124.8000 73.0000 125.1000 ;
	    RECT 83.8000 125.1000 84.2000 125.2000 ;
	    RECT 86.2000 125.1000 86.6000 125.2000 ;
	    RECT 95.8000 125.1000 96.2000 125.2000 ;
	    RECT 83.8000 124.8000 96.2000 125.1000 ;
	    RECT 98.2000 125.1000 98.6000 125.2000 ;
	    RECT 102.2000 125.1000 102.6000 125.2000 ;
	    RECT 98.2000 124.8000 102.6000 125.1000 ;
	    RECT 103.8000 125.1000 104.2000 125.2000 ;
	    RECT 121.4000 125.1000 121.8000 125.2000 ;
	    RECT 123.8000 125.1000 124.2000 125.2000 ;
	    RECT 103.8000 124.8000 124.2000 125.1000 ;
	    RECT 160.6000 125.1000 161.0000 125.2000 ;
	    RECT 161.4000 125.1000 161.8000 125.2000 ;
	    RECT 160.6000 124.8000 161.8000 125.1000 ;
	    RECT 71.0000 124.2000 71.3000 124.8000 ;
	    RECT 16.6000 124.1000 17.0000 124.2000 ;
	    RECT 19.8000 124.1000 20.2000 124.2000 ;
	    RECT 16.6000 123.8000 20.2000 124.1000 ;
	    RECT 28.6000 124.1000 29.0000 124.2000 ;
	    RECT 29.4000 124.1000 29.8000 124.2000 ;
	    RECT 38.2000 124.1000 38.6000 124.2000 ;
	    RECT 28.6000 123.8000 29.8000 124.1000 ;
	    RECT 35.8000 123.8000 38.6000 124.1000 ;
	    RECT 43.0000 124.1000 43.4000 124.2000 ;
	    RECT 47.0000 124.1000 47.4000 124.2000 ;
	    RECT 43.0000 123.8000 47.4000 124.1000 ;
	    RECT 59.0000 124.1000 59.4000 124.2000 ;
	    RECT 60.6000 124.1000 61.0000 124.2000 ;
	    RECT 59.0000 123.8000 61.0000 124.1000 ;
	    RECT 71.0000 123.8000 71.4000 124.2000 ;
	    RECT 98.2000 124.1000 98.6000 124.2000 ;
	    RECT 115.0000 124.1000 115.4000 124.2000 ;
	    RECT 98.2000 123.8000 115.4000 124.1000 ;
	    RECT 120.6000 124.1000 121.0000 124.2000 ;
	    RECT 156.6000 124.1000 157.0000 124.2000 ;
	    RECT 161.4000 124.1000 161.8000 124.2000 ;
	    RECT 120.6000 123.8000 161.8000 124.1000 ;
	    RECT 35.8000 123.2000 36.1000 123.8000 ;
	    RECT 35.8000 122.8000 36.2000 123.2000 ;
	    RECT 55.0000 123.1000 55.4000 123.2000 ;
	    RECT 62.2000 123.1000 62.6000 123.2000 ;
	    RECT 55.0000 122.8000 62.6000 123.1000 ;
	    RECT 71.8000 123.1000 72.2000 123.2000 ;
	    RECT 104.6000 123.1000 105.0000 123.2000 ;
	    RECT 126.2000 123.1000 126.6000 123.2000 ;
	    RECT 71.8000 122.8000 126.6000 123.1000 ;
	    RECT 134.2000 123.1000 134.6000 123.2000 ;
	    RECT 139.8000 123.1000 140.2000 123.2000 ;
	    RECT 144.6000 123.1000 145.0000 123.2000 ;
	    RECT 134.2000 122.8000 145.0000 123.1000 ;
	    RECT 2.2000 122.1000 2.6000 122.2000 ;
	    RECT 1.4000 121.8000 2.6000 122.1000 ;
	    RECT 13.4000 122.1000 13.8000 122.2000 ;
	    RECT 17.4000 122.1000 17.8000 122.2000 ;
	    RECT 26.2000 122.1000 26.6000 122.2000 ;
	    RECT 30.2000 122.1000 30.6000 122.2000 ;
	    RECT 34.2000 122.1000 34.6000 122.2000 ;
	    RECT 13.4000 121.8000 34.6000 122.1000 ;
	    RECT 114.2000 122.1000 114.6000 122.2000 ;
	    RECT 122.2000 122.1000 122.6000 122.2000 ;
	    RECT 114.2000 121.8000 122.6000 122.1000 ;
	    RECT 124.6000 122.1000 125.0000 122.2000 ;
	    RECT 128.6000 122.1000 129.0000 122.2000 ;
	    RECT 137.4000 122.1000 137.8000 122.2000 ;
	    RECT 124.6000 121.8000 137.8000 122.1000 ;
	    RECT 1.4000 121.2000 1.7000 121.8000 ;
	    RECT 1.4000 120.8000 1.8000 121.2000 ;
	    RECT 31.8000 121.1000 32.2000 121.2000 ;
	    RECT 41.4000 121.1000 41.8000 121.2000 ;
	    RECT 31.8000 120.8000 41.8000 121.1000 ;
	    RECT 19.8000 119.1000 20.2000 119.2000 ;
	    RECT 32.6000 119.1000 33.0000 119.2000 ;
	    RECT 19.8000 118.8000 33.0000 119.1000 ;
	    RECT 52.6000 118.8000 53.0000 119.2000 ;
	    RECT 91.8000 119.1000 92.2000 119.2000 ;
	    RECT 95.0000 119.1000 95.4000 119.2000 ;
	    RECT 91.8000 118.8000 95.4000 119.1000 ;
	    RECT 11.0000 118.1000 11.4000 118.2000 ;
	    RECT 21.4000 118.1000 21.8000 118.2000 ;
	    RECT 11.0000 117.8000 21.8000 118.1000 ;
	    RECT 52.6000 118.1000 52.9000 118.8000 ;
	    RECT 57.4000 118.1000 57.8000 118.2000 ;
	    RECT 52.6000 117.8000 57.8000 118.1000 ;
	    RECT 69.4000 117.8000 69.8000 118.2000 ;
	    RECT 69.4000 117.2000 69.7000 117.8000 ;
	    RECT 11.0000 117.1000 11.4000 117.2000 ;
	    RECT 11.8000 117.1000 12.2000 117.2000 ;
	    RECT 11.0000 116.8000 12.2000 117.1000 ;
	    RECT 30.2000 117.1000 30.6000 117.2000 ;
	    RECT 31.8000 117.1000 32.2000 117.2000 ;
	    RECT 30.2000 116.8000 32.2000 117.1000 ;
	    RECT 33.4000 117.1000 33.8000 117.2000 ;
	    RECT 37.4000 117.1000 37.8000 117.2000 ;
	    RECT 33.4000 116.8000 37.8000 117.1000 ;
	    RECT 39.0000 117.1000 39.4000 117.2000 ;
	    RECT 45.4000 117.1000 45.8000 117.2000 ;
	    RECT 39.0000 116.8000 45.8000 117.1000 ;
	    RECT 48.6000 117.1000 49.0000 117.2000 ;
	    RECT 68.6000 117.1000 69.0000 117.2000 ;
	    RECT 48.6000 116.8000 69.0000 117.1000 ;
	    RECT 69.4000 116.8000 69.8000 117.2000 ;
	    RECT 147.0000 116.8000 147.4000 117.2000 ;
	    RECT 149.4000 117.1000 149.8000 117.2000 ;
	    RECT 151.8000 117.1000 152.2000 117.2000 ;
	    RECT 152.6000 117.1000 153.0000 117.2000 ;
	    RECT 149.4000 116.8000 153.0000 117.1000 ;
	    RECT 158.2000 116.8000 158.6000 117.2000 ;
	    RECT 7.0000 116.1000 7.4000 116.2000 ;
	    RECT 12.6000 116.1000 13.0000 116.2000 ;
	    RECT 7.0000 115.8000 13.0000 116.1000 ;
	    RECT 14.2000 116.1000 14.6000 116.2000 ;
	    RECT 15.8000 116.1000 16.2000 116.2000 ;
	    RECT 14.2000 115.8000 16.2000 116.1000 ;
	    RECT 47.8000 116.1000 48.2000 116.2000 ;
	    RECT 48.6000 116.1000 49.0000 116.2000 ;
	    RECT 47.8000 115.8000 49.0000 116.1000 ;
	    RECT 87.0000 115.8000 87.4000 116.2000 ;
	    RECT 123.8000 116.1000 124.2000 116.2000 ;
	    RECT 127.8000 116.1000 128.2000 116.2000 ;
	    RECT 130.2000 116.1000 130.6000 116.2000 ;
	    RECT 135.8000 116.1000 136.2000 116.2000 ;
	    RECT 123.8000 115.8000 136.2000 116.1000 ;
	    RECT 139.0000 116.1000 139.4000 116.2000 ;
	    RECT 147.0000 116.1000 147.3000 116.8000 ;
	    RECT 139.0000 115.8000 147.3000 116.1000 ;
	    RECT 151.8000 116.1000 152.2000 116.2000 ;
	    RECT 158.2000 116.1000 158.5000 116.8000 ;
	    RECT 151.8000 115.8000 158.5000 116.1000 ;
	    RECT 160.6000 115.8000 161.0000 116.2000 ;
	    RECT 32.6000 115.1000 33.0000 115.2000 ;
	    RECT 38.2000 115.1000 38.6000 115.2000 ;
	    RECT 32.6000 114.8000 38.6000 115.1000 ;
	    RECT 78.2000 114.8000 78.6000 115.2000 ;
	    RECT 83.8000 114.8000 84.2000 115.2000 ;
	    RECT 87.0000 115.1000 87.3000 115.8000 ;
	    RECT 92.6000 115.1000 93.0000 115.2000 ;
	    RECT 87.0000 114.8000 93.0000 115.1000 ;
	    RECT 116.6000 115.1000 117.0000 115.2000 ;
	    RECT 120.6000 115.1000 121.0000 115.2000 ;
	    RECT 116.6000 114.8000 121.0000 115.1000 ;
	    RECT 129.4000 115.1000 129.8000 115.2000 ;
	    RECT 132.6000 115.1000 133.0000 115.2000 ;
	    RECT 129.4000 114.8000 133.0000 115.1000 ;
	    RECT 135.8000 115.1000 136.2000 115.2000 ;
	    RECT 140.6000 115.1000 141.0000 115.2000 ;
	    RECT 135.8000 114.8000 141.0000 115.1000 ;
	    RECT 147.8000 115.1000 148.2000 115.2000 ;
	    RECT 160.6000 115.1000 160.9000 115.8000 ;
	    RECT 147.8000 114.8000 160.9000 115.1000 ;
	    RECT 167.8000 115.1000 168.2000 115.2000 ;
	    RECT 171.8000 115.1000 172.2000 115.2000 ;
	    RECT 167.8000 114.8000 172.2000 115.1000 ;
	    RECT 78.2000 114.2000 78.5000 114.8000 ;
	    RECT 83.8000 114.2000 84.1000 114.8000 ;
	    RECT 47.0000 114.1000 47.4000 114.2000 ;
	    RECT 56.6000 114.1000 57.0000 114.2000 ;
	    RECT 44.6000 113.8000 47.4000 114.1000 ;
	    RECT 51.0000 113.8000 57.0000 114.1000 ;
	    RECT 78.2000 113.8000 78.6000 114.2000 ;
	    RECT 83.8000 113.8000 84.2000 114.2000 ;
	    RECT 139.8000 114.1000 140.2000 114.2000 ;
	    RECT 151.8000 114.1000 152.2000 114.2000 ;
	    RECT 154.2000 114.1000 154.6000 114.2000 ;
	    RECT 156.6000 114.1000 157.0000 114.2000 ;
	    RECT 159.8000 114.1000 160.2000 114.2000 ;
	    RECT 139.8000 113.8000 144.9000 114.1000 ;
	    RECT 151.8000 113.8000 160.2000 114.1000 ;
	    RECT 160.6000 114.1000 161.0000 114.2000 ;
	    RECT 161.4000 114.1000 161.8000 114.2000 ;
	    RECT 160.6000 113.8000 161.8000 114.1000 ;
	    RECT 44.6000 113.2000 44.9000 113.8000 ;
	    RECT 51.0000 113.2000 51.3000 113.8000 ;
	    RECT 144.6000 113.2000 144.9000 113.8000 ;
	    RECT 1.4000 113.1000 1.8000 113.2000 ;
	    RECT 2.2000 113.1000 2.6000 113.2000 ;
	    RECT 3.8000 113.1000 4.2000 113.2000 ;
	    RECT 1.4000 112.8000 4.2000 113.1000 ;
	    RECT 44.6000 112.8000 45.0000 113.2000 ;
	    RECT 51.0000 112.8000 51.4000 113.2000 ;
	    RECT 51.8000 113.1000 52.2000 113.2000 ;
	    RECT 59.0000 113.1000 59.4000 113.2000 ;
	    RECT 51.8000 112.8000 59.4000 113.1000 ;
	    RECT 140.6000 113.1000 141.0000 113.2000 ;
	    RECT 142.2000 113.1000 142.6000 113.2000 ;
	    RECT 140.6000 112.8000 142.6000 113.1000 ;
	    RECT 144.6000 112.8000 145.0000 113.2000 ;
	    RECT 150.2000 113.1000 150.6000 113.2000 ;
	    RECT 152.6000 113.1000 153.0000 113.2000 ;
	    RECT 155.0000 113.1000 155.4000 113.2000 ;
	    RECT 157.4000 113.1000 157.8000 113.2000 ;
	    RECT 150.2000 112.8000 157.8000 113.1000 ;
	    RECT 11.0000 112.1000 11.4000 112.2000 ;
	    RECT 13.4000 112.1000 13.8000 112.2000 ;
	    RECT 17.4000 112.1000 17.8000 112.2000 ;
	    RECT 19.8000 112.1000 20.2000 112.2000 ;
	    RECT 23.8000 112.1000 24.2000 112.2000 ;
	    RECT 31.0000 112.1000 31.4000 112.2000 ;
	    RECT 11.0000 111.8000 31.4000 112.1000 ;
	    RECT 39.0000 112.1000 39.4000 112.2000 ;
	    RECT 41.4000 112.1000 41.8000 112.2000 ;
	    RECT 48.6000 112.1000 49.0000 112.2000 ;
	    RECT 51.8000 112.1000 52.2000 112.2000 ;
	    RECT 39.0000 111.8000 52.2000 112.1000 ;
	    RECT 79.8000 112.1000 80.2000 112.2000 ;
	    RECT 90.2000 112.1000 90.6000 112.2000 ;
	    RECT 79.8000 111.8000 90.6000 112.1000 ;
	    RECT 123.8000 112.1000 124.2000 112.2000 ;
	    RECT 127.0000 112.1000 127.4000 112.2000 ;
	    RECT 131.8000 112.1000 132.2000 112.2000 ;
	    RECT 138.2000 112.1000 138.6000 112.2000 ;
	    RECT 142.2000 112.1000 142.6000 112.2000 ;
	    RECT 146.2000 112.1000 146.6000 112.2000 ;
	    RECT 123.8000 111.8000 146.6000 112.1000 ;
	    RECT 67.0000 111.1000 67.4000 111.2000 ;
	    RECT 96.6000 111.1000 97.0000 111.2000 ;
	    RECT 67.0000 110.8000 97.0000 111.1000 ;
	    RECT 97.4000 111.1000 97.8000 111.2000 ;
	    RECT 103.0000 111.1000 103.4000 111.2000 ;
	    RECT 97.4000 110.8000 103.4000 111.1000 ;
	    RECT 169.4000 111.1000 169.8000 111.2000 ;
	    RECT 171.0000 111.1000 171.4000 111.2000 ;
	    RECT 169.4000 110.8000 171.4000 111.1000 ;
	    RECT 47.0000 110.1000 47.4000 110.2000 ;
	    RECT 64.6000 110.1000 65.0000 110.2000 ;
	    RECT 75.8000 110.1000 76.2000 110.2000 ;
	    RECT 47.0000 109.8000 64.1000 110.1000 ;
	    RECT 64.6000 109.8000 76.2000 110.1000 ;
	    RECT 80.6000 110.1000 81.0000 110.2000 ;
	    RECT 81.4000 110.1000 81.8000 110.2000 ;
	    RECT 80.6000 109.8000 81.8000 110.1000 ;
	    RECT 63.8000 109.1000 64.1000 109.8000 ;
	    RECT 67.0000 109.1000 67.4000 109.2000 ;
	    RECT 63.8000 108.8000 67.4000 109.1000 ;
	    RECT 70.2000 109.1000 70.6000 109.2000 ;
	    RECT 91.0000 109.1000 91.4000 109.2000 ;
	    RECT 104.6000 109.1000 105.0000 109.2000 ;
	    RECT 70.2000 108.8000 91.4000 109.1000 ;
	    RECT 102.2000 108.8000 105.0000 109.1000 ;
	    RECT 111.8000 109.1000 112.2000 109.2000 ;
	    RECT 117.4000 109.1000 117.8000 109.2000 ;
	    RECT 111.8000 108.8000 117.8000 109.1000 ;
	    RECT 141.4000 108.8000 141.8000 109.2000 ;
	    RECT 102.2000 108.2000 102.5000 108.8000 ;
	    RECT 22.2000 107.8000 22.6000 108.2000 ;
	    RECT 62.2000 108.1000 62.6000 108.2000 ;
	    RECT 92.6000 108.1000 93.0000 108.2000 ;
	    RECT 62.2000 107.8000 93.0000 108.1000 ;
	    RECT 102.2000 107.8000 102.6000 108.2000 ;
	    RECT 127.8000 108.1000 128.2000 108.2000 ;
	    RECT 130.2000 108.1000 130.6000 108.2000 ;
	    RECT 127.8000 107.8000 130.6000 108.1000 ;
	    RECT 138.2000 108.1000 138.6000 108.2000 ;
	    RECT 141.4000 108.1000 141.7000 108.8000 ;
	    RECT 138.2000 107.8000 141.7000 108.1000 ;
	    RECT 9.4000 106.8000 9.8000 107.2000 ;
	    RECT 11.0000 106.8000 11.4000 107.2000 ;
	    RECT 15.8000 107.1000 16.2000 107.2000 ;
	    RECT 19.8000 107.1000 20.2000 107.2000 ;
	    RECT 15.8000 106.8000 20.2000 107.1000 ;
	    RECT 22.2000 107.1000 22.5000 107.8000 ;
	    RECT 24.6000 107.1000 25.0000 107.2000 ;
	    RECT 22.2000 106.8000 25.0000 107.1000 ;
	    RECT 43.8000 106.8000 44.2000 107.2000 ;
	    RECT 54.2000 106.8000 54.6000 107.2000 ;
	    RECT 57.4000 107.1000 57.8000 107.2000 ;
	    RECT 62.2000 107.1000 62.6000 107.2000 ;
	    RECT 57.4000 106.8000 62.6000 107.1000 ;
	    RECT 81.4000 107.1000 81.8000 107.2000 ;
	    RECT 82.2000 107.1000 82.6000 107.2000 ;
	    RECT 81.4000 106.8000 82.6000 107.1000 ;
	    RECT 89.4000 106.8000 89.8000 107.2000 ;
	    RECT 107.0000 107.1000 107.4000 107.2000 ;
	    RECT 123.0000 107.1000 123.4000 107.2000 ;
	    RECT 107.0000 106.8000 123.4000 107.1000 ;
	    RECT 136.6000 107.1000 137.0000 107.2000 ;
	    RECT 139.0000 107.1000 139.4000 107.2000 ;
	    RECT 139.8000 107.1000 140.2000 107.2000 ;
	    RECT 136.6000 106.8000 140.2000 107.1000 ;
	    RECT 3.8000 106.1000 4.2000 106.2000 ;
	    RECT 5.4000 106.1000 5.8000 106.2000 ;
	    RECT 3.8000 105.8000 5.8000 106.1000 ;
	    RECT 9.4000 106.1000 9.7000 106.8000 ;
	    RECT 11.0000 106.1000 11.3000 106.8000 ;
	    RECT 9.4000 105.8000 11.3000 106.1000 ;
	    RECT 11.8000 106.1000 12.2000 106.2000 ;
	    RECT 15.0000 106.1000 15.4000 106.2000 ;
	    RECT 11.8000 105.8000 15.4000 106.1000 ;
	    RECT 22.2000 106.1000 22.6000 106.2000 ;
	    RECT 27.8000 106.1000 28.2000 106.2000 ;
	    RECT 22.2000 105.8000 28.2000 106.1000 ;
	    RECT 31.0000 106.1000 31.4000 106.2000 ;
	    RECT 35.8000 106.1000 36.2000 106.2000 ;
	    RECT 31.0000 105.8000 36.2000 106.1000 ;
	    RECT 39.0000 106.1000 39.4000 106.2000 ;
	    RECT 39.8000 106.1000 40.2000 106.2000 ;
	    RECT 39.0000 105.8000 40.2000 106.1000 ;
	    RECT 43.8000 106.1000 44.1000 106.8000 ;
	    RECT 49.4000 106.1000 49.8000 106.2000 ;
	    RECT 43.8000 105.8000 49.8000 106.1000 ;
	    RECT 54.2000 106.1000 54.5000 106.8000 ;
	    RECT 55.0000 106.1000 55.4000 106.2000 ;
	    RECT 54.2000 105.8000 55.4000 106.1000 ;
	    RECT 57.4000 106.1000 57.8000 106.2000 ;
	    RECT 63.0000 106.1000 63.4000 106.2000 ;
	    RECT 57.4000 105.8000 63.4000 106.1000 ;
	    RECT 64.6000 106.1000 65.0000 106.2000 ;
	    RECT 67.8000 106.1000 68.2000 106.2000 ;
	    RECT 64.6000 105.8000 68.2000 106.1000 ;
	    RECT 75.8000 106.1000 76.2000 106.2000 ;
	    RECT 83.8000 106.1000 84.2000 106.2000 ;
	    RECT 87.0000 106.1000 87.4000 106.2000 ;
	    RECT 75.8000 105.8000 87.4000 106.1000 ;
	    RECT 89.4000 106.1000 89.7000 106.8000 ;
	    RECT 91.0000 106.1000 91.4000 106.2000 ;
	    RECT 101.4000 106.1000 101.8000 106.2000 ;
	    RECT 89.4000 105.8000 91.4000 106.1000 ;
	    RECT 99.0000 105.8000 101.8000 106.1000 ;
	    RECT 110.2000 106.1000 110.6000 106.2000 ;
	    RECT 115.0000 106.1000 115.4000 106.2000 ;
	    RECT 110.2000 105.8000 115.4000 106.1000 ;
	    RECT 116.6000 105.8000 117.0000 106.2000 ;
	    RECT 125.4000 106.1000 125.8000 106.2000 ;
	    RECT 127.0000 106.1000 127.4000 106.2000 ;
	    RECT 125.4000 105.8000 127.4000 106.1000 ;
	    RECT 130.2000 106.1000 130.6000 106.2000 ;
	    RECT 132.6000 106.1000 133.0000 106.2000 ;
	    RECT 130.2000 105.8000 133.0000 106.1000 ;
	    RECT 163.8000 106.1000 164.2000 106.2000 ;
	    RECT 163.8000 105.8000 164.9000 106.1000 ;
	    RECT 1.4000 105.1000 1.8000 105.2000 ;
	    RECT 1.4000 104.8000 5.7000 105.1000 ;
	    RECT 5.4000 104.2000 5.7000 104.8000 ;
	    RECT 8.6000 104.8000 9.0000 105.2000 ;
	    RECT 35.8000 104.8000 36.2000 105.2000 ;
	    RECT 37.4000 105.1000 37.8000 105.2000 ;
	    RECT 39.8000 105.1000 40.2000 105.2000 ;
	    RECT 37.4000 104.8000 40.2000 105.1000 ;
	    RECT 63.8000 105.1000 64.2000 105.2000 ;
	    RECT 67.8000 105.1000 68.2000 105.2000 ;
	    RECT 63.8000 104.8000 68.2000 105.1000 ;
	    RECT 68.6000 105.1000 69.0000 105.2000 ;
	    RECT 75.8000 105.1000 76.1000 105.8000 ;
	    RECT 99.0000 105.2000 99.3000 105.8000 ;
	    RECT 116.6000 105.2000 116.9000 105.8000 ;
	    RECT 164.6000 105.2000 164.9000 105.8000 ;
	    RECT 68.6000 104.8000 76.1000 105.1000 ;
	    RECT 80.6000 105.1000 81.0000 105.2000 ;
	    RECT 82.2000 105.1000 82.6000 105.2000 ;
	    RECT 92.6000 105.1000 93.0000 105.2000 ;
	    RECT 80.6000 104.8000 93.0000 105.1000 ;
	    RECT 99.0000 104.8000 99.4000 105.2000 ;
	    RECT 100.6000 105.1000 101.0000 105.2000 ;
	    RECT 107.0000 105.1000 107.4000 105.2000 ;
	    RECT 100.6000 104.8000 107.4000 105.1000 ;
	    RECT 116.6000 104.8000 117.0000 105.2000 ;
	    RECT 119.0000 105.1000 119.4000 105.2000 ;
	    RECT 130.2000 105.1000 130.6000 105.2000 ;
	    RECT 119.0000 104.8000 130.6000 105.1000 ;
	    RECT 137.4000 105.1000 137.8000 105.2000 ;
	    RECT 139.0000 105.1000 139.4000 105.2000 ;
	    RECT 137.4000 104.8000 139.4000 105.1000 ;
	    RECT 164.6000 104.8000 165.0000 105.2000 ;
	    RECT 5.4000 103.8000 5.8000 104.2000 ;
	    RECT 7.0000 104.1000 7.4000 104.2000 ;
	    RECT 8.6000 104.1000 8.9000 104.8000 ;
	    RECT 7.0000 103.8000 8.9000 104.1000 ;
	    RECT 9.4000 104.1000 9.8000 104.2000 ;
	    RECT 14.2000 104.1000 14.6000 104.2000 ;
	    RECT 9.4000 103.8000 14.6000 104.1000 ;
	    RECT 16.6000 104.1000 17.0000 104.2000 ;
	    RECT 26.2000 104.1000 26.6000 104.2000 ;
	    RECT 27.8000 104.1000 28.2000 104.2000 ;
	    RECT 16.6000 103.8000 28.2000 104.1000 ;
	    RECT 32.6000 104.1000 33.0000 104.2000 ;
	    RECT 35.8000 104.1000 36.1000 104.8000 ;
	    RECT 32.6000 103.8000 36.1000 104.1000 ;
	    RECT 47.8000 104.1000 48.2000 104.2000 ;
	    RECT 48.6000 104.1000 49.0000 104.2000 ;
	    RECT 47.8000 103.8000 49.0000 104.1000 ;
	    RECT 57.4000 104.1000 57.8000 104.2000 ;
	    RECT 58.2000 104.1000 58.6000 104.2000 ;
	    RECT 57.4000 103.8000 58.6000 104.1000 ;
	    RECT 76.6000 104.1000 77.0000 104.2000 ;
	    RECT 77.4000 104.1000 77.8000 104.2000 ;
	    RECT 76.6000 103.8000 77.8000 104.1000 ;
	    RECT 84.6000 104.1000 85.0000 104.2000 ;
	    RECT 85.4000 104.1000 85.8000 104.2000 ;
	    RECT 84.6000 103.8000 85.8000 104.1000 ;
	    RECT 90.2000 104.1000 90.6000 104.2000 ;
	    RECT 92.6000 104.1000 93.0000 104.2000 ;
	    RECT 99.0000 104.1000 99.4000 104.2000 ;
	    RECT 90.2000 103.8000 91.3000 104.1000 ;
	    RECT 92.6000 103.8000 99.4000 104.1000 ;
	    RECT 131.8000 104.1000 132.2000 104.2000 ;
	    RECT 145.4000 104.1000 145.8000 104.2000 ;
	    RECT 131.8000 103.8000 145.8000 104.1000 ;
	    RECT 159.0000 104.1000 159.4000 104.2000 ;
	    RECT 165.4000 104.1000 165.8000 104.2000 ;
	    RECT 159.0000 103.8000 165.8000 104.1000 ;
	    RECT 91.0000 103.2000 91.3000 103.8000 ;
	    RECT 2.2000 103.1000 2.6000 103.2000 ;
	    RECT 3.0000 103.1000 3.4000 103.2000 ;
	    RECT 2.2000 102.8000 3.4000 103.1000 ;
	    RECT 50.2000 103.1000 50.6000 103.2000 ;
	    RECT 66.2000 103.1000 66.6000 103.2000 ;
	    RECT 50.2000 102.8000 66.6000 103.1000 ;
	    RECT 67.0000 103.1000 67.4000 103.2000 ;
	    RECT 79.0000 103.1000 79.4000 103.2000 ;
	    RECT 67.0000 102.8000 79.4000 103.1000 ;
	    RECT 85.4000 103.1000 85.8000 103.2000 ;
	    RECT 87.8000 103.1000 88.2000 103.2000 ;
	    RECT 85.4000 102.8000 88.2000 103.1000 ;
	    RECT 91.0000 102.8000 91.4000 103.2000 ;
	    RECT 96.6000 103.1000 97.0000 103.2000 ;
	    RECT 108.6000 103.1000 109.0000 103.2000 ;
	    RECT 96.6000 102.8000 109.0000 103.1000 ;
	    RECT 133.4000 103.1000 133.8000 103.2000 ;
	    RECT 137.4000 103.1000 137.8000 103.2000 ;
	    RECT 133.4000 102.8000 137.8000 103.1000 ;
	    RECT 3.0000 102.2000 3.3000 102.8000 ;
	    RECT 3.0000 101.8000 3.4000 102.2000 ;
	    RECT 71.0000 102.1000 71.4000 102.2000 ;
	    RECT 97.4000 102.1000 97.8000 102.2000 ;
	    RECT 70.2000 101.8000 97.8000 102.1000 ;
	    RECT 123.8000 102.1000 124.2000 102.2000 ;
	    RECT 126.2000 102.1000 126.6000 102.2000 ;
	    RECT 135.8000 102.1000 136.2000 102.2000 ;
	    RECT 138.2000 102.1000 138.6000 102.2000 ;
	    RECT 123.8000 101.8000 138.6000 102.1000 ;
	    RECT 39.8000 101.1000 40.2000 101.2000 ;
	    RECT 57.4000 101.1000 57.8000 101.2000 ;
	    RECT 39.8000 100.8000 57.8000 101.1000 ;
	    RECT 82.2000 101.1000 82.6000 101.2000 ;
	    RECT 114.2000 101.1000 114.6000 101.2000 ;
	    RECT 82.2000 100.8000 114.6000 101.1000 ;
	    RECT 124.6000 101.1000 125.0000 101.2000 ;
	    RECT 136.6000 101.1000 137.0000 101.2000 ;
	    RECT 124.6000 100.8000 137.0000 101.1000 ;
	    RECT 47.8000 100.1000 48.2000 100.2000 ;
	    RECT 58.2000 100.1000 58.6000 100.2000 ;
	    RECT 47.8000 99.8000 58.6000 100.1000 ;
	    RECT 79.0000 100.1000 79.4000 100.2000 ;
	    RECT 88.6000 100.1000 89.0000 100.2000 ;
	    RECT 91.0000 100.1000 91.4000 100.2000 ;
	    RECT 79.0000 99.8000 88.1000 100.1000 ;
	    RECT 88.6000 99.8000 91.4000 100.1000 ;
	    RECT 122.2000 100.1000 122.6000 100.2000 ;
	    RECT 126.2000 100.1000 126.6000 100.2000 ;
	    RECT 122.2000 99.8000 126.6000 100.1000 ;
	    RECT 127.0000 99.8000 127.4000 100.2000 ;
	    RECT 36.6000 99.1000 37.0000 99.2000 ;
	    RECT 83.0000 99.1000 83.4000 99.2000 ;
	    RECT 84.6000 99.1000 85.0000 99.2000 ;
	    RECT 87.0000 99.1000 87.4000 99.2000 ;
	    RECT 36.6000 98.8000 83.4000 99.1000 ;
	    RECT 83.8000 98.8000 87.4000 99.1000 ;
	    RECT 87.8000 99.1000 88.1000 99.8000 ;
	    RECT 109.4000 99.1000 109.8000 99.2000 ;
	    RECT 87.8000 98.8000 109.8000 99.1000 ;
	    RECT 122.2000 99.1000 122.6000 99.2000 ;
	    RECT 127.0000 99.1000 127.3000 99.8000 ;
	    RECT 122.2000 98.8000 127.3000 99.1000 ;
	    RECT 138.2000 99.1000 138.6000 99.2000 ;
	    RECT 142.2000 99.1000 142.6000 99.2000 ;
	    RECT 138.2000 98.8000 142.6000 99.1000 ;
	    RECT 74.2000 97.8000 74.6000 98.2000 ;
	    RECT 85.4000 97.8000 85.8000 98.2000 ;
	    RECT 167.0000 98.1000 167.4000 98.2000 ;
	    RECT 167.8000 98.1000 168.2000 98.2000 ;
	    RECT 167.0000 97.8000 168.2000 98.1000 ;
	    RECT 10.2000 97.1000 10.6000 97.2000 ;
	    RECT 5.4000 96.8000 10.6000 97.1000 ;
	    RECT 17.4000 97.1000 17.8000 97.2000 ;
	    RECT 20.6000 97.1000 21.0000 97.2000 ;
	    RECT 17.4000 96.8000 21.0000 97.1000 ;
	    RECT 23.0000 96.8000 23.4000 97.2000 ;
	    RECT 28.6000 97.1000 29.0000 97.2000 ;
	    RECT 30.2000 97.1000 30.6000 97.2000 ;
	    RECT 28.6000 96.8000 30.6000 97.1000 ;
	    RECT 35.0000 97.1000 35.4000 97.2000 ;
	    RECT 35.8000 97.1000 36.2000 97.2000 ;
	    RECT 35.0000 96.8000 36.2000 97.1000 ;
	    RECT 42.2000 97.1000 42.6000 97.2000 ;
	    RECT 46.2000 97.1000 46.6000 97.2000 ;
	    RECT 42.2000 96.8000 46.6000 97.1000 ;
	    RECT 47.8000 96.8000 48.2000 97.2000 ;
	    RECT 52.6000 97.1000 53.0000 97.2000 ;
	    RECT 57.4000 97.1000 57.8000 97.2000 ;
	    RECT 52.6000 96.8000 57.8000 97.1000 ;
	    RECT 60.6000 97.1000 61.0000 97.2000 ;
	    RECT 69.4000 97.1000 69.8000 97.2000 ;
	    RECT 60.6000 96.8000 69.8000 97.1000 ;
	    RECT 71.8000 97.1000 72.2000 97.2000 ;
	    RECT 74.2000 97.1000 74.5000 97.8000 ;
	    RECT 71.8000 96.8000 74.5000 97.1000 ;
	    RECT 77.4000 97.1000 77.8000 97.2000 ;
	    RECT 81.4000 97.1000 81.8000 97.2000 ;
	    RECT 77.4000 96.8000 81.8000 97.1000 ;
	    RECT 83.8000 97.1000 84.2000 97.2000 ;
	    RECT 85.4000 97.1000 85.7000 97.8000 ;
	    RECT 83.8000 96.8000 85.7000 97.1000 ;
	    RECT 91.8000 97.1000 92.2000 97.2000 ;
	    RECT 106.2000 97.1000 106.6000 97.2000 ;
	    RECT 91.8000 96.8000 106.6000 97.1000 ;
	    RECT 5.4000 96.2000 5.7000 96.8000 ;
	    RECT 5.4000 95.8000 5.8000 96.2000 ;
	    RECT 13.4000 96.1000 13.8000 96.2000 ;
	    RECT 23.0000 96.1000 23.3000 96.8000 ;
	    RECT 47.8000 96.2000 48.1000 96.8000 ;
	    RECT 23.8000 96.1000 24.2000 96.2000 ;
	    RECT 25.4000 96.1000 25.8000 96.2000 ;
	    RECT 13.4000 95.8000 25.8000 96.1000 ;
	    RECT 27.0000 95.8000 27.4000 96.2000 ;
	    RECT 32.6000 95.8000 33.0000 96.2000 ;
	    RECT 45.4000 95.8000 45.8000 96.2000 ;
	    RECT 47.8000 96.1000 48.2000 96.2000 ;
	    RECT 55.8000 96.1000 56.2000 96.2000 ;
	    RECT 47.8000 95.8000 56.2000 96.1000 ;
	    RECT 66.2000 96.1000 66.6000 96.2000 ;
	    RECT 71.0000 96.1000 71.4000 96.2000 ;
	    RECT 66.2000 95.8000 71.4000 96.1000 ;
	    RECT 75.0000 96.1000 75.4000 96.2000 ;
	    RECT 76.6000 96.1000 77.0000 96.2000 ;
	    RECT 75.0000 95.8000 77.0000 96.1000 ;
	    RECT 80.6000 96.1000 81.0000 96.2000 ;
	    RECT 83.8000 96.1000 84.2000 96.2000 ;
	    RECT 80.6000 95.8000 84.2000 96.1000 ;
	    RECT 99.8000 95.8000 100.2000 96.2000 ;
	    RECT 144.6000 96.1000 145.0000 96.2000 ;
	    RECT 151.0000 96.1000 151.4000 96.2000 ;
	    RECT 144.6000 95.8000 151.4000 96.1000 ;
	    RECT 7.8000 95.1000 8.2000 95.2000 ;
	    RECT 13.4000 95.1000 13.8000 95.2000 ;
	    RECT 15.8000 95.1000 16.2000 95.2000 ;
	    RECT 17.4000 95.1000 17.8000 95.2000 ;
	    RECT 7.8000 94.8000 17.8000 95.1000 ;
	    RECT 24.6000 95.1000 25.0000 95.2000 ;
	    RECT 27.0000 95.1000 27.3000 95.8000 ;
	    RECT 29.4000 95.1000 29.8000 95.2000 ;
	    RECT 24.6000 94.8000 27.3000 95.1000 ;
	    RECT 28.6000 94.8000 29.8000 95.1000 ;
	    RECT 31.0000 95.1000 31.4000 95.2000 ;
	    RECT 32.6000 95.1000 32.9000 95.8000 ;
	    RECT 31.0000 94.8000 32.9000 95.1000 ;
	    RECT 36.6000 95.1000 37.0000 95.2000 ;
	    RECT 37.4000 95.1000 37.8000 95.2000 ;
	    RECT 36.6000 94.8000 37.8000 95.1000 ;
	    RECT 43.8000 94.8000 44.2000 95.2000 ;
	    RECT 45.4000 95.1000 45.7000 95.8000 ;
	    RECT 99.8000 95.2000 100.1000 95.8000 ;
	    RECT 47.0000 95.1000 47.4000 95.2000 ;
	    RECT 56.6000 95.1000 57.0000 95.2000 ;
	    RECT 45.4000 94.8000 47.4000 95.1000 ;
	    RECT 55.8000 94.8000 57.0000 95.1000 ;
	    RECT 68.6000 95.1000 69.0000 95.2000 ;
	    RECT 74.2000 95.1000 74.6000 95.2000 ;
	    RECT 68.6000 94.8000 74.6000 95.1000 ;
	    RECT 79.8000 95.1000 80.2000 95.2000 ;
	    RECT 81.4000 95.1000 81.8000 95.2000 ;
	    RECT 79.8000 94.8000 81.8000 95.1000 ;
	    RECT 86.2000 95.1000 86.6000 95.2000 ;
	    RECT 97.4000 95.1000 97.8000 95.2000 ;
	    RECT 86.2000 94.8000 97.8000 95.1000 ;
	    RECT 99.8000 94.8000 100.2000 95.2000 ;
	    RECT 102.2000 95.1000 102.6000 95.2000 ;
	    RECT 102.2000 94.8000 121.0000 95.1000 ;
	    RECT 28.6000 94.2000 28.9000 94.8000 ;
	    RECT 11.8000 94.1000 12.2000 94.2000 ;
	    RECT 22.2000 94.1000 22.6000 94.2000 ;
	    RECT 9.4000 93.8000 12.2000 94.1000 ;
	    RECT 15.8000 93.8000 22.6000 94.1000 ;
	    RECT 25.4000 93.8000 25.8000 94.2000 ;
	    RECT 28.6000 93.8000 29.0000 94.2000 ;
	    RECT 37.4000 94.1000 37.8000 94.2000 ;
	    RECT 42.2000 94.1000 42.6000 94.2000 ;
	    RECT 37.4000 93.8000 42.6000 94.1000 ;
	    RECT 43.8000 94.1000 44.1000 94.8000 ;
	    RECT 55.8000 94.2000 56.1000 94.8000 ;
	    RECT 120.6000 94.7000 121.0000 94.8000 ;
	    RECT 135.0000 94.8000 135.4000 95.2000 ;
	    RECT 151.0000 94.8000 151.4000 95.2000 ;
	    RECT 152.6000 95.1000 153.0000 95.2000 ;
	    RECT 155.8000 95.1000 156.2000 95.2000 ;
	    RECT 152.6000 94.8000 156.2000 95.1000 ;
	    RECT 44.6000 94.1000 45.0000 94.2000 ;
	    RECT 51.8000 94.1000 52.2000 94.2000 ;
	    RECT 43.8000 93.8000 52.2000 94.1000 ;
	    RECT 55.8000 93.8000 56.2000 94.2000 ;
	    RECT 70.2000 94.1000 70.6000 94.2000 ;
	    RECT 71.8000 94.1000 72.2000 94.2000 ;
	    RECT 69.4000 93.8000 72.2000 94.1000 ;
	    RECT 104.6000 94.1000 105.0000 94.2000 ;
	    RECT 105.4000 94.1000 105.8000 94.2000 ;
	    RECT 104.6000 93.8000 105.8000 94.1000 ;
	    RECT 109.4000 94.1000 109.8000 94.2000 ;
	    RECT 110.2000 94.1000 110.6000 94.2000 ;
	    RECT 109.4000 93.8000 110.6000 94.1000 ;
	    RECT 115.8000 94.1000 116.2000 94.2000 ;
	    RECT 132.6000 94.1000 133.0000 94.2000 ;
	    RECT 115.8000 93.8000 133.0000 94.1000 ;
	    RECT 135.0000 94.1000 135.3000 94.8000 ;
	    RECT 151.0000 94.1000 151.3000 94.8000 ;
	    RECT 152.6000 94.1000 152.9000 94.8000 ;
	    RECT 171.0000 94.1000 171.4000 94.2000 ;
	    RECT 135.0000 93.8000 152.9000 94.1000 ;
	    RECT 168.6000 93.8000 171.4000 94.1000 ;
	    RECT 9.4000 93.2000 9.7000 93.8000 ;
	    RECT 15.8000 93.2000 16.1000 93.8000 ;
	    RECT 9.4000 92.8000 9.8000 93.2000 ;
	    RECT 15.8000 92.8000 16.2000 93.2000 ;
	    RECT 25.4000 93.1000 25.7000 93.8000 ;
	    RECT 34.2000 93.1000 34.6000 93.2000 ;
	    RECT 25.4000 92.8000 34.6000 93.1000 ;
	    RECT 75.0000 93.1000 75.4000 93.2000 ;
	    RECT 75.8000 93.1000 76.2000 93.2000 ;
	    RECT 83.8000 93.1000 84.2000 93.2000 ;
	    RECT 86.2000 93.1000 86.6000 93.2000 ;
	    RECT 91.0000 93.1000 91.4000 93.2000 ;
	    RECT 92.6000 93.1000 93.0000 93.2000 ;
	    RECT 75.0000 92.8000 93.0000 93.1000 ;
	    RECT 103.8000 93.1000 104.2000 93.2000 ;
	    RECT 104.6000 93.1000 105.0000 93.2000 ;
	    RECT 103.8000 92.8000 105.0000 93.1000 ;
	    RECT 109.4000 93.1000 109.8000 93.2000 ;
	    RECT 113.4000 93.1000 113.8000 93.2000 ;
	    RECT 115.8000 93.1000 116.2000 93.2000 ;
	    RECT 109.4000 92.8000 116.2000 93.1000 ;
	    RECT 139.0000 93.1000 139.4000 93.2000 ;
	    RECT 139.8000 93.1000 140.2000 93.2000 ;
	    RECT 151.8000 93.1000 152.2000 93.2000 ;
	    RECT 163.0000 93.1000 163.4000 93.2000 ;
	    RECT 168.6000 93.1000 168.9000 93.8000 ;
	    RECT 139.0000 92.8000 140.2000 93.1000 ;
	    RECT 142.2000 92.8000 168.9000 93.1000 ;
	    RECT 171.8000 92.8000 172.2000 93.2000 ;
	    RECT 142.2000 92.2000 142.5000 92.8000 ;
	    RECT 171.8000 92.2000 172.1000 92.8000 ;
	    RECT 86.2000 92.1000 86.6000 92.2000 ;
	    RECT 87.8000 92.1000 88.2000 92.2000 ;
	    RECT 86.2000 91.8000 88.2000 92.1000 ;
	    RECT 99.0000 92.1000 99.4000 92.2000 ;
	    RECT 99.8000 92.1000 100.2000 92.2000 ;
	    RECT 111.8000 92.1000 112.2000 92.2000 ;
	    RECT 115.8000 92.1000 116.2000 92.2000 ;
	    RECT 99.0000 91.8000 100.2000 92.1000 ;
	    RECT 111.0000 91.8000 116.2000 92.1000 ;
	    RECT 116.6000 91.8000 117.0000 92.2000 ;
	    RECT 142.2000 91.8000 142.6000 92.2000 ;
	    RECT 151.0000 92.1000 151.4000 92.2000 ;
	    RECT 163.0000 92.1000 163.4000 92.2000 ;
	    RECT 151.0000 91.8000 163.4000 92.1000 ;
	    RECT 171.8000 91.8000 172.2000 92.2000 ;
	    RECT 116.6000 91.2000 116.9000 91.8000 ;
	    RECT 116.6000 90.8000 117.0000 91.2000 ;
	    RECT 115.8000 90.1000 116.2000 90.2000 ;
	    RECT 125.4000 90.1000 125.8000 90.2000 ;
	    RECT 115.8000 89.8000 125.8000 90.1000 ;
	    RECT 128.6000 90.1000 129.0000 90.2000 ;
	    RECT 142.2000 90.1000 142.6000 90.2000 ;
	    RECT 128.6000 89.8000 142.6000 90.1000 ;
	    RECT 146.2000 90.1000 146.6000 90.2000 ;
	    RECT 152.6000 90.1000 153.0000 90.2000 ;
	    RECT 146.2000 89.8000 153.0000 90.1000 ;
	    RECT 155.0000 90.1000 155.4000 90.2000 ;
	    RECT 171.0000 90.1000 171.4000 90.2000 ;
	    RECT 155.0000 89.8000 171.4000 90.1000 ;
	    RECT 6.2000 88.8000 6.6000 89.2000 ;
	    RECT 11.8000 89.1000 12.2000 89.2000 ;
	    RECT 23.8000 89.1000 24.2000 89.2000 ;
	    RECT 11.8000 88.8000 24.2000 89.1000 ;
	    RECT 118.2000 89.1000 118.6000 89.2000 ;
	    RECT 119.0000 89.1000 119.4000 89.2000 ;
	    RECT 118.2000 88.8000 119.4000 89.1000 ;
	    RECT 136.6000 89.1000 137.0000 89.2000 ;
	    RECT 140.6000 89.1000 141.0000 89.2000 ;
	    RECT 136.6000 88.8000 141.0000 89.1000 ;
	    RECT 170.2000 89.1000 170.6000 89.2000 ;
	    RECT 172.6000 89.1000 173.0000 89.2000 ;
	    RECT 170.2000 88.8000 173.0000 89.1000 ;
	    RECT 2.2000 88.1000 2.6000 88.2000 ;
	    RECT 6.2000 88.1000 6.5000 88.8000 ;
	    RECT 2.2000 87.8000 6.5000 88.1000 ;
	    RECT 8.6000 87.8000 9.0000 88.2000 ;
	    RECT 17.4000 88.1000 17.8000 88.2000 ;
	    RECT 19.0000 88.1000 19.4000 88.2000 ;
	    RECT 17.4000 87.8000 19.4000 88.1000 ;
	    RECT 23.0000 88.1000 23.4000 88.2000 ;
	    RECT 26.2000 88.1000 26.6000 88.2000 ;
	    RECT 23.0000 87.8000 26.6000 88.1000 ;
	    RECT 31.0000 88.1000 31.4000 88.2000 ;
	    RECT 32.6000 88.1000 33.0000 88.2000 ;
	    RECT 31.0000 87.8000 33.0000 88.1000 ;
	    RECT 34.2000 88.1000 34.6000 88.2000 ;
	    RECT 35.8000 88.1000 36.2000 88.2000 ;
	    RECT 36.6000 88.1000 37.0000 88.2000 ;
	    RECT 34.2000 87.8000 37.0000 88.1000 ;
	    RECT 38.2000 88.1000 38.6000 88.2000 ;
	    RECT 43.8000 88.1000 44.2000 88.2000 ;
	    RECT 38.2000 87.8000 44.2000 88.1000 ;
	    RECT 48.6000 88.1000 49.0000 88.2000 ;
	    RECT 51.8000 88.1000 52.2000 88.2000 ;
	    RECT 58.2000 88.1000 58.6000 88.2000 ;
	    RECT 66.2000 88.1000 66.6000 88.2000 ;
	    RECT 48.6000 87.8000 66.6000 88.1000 ;
	    RECT 75.0000 88.1000 75.4000 88.2000 ;
	    RECT 93.4000 88.1000 93.8000 88.2000 ;
	    RECT 75.0000 87.8000 93.8000 88.1000 ;
	    RECT 96.6000 88.1000 97.0000 88.2000 ;
	    RECT 99.0000 88.1000 99.4000 88.2000 ;
	    RECT 96.6000 87.8000 99.4000 88.1000 ;
	    RECT 101.4000 88.1000 101.8000 88.2000 ;
	    RECT 103.8000 88.1000 104.2000 88.2000 ;
	    RECT 117.4000 88.1000 117.8000 88.2000 ;
	    RECT 101.4000 87.8000 117.8000 88.1000 ;
	    RECT 129.4000 87.8000 129.8000 88.2000 ;
	    RECT 143.8000 87.8000 144.2000 88.2000 ;
	    RECT 158.2000 88.1000 158.6000 88.2000 ;
	    RECT 172.6000 88.1000 173.0000 88.2000 ;
	    RECT 158.2000 87.8000 173.0000 88.1000 ;
	    RECT 8.6000 87.1000 8.9000 87.8000 ;
	    RECT 11.0000 87.1000 11.4000 87.2000 ;
	    RECT 8.6000 86.8000 11.4000 87.1000 ;
	    RECT 19.0000 87.1000 19.4000 87.2000 ;
	    RECT 19.8000 87.1000 20.2000 87.2000 ;
	    RECT 19.0000 86.8000 20.2000 87.1000 ;
	    RECT 22.2000 86.8000 22.6000 87.2000 ;
	    RECT 41.4000 86.8000 41.8000 87.2000 ;
	    RECT 53.4000 86.8000 53.8000 87.2000 ;
	    RECT 72.6000 87.1000 73.0000 87.2000 ;
	    RECT 75.8000 87.1000 76.2000 87.2000 ;
	    RECT 72.6000 86.8000 76.2000 87.1000 ;
	    RECT 82.2000 87.1000 82.6000 87.2000 ;
	    RECT 99.8000 87.1000 100.2000 87.2000 ;
	    RECT 82.2000 86.8000 100.2000 87.1000 ;
	    RECT 100.6000 86.8000 101.0000 87.2000 ;
	    RECT 113.4000 87.1000 113.8000 87.2000 ;
	    RECT 119.8000 87.1000 120.2000 87.2000 ;
	    RECT 123.0000 87.1000 123.4000 87.2000 ;
	    RECT 129.4000 87.1000 129.7000 87.8000 ;
	    RECT 113.4000 86.8000 129.7000 87.1000 ;
	    RECT 143.8000 87.1000 144.1000 87.8000 ;
	    RECT 147.8000 87.1000 148.2000 87.2000 ;
	    RECT 143.8000 86.8000 148.2000 87.1000 ;
	    RECT 158.2000 87.1000 158.6000 87.2000 ;
	    RECT 163.0000 87.1000 163.4000 87.2000 ;
	    RECT 167.0000 87.1000 167.4000 87.2000 ;
	    RECT 158.2000 86.8000 167.4000 87.1000 ;
	    RECT 3.8000 86.1000 4.2000 86.2000 ;
	    RECT 13.4000 86.1000 13.8000 86.2000 ;
	    RECT 3.8000 85.8000 13.8000 86.1000 ;
	    RECT 22.2000 85.8000 22.5000 86.8000 ;
	    RECT 24.6000 86.1000 25.0000 86.2000 ;
	    RECT 25.4000 86.1000 25.8000 86.2000 ;
	    RECT 24.6000 85.8000 25.8000 86.1000 ;
	    RECT 26.2000 86.1000 26.6000 86.2000 ;
	    RECT 27.8000 86.1000 28.2000 86.2000 ;
	    RECT 26.2000 85.8000 28.2000 86.1000 ;
	    RECT 29.4000 86.1000 29.8000 86.2000 ;
	    RECT 30.2000 86.1000 30.6000 86.2000 ;
	    RECT 29.4000 85.8000 30.6000 86.1000 ;
	    RECT 31.8000 86.1000 32.2000 86.2000 ;
	    RECT 34.2000 86.1000 34.6000 86.2000 ;
	    RECT 31.8000 85.8000 34.6000 86.1000 ;
	    RECT 35.0000 86.1000 35.4000 86.2000 ;
	    RECT 41.4000 86.1000 41.7000 86.8000 ;
	    RECT 35.0000 85.8000 41.7000 86.1000 ;
	    RECT 43.8000 86.1000 44.2000 86.2000 ;
	    RECT 53.4000 86.1000 53.7000 86.8000 ;
	    RECT 100.6000 86.2000 100.9000 86.8000 ;
	    RECT 55.0000 86.1000 55.4000 86.2000 ;
	    RECT 43.8000 85.8000 44.9000 86.1000 ;
	    RECT 53.4000 85.8000 55.4000 86.1000 ;
	    RECT 62.2000 86.1000 62.6000 86.2000 ;
	    RECT 71.8000 86.1000 72.2000 86.2000 ;
	    RECT 62.2000 85.8000 72.2000 86.1000 ;
	    RECT 74.2000 86.1000 74.6000 86.2000 ;
	    RECT 75.0000 86.1000 75.4000 86.2000 ;
	    RECT 74.2000 85.8000 75.4000 86.1000 ;
	    RECT 76.6000 85.8000 77.0000 86.2000 ;
	    RECT 78.2000 86.1000 78.6000 86.2000 ;
	    RECT 79.0000 86.1000 79.4000 86.2000 ;
	    RECT 78.2000 85.8000 79.4000 86.1000 ;
	    RECT 81.4000 85.8000 81.8000 86.2000 ;
	    RECT 83.0000 86.1000 83.4000 86.2000 ;
	    RECT 83.8000 86.1000 84.2000 86.2000 ;
	    RECT 83.0000 85.8000 84.2000 86.1000 ;
	    RECT 87.0000 85.8000 87.4000 86.2000 ;
	    RECT 95.8000 86.1000 96.2000 86.2000 ;
	    RECT 96.6000 86.1000 97.0000 86.2000 ;
	    RECT 95.8000 85.8000 97.0000 86.1000 ;
	    RECT 100.6000 85.8000 101.0000 86.2000 ;
	    RECT 111.8000 86.1000 112.2000 86.2000 ;
	    RECT 129.4000 86.1000 129.8000 86.2000 ;
	    RECT 111.8000 85.8000 129.8000 86.1000 ;
	    RECT 165.4000 85.8000 165.8000 86.2000 ;
	    RECT 167.8000 86.1000 168.2000 86.2000 ;
	    RECT 170.2000 86.1000 170.6000 86.2000 ;
	    RECT 167.8000 85.8000 170.6000 86.1000 ;
	    RECT 44.6000 85.2000 44.9000 85.8000 ;
	    RECT 76.6000 85.2000 76.9000 85.8000 ;
	    RECT 81.4000 85.2000 81.7000 85.8000 ;
	    RECT 87.0000 85.2000 87.3000 85.8000 ;
	    RECT 165.4000 85.2000 165.7000 85.8000 ;
	    RECT 3.0000 84.8000 3.4000 85.2000 ;
	    RECT 17.4000 85.1000 17.8000 85.2000 ;
	    RECT 18.2000 85.1000 18.6000 85.2000 ;
	    RECT 17.4000 84.8000 18.6000 85.1000 ;
	    RECT 23.8000 85.1000 24.2000 85.2000 ;
	    RECT 31.0000 85.1000 31.4000 85.2000 ;
	    RECT 23.8000 84.8000 31.4000 85.1000 ;
	    RECT 44.6000 84.8000 45.0000 85.2000 ;
	    RECT 48.6000 85.1000 49.0000 85.2000 ;
	    RECT 49.4000 85.1000 49.8000 85.2000 ;
	    RECT 48.6000 84.8000 49.8000 85.1000 ;
	    RECT 51.0000 85.1000 51.4000 85.2000 ;
	    RECT 57.4000 85.1000 57.8000 85.2000 ;
	    RECT 73.4000 85.1000 73.8000 85.2000 ;
	    RECT 51.0000 84.8000 73.8000 85.1000 ;
	    RECT 76.6000 85.1000 77.0000 85.2000 ;
	    RECT 79.0000 85.1000 79.4000 85.2000 ;
	    RECT 76.6000 84.8000 79.4000 85.1000 ;
	    RECT 81.4000 84.8000 81.8000 85.2000 ;
	    RECT 87.0000 84.8000 87.4000 85.2000 ;
	    RECT 91.0000 85.1000 91.4000 85.2000 ;
	    RECT 92.6000 85.1000 93.0000 85.2000 ;
	    RECT 91.0000 84.8000 93.0000 85.1000 ;
	    RECT 95.0000 85.1000 95.4000 85.2000 ;
	    RECT 97.4000 85.1000 97.8000 85.2000 ;
	    RECT 95.0000 84.8000 97.8000 85.1000 ;
	    RECT 126.2000 85.1000 126.6000 85.2000 ;
	    RECT 135.0000 85.1000 135.4000 85.2000 ;
	    RECT 126.2000 84.8000 135.4000 85.1000 ;
	    RECT 144.6000 85.1000 145.0000 85.2000 ;
	    RECT 148.6000 85.1000 149.0000 85.2000 ;
	    RECT 144.6000 84.8000 149.0000 85.1000 ;
	    RECT 165.4000 84.8000 165.8000 85.2000 ;
	    RECT 3.0000 84.1000 3.3000 84.8000 ;
	    RECT 9.4000 84.1000 9.8000 84.2000 ;
	    RECT 3.0000 83.8000 9.8000 84.1000 ;
	    RECT 49.4000 84.1000 49.8000 84.2000 ;
	    RECT 55.8000 84.1000 56.2000 84.2000 ;
	    RECT 49.4000 83.8000 56.2000 84.1000 ;
	    RECT 63.0000 84.1000 63.4000 84.2000 ;
	    RECT 67.8000 84.1000 68.2000 84.2000 ;
	    RECT 63.0000 83.8000 68.2000 84.1000 ;
	    RECT 72.6000 84.1000 73.0000 84.2000 ;
	    RECT 84.6000 84.1000 85.0000 84.2000 ;
	    RECT 88.6000 84.1000 89.0000 84.2000 ;
	    RECT 72.6000 83.8000 78.5000 84.1000 ;
	    RECT 84.6000 83.8000 89.0000 84.1000 ;
	    RECT 92.6000 84.1000 93.0000 84.2000 ;
	    RECT 95.0000 84.1000 95.4000 84.2000 ;
	    RECT 92.6000 83.8000 95.4000 84.1000 ;
	    RECT 78.2000 83.2000 78.5000 83.8000 ;
	    RECT 71.8000 83.1000 72.2000 83.2000 ;
	    RECT 67.0000 82.8000 72.2000 83.1000 ;
	    RECT 78.2000 82.8000 78.6000 83.2000 ;
	    RECT 86.2000 83.1000 86.6000 83.2000 ;
	    RECT 89.4000 83.1000 89.8000 83.2000 ;
	    RECT 86.2000 82.8000 89.8000 83.1000 ;
	    RECT 91.8000 83.1000 92.2000 83.2000 ;
	    RECT 92.6000 83.1000 93.0000 83.2000 ;
	    RECT 91.8000 82.8000 93.0000 83.1000 ;
	    RECT 127.8000 83.1000 128.2000 83.2000 ;
	    RECT 133.4000 83.1000 133.8000 83.2000 ;
	    RECT 127.8000 82.8000 133.8000 83.1000 ;
	    RECT 67.0000 82.2000 67.3000 82.8000 ;
	    RECT 10.2000 82.1000 10.6000 82.2000 ;
	    RECT 13.4000 82.1000 13.8000 82.2000 ;
	    RECT 10.2000 81.8000 13.8000 82.1000 ;
	    RECT 37.4000 82.1000 37.8000 82.2000 ;
	    RECT 39.8000 82.1000 40.2000 82.2000 ;
	    RECT 37.4000 81.8000 40.2000 82.1000 ;
	    RECT 50.2000 82.1000 50.6000 82.2000 ;
	    RECT 64.6000 82.1000 65.0000 82.2000 ;
	    RECT 50.2000 81.8000 65.0000 82.1000 ;
	    RECT 67.0000 81.8000 67.4000 82.2000 ;
	    RECT 67.8000 82.1000 68.2000 82.2000 ;
	    RECT 68.6000 82.1000 69.0000 82.2000 ;
	    RECT 67.8000 81.8000 69.0000 82.1000 ;
	    RECT 69.4000 82.1000 69.8000 82.2000 ;
	    RECT 81.4000 82.1000 81.8000 82.2000 ;
	    RECT 69.4000 81.8000 81.8000 82.1000 ;
	    RECT 39.0000 81.1000 39.4000 81.2000 ;
	    RECT 42.2000 81.1000 42.6000 81.2000 ;
	    RECT 39.0000 80.8000 42.6000 81.1000 ;
	    RECT 99.8000 81.1000 100.2000 81.2000 ;
	    RECT 147.0000 81.1000 147.4000 81.2000 ;
	    RECT 99.8000 80.8000 147.4000 81.1000 ;
	    RECT 39.8000 80.1000 40.2000 80.2000 ;
	    RECT 43.8000 80.1000 44.2000 80.2000 ;
	    RECT 39.8000 79.8000 44.2000 80.1000 ;
	    RECT 46.2000 80.1000 46.6000 80.2000 ;
	    RECT 59.0000 80.1000 59.4000 80.2000 ;
	    RECT 75.0000 80.1000 75.4000 80.2000 ;
	    RECT 46.2000 79.8000 59.4000 80.1000 ;
	    RECT 63.8000 79.8000 75.4000 80.1000 ;
	    RECT 93.4000 80.1000 93.8000 80.2000 ;
	    RECT 143.8000 80.1000 144.2000 80.2000 ;
	    RECT 93.4000 79.8000 144.2000 80.1000 ;
	    RECT 59.8000 79.1000 60.2000 79.2000 ;
	    RECT 63.8000 79.1000 64.1000 79.8000 ;
	    RECT 59.0000 78.8000 64.1000 79.1000 ;
	    RECT 64.6000 79.1000 65.0000 79.2000 ;
	    RECT 69.4000 79.1000 69.8000 79.2000 ;
	    RECT 64.6000 78.8000 69.8000 79.1000 ;
	    RECT 70.2000 79.1000 70.6000 79.2000 ;
	    RECT 73.4000 79.1000 73.8000 79.2000 ;
	    RECT 70.2000 78.8000 73.8000 79.1000 ;
	    RECT 98.2000 79.1000 98.6000 79.2000 ;
	    RECT 99.8000 79.1000 100.2000 79.2000 ;
	    RECT 98.2000 78.8000 100.2000 79.1000 ;
	    RECT 136.6000 79.1000 137.0000 79.2000 ;
	    RECT 139.8000 79.1000 140.2000 79.2000 ;
	    RECT 136.6000 78.8000 140.2000 79.1000 ;
	    RECT 166.2000 79.1000 166.6000 79.2000 ;
	    RECT 169.4000 79.1000 169.8000 79.2000 ;
	    RECT 166.2000 78.8000 169.8000 79.1000 ;
	    RECT 95.0000 78.1000 95.4000 78.2000 ;
	    RECT 139.0000 78.1000 139.4000 78.2000 ;
	    RECT 95.0000 77.8000 139.4000 78.1000 ;
	    RECT 3.8000 77.1000 4.2000 77.2000 ;
	    RECT 4.6000 77.1000 5.0000 77.2000 ;
	    RECT 3.8000 76.8000 5.0000 77.1000 ;
	    RECT 44.6000 77.1000 45.0000 77.2000 ;
	    RECT 48.6000 77.1000 49.0000 77.2000 ;
	    RECT 44.6000 76.8000 49.0000 77.1000 ;
	    RECT 55.8000 77.1000 56.2000 77.2000 ;
	    RECT 63.8000 77.1000 64.2000 77.2000 ;
	    RECT 55.8000 76.8000 64.2000 77.1000 ;
	    RECT 67.8000 77.1000 68.2000 77.2000 ;
	    RECT 72.6000 77.1000 73.0000 77.2000 ;
	    RECT 67.8000 76.8000 73.0000 77.1000 ;
	    RECT 93.4000 77.1000 93.8000 77.2000 ;
	    RECT 94.2000 77.1000 94.6000 77.2000 ;
	    RECT 93.4000 76.8000 94.6000 77.1000 ;
	    RECT 95.8000 77.1000 96.2000 77.2000 ;
	    RECT 97.4000 77.1000 97.8000 77.2000 ;
	    RECT 100.6000 77.1000 101.0000 77.2000 ;
	    RECT 103.0000 77.1000 103.4000 77.2000 ;
	    RECT 95.8000 76.8000 103.4000 77.1000 ;
	    RECT 146.2000 76.8000 146.6000 77.2000 ;
	    RECT 47.8000 75.8000 48.2000 76.2000 ;
	    RECT 55.0000 76.1000 55.4000 76.2000 ;
	    RECT 59.0000 76.1000 59.4000 76.2000 ;
	    RECT 54.2000 75.8000 59.4000 76.1000 ;
	    RECT 83.0000 76.1000 83.4000 76.2000 ;
	    RECT 96.6000 76.1000 97.0000 76.2000 ;
	    RECT 136.6000 76.1000 137.0000 76.2000 ;
	    RECT 83.0000 75.8000 96.1000 76.1000 ;
	    RECT 96.6000 75.8000 137.0000 76.1000 ;
	    RECT 146.2000 76.1000 146.5000 76.8000 ;
	    RECT 155.8000 76.1000 156.2000 76.2000 ;
	    RECT 146.2000 75.8000 156.2000 76.1000 ;
	    RECT 14.2000 75.1000 14.6000 75.2000 ;
	    RECT 16.6000 75.1000 17.0000 75.2000 ;
	    RECT 14.2000 74.8000 17.0000 75.1000 ;
	    RECT 29.4000 75.1000 29.8000 75.2000 ;
	    RECT 35.8000 75.1000 36.2000 75.2000 ;
	    RECT 29.4000 74.8000 36.2000 75.1000 ;
	    RECT 47.8000 75.1000 48.1000 75.8000 ;
	    RECT 95.8000 75.2000 96.1000 75.8000 ;
	    RECT 49.4000 75.1000 49.8000 75.2000 ;
	    RECT 47.8000 74.8000 49.8000 75.1000 ;
	    RECT 73.4000 75.1000 73.8000 75.2000 ;
	    RECT 75.0000 75.1000 75.4000 75.2000 ;
	    RECT 73.4000 74.8000 75.4000 75.1000 ;
	    RECT 79.0000 75.1000 79.4000 75.2000 ;
	    RECT 94.2000 75.1000 94.6000 75.2000 ;
	    RECT 79.0000 74.8000 94.6000 75.1000 ;
	    RECT 95.8000 74.8000 96.2000 75.2000 ;
	    RECT 98.2000 75.1000 98.6000 75.2000 ;
	    RECT 139.0000 75.1000 139.4000 75.2000 ;
	    RECT 151.8000 75.1000 152.2000 75.2000 ;
	    RECT 98.2000 74.8000 116.9000 75.1000 ;
	    RECT 139.0000 74.8000 152.2000 75.1000 ;
	    RECT 116.6000 74.2000 116.9000 74.8000 ;
	    RECT 13.4000 74.1000 13.8000 74.2000 ;
	    RECT 17.4000 74.1000 17.8000 74.2000 ;
	    RECT 23.0000 74.1000 23.4000 74.2000 ;
	    RECT 10.2000 73.8000 23.4000 74.1000 ;
	    RECT 99.0000 74.1000 99.4000 74.2000 ;
	    RECT 102.2000 74.1000 102.6000 74.2000 ;
	    RECT 99.0000 73.8000 102.6000 74.1000 ;
	    RECT 116.6000 73.8000 117.0000 74.2000 ;
	    RECT 143.0000 74.1000 143.4000 74.2000 ;
	    RECT 149.4000 74.1000 149.8000 74.2000 ;
	    RECT 143.0000 73.8000 149.8000 74.1000 ;
	    RECT 152.6000 74.1000 153.0000 74.2000 ;
	    RECT 153.4000 74.1000 153.8000 74.2000 ;
	    RECT 152.6000 73.8000 153.8000 74.1000 ;
	    RECT 10.2000 73.2000 10.5000 73.8000 ;
	    RECT 2.2000 73.1000 2.6000 73.2000 ;
	    RECT 4.6000 73.1000 5.0000 73.2000 ;
	    RECT 2.2000 72.8000 5.0000 73.1000 ;
	    RECT 10.2000 72.8000 10.6000 73.2000 ;
	    RECT 31.8000 73.1000 32.2000 73.2000 ;
	    RECT 33.4000 73.1000 33.8000 73.2000 ;
	    RECT 31.8000 72.8000 33.8000 73.1000 ;
	    RECT 46.2000 73.1000 46.6000 73.2000 ;
	    RECT 48.6000 73.1000 49.0000 73.2000 ;
	    RECT 52.6000 73.1000 53.0000 73.2000 ;
	    RECT 59.0000 73.1000 59.4000 73.2000 ;
	    RECT 63.0000 73.1000 63.4000 73.2000 ;
	    RECT 46.2000 72.8000 55.3000 73.1000 ;
	    RECT 59.0000 72.8000 63.4000 73.1000 ;
	    RECT 64.6000 73.1000 65.0000 73.2000 ;
	    RECT 68.6000 73.1000 69.0000 73.2000 ;
	    RECT 64.6000 72.8000 69.0000 73.1000 ;
	    RECT 78.2000 73.1000 78.6000 73.2000 ;
	    RECT 79.8000 73.1000 80.2000 73.2000 ;
	    RECT 78.2000 72.8000 80.2000 73.1000 ;
	    RECT 103.0000 73.1000 103.4000 73.2000 ;
	    RECT 111.0000 73.1000 111.4000 73.2000 ;
	    RECT 103.0000 72.8000 111.4000 73.1000 ;
	    RECT 139.8000 73.1000 140.2000 73.2000 ;
	    RECT 143.0000 73.1000 143.3000 73.8000 ;
	    RECT 145.4000 73.1000 145.8000 73.2000 ;
	    RECT 139.8000 72.8000 145.8000 73.1000 ;
	    RECT 147.8000 73.1000 148.2000 73.2000 ;
	    RECT 148.6000 73.1000 149.0000 73.2000 ;
	    RECT 147.8000 72.8000 149.0000 73.1000 ;
	    RECT 55.0000 72.2000 55.3000 72.8000 ;
	    RECT 4.6000 72.1000 5.0000 72.2000 ;
	    RECT 15.0000 72.1000 15.4000 72.2000 ;
	    RECT 4.6000 71.8000 15.4000 72.1000 ;
	    RECT 55.0000 71.8000 55.4000 72.2000 ;
	    RECT 75.8000 72.1000 76.2000 72.2000 ;
	    RECT 82.2000 72.1000 82.6000 72.2000 ;
	    RECT 75.8000 71.8000 82.6000 72.1000 ;
	    RECT 100.6000 72.1000 101.0000 72.2000 ;
	    RECT 116.6000 72.1000 117.0000 72.2000 ;
	    RECT 100.6000 71.8000 117.0000 72.1000 ;
	    RECT 170.2000 72.1000 170.6000 72.2000 ;
	    RECT 171.0000 72.1000 171.4000 72.2000 ;
	    RECT 170.2000 71.8000 171.4000 72.1000 ;
	    RECT 5.4000 71.1000 5.8000 71.2000 ;
	    RECT 10.2000 71.1000 10.6000 71.2000 ;
	    RECT 5.4000 70.8000 10.6000 71.1000 ;
	    RECT 25.4000 71.1000 25.8000 71.2000 ;
	    RECT 30.2000 71.1000 30.6000 71.2000 ;
	    RECT 25.4000 70.8000 30.6000 71.1000 ;
	    RECT 46.2000 71.1000 46.6000 71.2000 ;
	    RECT 67.8000 71.1000 68.2000 71.2000 ;
	    RECT 46.2000 70.8000 68.2000 71.1000 ;
	    RECT 96.6000 71.1000 97.0000 71.2000 ;
	    RECT 97.4000 71.1000 97.8000 71.2000 ;
	    RECT 96.6000 70.8000 97.8000 71.1000 ;
	    RECT 95.0000 69.1000 95.4000 69.2000 ;
	    RECT 101.4000 69.1000 101.8000 69.2000 ;
	    RECT 95.0000 68.8000 101.8000 69.1000 ;
	    RECT 109.4000 69.1000 109.8000 69.2000 ;
	    RECT 111.8000 69.1000 112.2000 69.2000 ;
	    RECT 109.4000 68.8000 112.2000 69.1000 ;
	    RECT 142.2000 69.1000 142.6000 69.2000 ;
	    RECT 155.0000 69.1000 155.4000 69.2000 ;
	    RECT 158.2000 69.1000 158.6000 69.2000 ;
	    RECT 142.2000 68.8000 158.6000 69.1000 ;
	    RECT 7.8000 68.1000 8.2000 68.2000 ;
	    RECT 11.0000 68.1000 11.4000 68.2000 ;
	    RECT 7.8000 67.8000 11.4000 68.1000 ;
	    RECT 13.4000 68.1000 13.8000 68.2000 ;
	    RECT 21.4000 68.1000 21.8000 68.2000 ;
	    RECT 13.4000 67.8000 21.8000 68.1000 ;
	    RECT 23.0000 68.1000 23.4000 68.2000 ;
	    RECT 26.2000 68.1000 26.6000 68.2000 ;
	    RECT 23.0000 67.8000 26.6000 68.1000 ;
	    RECT 67.0000 68.1000 67.4000 68.2000 ;
	    RECT 71.8000 68.1000 72.2000 68.2000 ;
	    RECT 76.6000 68.1000 77.0000 68.2000 ;
	    RECT 67.0000 67.8000 77.0000 68.1000 ;
	    RECT 77.4000 68.1000 77.8000 68.2000 ;
	    RECT 80.6000 68.1000 81.0000 68.2000 ;
	    RECT 89.4000 68.1000 89.8000 68.2000 ;
	    RECT 96.6000 68.1000 97.0000 68.2000 ;
	    RECT 98.2000 68.1000 98.6000 68.2000 ;
	    RECT 110.2000 68.1000 110.6000 68.2000 ;
	    RECT 77.4000 67.8000 110.6000 68.1000 ;
	    RECT 120.6000 68.1000 121.0000 68.2000 ;
	    RECT 127.8000 68.1000 128.2000 68.2000 ;
	    RECT 133.4000 68.1000 133.8000 68.2000 ;
	    RECT 120.6000 67.8000 133.8000 68.1000 ;
	    RECT 153.4000 67.8000 153.8000 68.2000 ;
	    RECT 8.6000 67.1000 9.0000 67.2000 ;
	    RECT 9.4000 67.1000 9.8000 67.2000 ;
	    RECT 7.8000 66.8000 9.8000 67.1000 ;
	    RECT 10.2000 67.1000 10.6000 67.2000 ;
	    RECT 12.6000 67.1000 13.0000 67.2000 ;
	    RECT 10.2000 66.8000 13.0000 67.1000 ;
	    RECT 19.8000 66.8000 20.2000 67.2000 ;
	    RECT 29.4000 66.8000 29.8000 67.2000 ;
	    RECT 42.2000 67.1000 42.6000 67.2000 ;
	    RECT 44.6000 67.1000 45.0000 67.2000 ;
	    RECT 42.2000 66.8000 45.0000 67.1000 ;
	    RECT 50.2000 67.1000 50.6000 67.2000 ;
	    RECT 72.6000 67.1000 73.0000 67.2000 ;
	    RECT 93.4000 67.1000 93.8000 67.2000 ;
	    RECT 50.2000 66.8000 53.7000 67.1000 ;
	    RECT 72.6000 66.8000 93.8000 67.1000 ;
	    RECT 95.8000 67.1000 96.2000 67.2000 ;
	    RECT 99.0000 67.1000 99.4000 67.2000 ;
	    RECT 95.8000 66.8000 99.4000 67.1000 ;
	    RECT 110.2000 67.1000 110.6000 67.2000 ;
	    RECT 115.0000 67.1000 115.4000 67.2000 ;
	    RECT 110.2000 66.8000 115.4000 67.1000 ;
	    RECT 118.2000 67.1000 118.6000 67.2000 ;
	    RECT 120.6000 67.1000 120.9000 67.8000 ;
	    RECT 118.2000 66.8000 120.9000 67.1000 ;
	    RECT 128.6000 66.8000 129.0000 67.2000 ;
	    RECT 142.2000 67.1000 142.6000 67.2000 ;
	    RECT 131.8000 66.8000 142.6000 67.1000 ;
	    RECT 153.4000 67.1000 153.7000 67.8000 ;
	    RECT 159.0000 67.1000 159.4000 67.2000 ;
	    RECT 153.4000 66.8000 159.4000 67.1000 ;
	    RECT 15.0000 66.1000 15.4000 66.2000 ;
	    RECT 15.8000 66.1000 16.2000 66.2000 ;
	    RECT 15.0000 65.8000 16.2000 66.1000 ;
	    RECT 17.4000 66.1000 17.8000 66.2000 ;
	    RECT 19.8000 66.1000 20.1000 66.8000 ;
	    RECT 17.4000 65.8000 20.1000 66.1000 ;
	    RECT 29.4000 66.1000 29.7000 66.8000 ;
	    RECT 44.6000 66.2000 44.9000 66.8000 ;
	    RECT 53.4000 66.2000 53.7000 66.8000 ;
	    RECT 97.4000 66.2000 97.7000 66.8000 ;
	    RECT 30.2000 66.1000 30.6000 66.2000 ;
	    RECT 29.4000 65.8000 30.6000 66.1000 ;
	    RECT 34.2000 65.8000 34.6000 66.2000 ;
	    RECT 44.6000 65.8000 45.0000 66.2000 ;
	    RECT 53.4000 65.8000 53.8000 66.2000 ;
	    RECT 58.2000 66.1000 58.6000 66.2000 ;
	    RECT 55.0000 65.8000 58.6000 66.1000 ;
	    RECT 59.0000 66.1000 59.4000 66.2000 ;
	    RECT 92.6000 66.1000 93.0000 66.2000 ;
	    RECT 59.0000 65.8000 93.0000 66.1000 ;
	    RECT 95.8000 65.8000 96.2000 66.2000 ;
	    RECT 97.4000 65.8000 97.8000 66.2000 ;
	    RECT 99.8000 66.1000 100.2000 66.2000 ;
	    RECT 104.6000 66.1000 105.0000 66.3000 ;
	    RECT 99.8000 65.9000 105.0000 66.1000 ;
	    RECT 128.6000 66.1000 128.9000 66.8000 ;
	    RECT 131.8000 66.2000 132.1000 66.8000 ;
	    RECT 159.0000 66.2000 159.3000 66.8000 ;
	    RECT 130.2000 66.1000 130.6000 66.2000 ;
	    RECT 99.8000 65.8000 104.9000 65.9000 ;
	    RECT 128.6000 65.8000 130.6000 66.1000 ;
	    RECT 131.8000 65.8000 132.2000 66.2000 ;
	    RECT 136.6000 66.1000 137.0000 66.2000 ;
	    RECT 138.2000 66.1000 138.6000 66.2000 ;
	    RECT 136.6000 65.8000 138.6000 66.1000 ;
	    RECT 147.0000 66.1000 147.4000 66.2000 ;
	    RECT 155.0000 66.1000 155.4000 66.2000 ;
	    RECT 147.0000 65.8000 155.4000 66.1000 ;
	    RECT 159.0000 65.8000 159.4000 66.2000 ;
	    RECT 3.0000 65.1000 3.4000 65.2000 ;
	    RECT 3.8000 65.1000 4.2000 65.2000 ;
	    RECT 9.4000 65.1000 9.8000 65.2000 ;
	    RECT 26.2000 65.1000 26.6000 65.2000 ;
	    RECT 29.4000 65.1000 29.8000 65.2000 ;
	    RECT 3.0000 64.8000 29.8000 65.1000 ;
	    RECT 31.8000 65.1000 32.2000 65.2000 ;
	    RECT 34.2000 65.1000 34.5000 65.8000 ;
	    RECT 31.8000 64.8000 34.5000 65.1000 ;
	    RECT 49.4000 65.1000 49.8000 65.2000 ;
	    RECT 50.2000 65.1000 50.6000 65.2000 ;
	    RECT 55.0000 65.1000 55.3000 65.8000 ;
	    RECT 49.4000 64.8000 50.6000 65.1000 ;
	    RECT 52.6000 64.8000 55.3000 65.1000 ;
	    RECT 55.8000 65.1000 56.2000 65.2000 ;
	    RECT 78.2000 65.1000 78.6000 65.2000 ;
	    RECT 55.8000 64.8000 78.6000 65.1000 ;
	    RECT 95.8000 65.1000 96.1000 65.8000 ;
	    RECT 122.2000 65.1000 122.6000 65.2000 ;
	    RECT 95.8000 64.8000 122.6000 65.1000 ;
	    RECT 148.6000 65.1000 149.0000 65.2000 ;
	    RECT 160.6000 65.1000 161.0000 65.2000 ;
	    RECT 148.6000 64.8000 161.0000 65.1000 ;
	    RECT 52.6000 64.2000 52.9000 64.8000 ;
	    RECT 42.2000 64.1000 42.6000 64.2000 ;
	    RECT 46.2000 64.1000 46.6000 64.2000 ;
	    RECT 42.2000 63.8000 46.6000 64.1000 ;
	    RECT 52.6000 63.8000 53.0000 64.2000 ;
	    RECT 55.0000 64.1000 55.4000 64.2000 ;
	    RECT 57.4000 64.1000 57.8000 64.2000 ;
	    RECT 55.0000 63.8000 57.8000 64.1000 ;
	    RECT 58.2000 64.1000 58.6000 64.2000 ;
	    RECT 67.0000 64.1000 67.4000 64.2000 ;
	    RECT 58.2000 63.8000 67.4000 64.1000 ;
	    RECT 70.2000 64.1000 70.6000 64.2000 ;
	    RECT 81.4000 64.1000 81.8000 64.2000 ;
	    RECT 70.2000 63.8000 81.8000 64.1000 ;
	    RECT 99.0000 64.1000 99.4000 64.2000 ;
	    RECT 99.8000 64.1000 100.2000 64.2000 ;
	    RECT 99.0000 63.8000 100.2000 64.1000 ;
	    RECT 26.2000 63.1000 26.6000 63.2000 ;
	    RECT 31.0000 63.1000 31.4000 63.2000 ;
	    RECT 26.2000 62.8000 31.4000 63.1000 ;
	    RECT 31.8000 63.1000 32.2000 63.2000 ;
	    RECT 33.4000 63.1000 33.8000 63.2000 ;
	    RECT 31.8000 62.8000 33.8000 63.1000 ;
	    RECT 75.8000 63.1000 76.2000 63.2000 ;
	    RECT 97.4000 63.1000 97.8000 63.2000 ;
	    RECT 75.8000 62.8000 97.8000 63.1000 ;
	    RECT 101.4000 63.1000 101.8000 63.2000 ;
	    RECT 110.2000 63.1000 110.6000 63.2000 ;
	    RECT 101.4000 62.8000 110.6000 63.1000 ;
	    RECT 3.0000 62.1000 3.4000 62.2000 ;
	    RECT 3.8000 62.1000 4.2000 62.2000 ;
	    RECT 3.0000 61.8000 4.2000 62.1000 ;
	    RECT 79.8000 62.1000 80.2000 62.2000 ;
	    RECT 104.6000 62.1000 105.0000 62.2000 ;
	    RECT 79.8000 61.8000 105.0000 62.1000 ;
	    RECT 11.8000 61.1000 12.2000 61.2000 ;
	    RECT 13.4000 61.1000 13.8000 61.2000 ;
	    RECT 11.8000 60.8000 13.8000 61.1000 ;
	    RECT 18.2000 61.1000 18.6000 61.2000 ;
	    RECT 23.8000 61.1000 24.2000 61.2000 ;
	    RECT 18.2000 60.8000 24.2000 61.1000 ;
	    RECT 62.2000 60.1000 62.6000 60.2000 ;
	    RECT 86.2000 60.1000 86.6000 60.2000 ;
	    RECT 62.2000 59.8000 86.6000 60.1000 ;
	    RECT 20.6000 59.1000 21.0000 59.2000 ;
	    RECT 23.0000 59.1000 23.4000 59.2000 ;
	    RECT 24.6000 59.1000 25.0000 59.2000 ;
	    RECT 27.8000 59.1000 28.2000 59.2000 ;
	    RECT 20.6000 58.8000 24.1000 59.1000 ;
	    RECT 24.6000 58.8000 28.2000 59.1000 ;
	    RECT 44.6000 59.1000 45.0000 59.2000 ;
	    RECT 45.4000 59.1000 45.8000 59.2000 ;
	    RECT 44.6000 58.8000 45.8000 59.1000 ;
	    RECT 46.2000 59.1000 46.6000 59.2000 ;
	    RECT 77.4000 59.1000 77.8000 59.2000 ;
	    RECT 46.2000 58.8000 77.8000 59.1000 ;
	    RECT 103.0000 59.1000 103.4000 59.2000 ;
	    RECT 134.2000 59.1000 134.6000 59.2000 ;
	    RECT 103.0000 58.8000 134.6000 59.1000 ;
	    RECT 148.6000 58.8000 149.0000 59.2000 ;
	    RECT 3.8000 57.8000 4.2000 58.2000 ;
	    RECT 6.2000 58.1000 6.6000 58.2000 ;
	    RECT 8.6000 58.1000 9.0000 58.2000 ;
	    RECT 15.8000 58.1000 16.2000 58.2000 ;
	    RECT 17.4000 58.1000 17.8000 58.2000 ;
	    RECT 19.8000 58.1000 20.2000 58.2000 ;
	    RECT 6.2000 57.8000 20.2000 58.1000 ;
	    RECT 21.4000 58.1000 21.8000 58.2000 ;
	    RECT 22.2000 58.1000 22.6000 58.2000 ;
	    RECT 35.8000 58.1000 36.2000 58.2000 ;
	    RECT 21.4000 57.8000 22.6000 58.1000 ;
	    RECT 23.0000 57.8000 36.2000 58.1000 ;
	    RECT 52.6000 58.1000 53.0000 58.2000 ;
	    RECT 67.0000 58.1000 67.4000 58.2000 ;
	    RECT 135.8000 58.1000 136.2000 58.2000 ;
	    RECT 142.2000 58.1000 142.6000 58.2000 ;
	    RECT 52.6000 57.8000 86.5000 58.1000 ;
	    RECT 135.8000 57.8000 142.6000 58.1000 ;
	    RECT 143.0000 58.1000 143.4000 58.2000 ;
	    RECT 145.4000 58.1000 145.8000 58.2000 ;
	    RECT 143.0000 57.8000 145.8000 58.1000 ;
	    RECT 146.2000 58.1000 146.6000 58.2000 ;
	    RECT 148.6000 58.1000 148.9000 58.8000 ;
	    RECT 146.2000 57.8000 148.9000 58.1000 ;
	    RECT 3.8000 57.2000 4.1000 57.8000 ;
	    RECT 3.8000 56.8000 4.2000 57.2000 ;
	    RECT 5.4000 57.1000 5.8000 57.2000 ;
	    RECT 12.6000 57.1000 13.0000 57.2000 ;
	    RECT 5.4000 56.8000 13.0000 57.1000 ;
	    RECT 15.0000 57.1000 15.4000 57.2000 ;
	    RECT 15.8000 57.1000 16.2000 57.2000 ;
	    RECT 15.0000 56.8000 16.2000 57.1000 ;
	    RECT 16.6000 57.1000 17.0000 57.2000 ;
	    RECT 23.0000 57.1000 23.3000 57.8000 ;
	    RECT 86.2000 57.2000 86.5000 57.8000 ;
	    RECT 16.6000 56.8000 23.3000 57.1000 ;
	    RECT 27.0000 57.1000 27.4000 57.2000 ;
	    RECT 27.8000 57.1000 28.2000 57.2000 ;
	    RECT 27.0000 56.8000 28.2000 57.1000 ;
	    RECT 35.0000 56.8000 35.4000 57.2000 ;
	    RECT 38.2000 56.8000 38.6000 57.2000 ;
	    RECT 41.4000 56.8000 41.8000 57.2000 ;
	    RECT 70.2000 57.1000 70.6000 57.2000 ;
	    RECT 71.0000 57.1000 71.4000 57.2000 ;
	    RECT 70.2000 56.8000 71.4000 57.1000 ;
	    RECT 74.2000 57.1000 74.6000 57.2000 ;
	    RECT 75.0000 57.1000 75.4000 57.2000 ;
	    RECT 74.2000 56.8000 75.4000 57.1000 ;
	    RECT 86.2000 57.1000 86.6000 57.2000 ;
	    RECT 88.6000 57.1000 89.0000 57.2000 ;
	    RECT 95.8000 57.1000 96.2000 57.2000 ;
	    RECT 102.2000 57.1000 102.6000 57.2000 ;
	    RECT 86.2000 56.8000 102.6000 57.1000 ;
	    RECT 108.6000 57.1000 109.0000 57.2000 ;
	    RECT 109.4000 57.1000 109.8000 57.2000 ;
	    RECT 108.6000 56.8000 109.8000 57.1000 ;
	    RECT 117.4000 57.1000 117.8000 57.2000 ;
	    RECT 118.2000 57.1000 118.6000 57.2000 ;
	    RECT 117.4000 56.8000 118.6000 57.1000 ;
	    RECT 29.4000 55.8000 29.8000 56.2000 ;
	    RECT 35.0000 56.1000 35.3000 56.8000 ;
	    RECT 36.6000 56.1000 37.0000 56.2000 ;
	    RECT 35.0000 55.8000 37.0000 56.1000 ;
	    RECT 38.2000 56.1000 38.5000 56.8000 ;
	    RECT 40.6000 56.1000 41.0000 56.2000 ;
	    RECT 38.2000 55.8000 41.0000 56.1000 ;
	    RECT 41.4000 56.1000 41.7000 56.8000 ;
	    RECT 41.4000 55.8000 72.9000 56.1000 ;
	    RECT 3.0000 55.1000 3.4000 55.2000 ;
	    RECT 19.8000 55.1000 20.2000 55.2000 ;
	    RECT 23.0000 55.1000 23.4000 55.2000 ;
	    RECT 3.0000 54.8000 23.4000 55.1000 ;
	    RECT 24.6000 55.1000 25.0000 55.2000 ;
	    RECT 26.2000 55.1000 26.6000 55.2000 ;
	    RECT 24.6000 54.8000 26.6000 55.1000 ;
	    RECT 27.8000 55.1000 28.2000 55.2000 ;
	    RECT 29.4000 55.1000 29.7000 55.8000 ;
	    RECT 27.8000 54.8000 29.7000 55.1000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 39.0000 55.1000 39.4000 55.2000 ;
	    RECT 38.2000 54.8000 39.4000 55.1000 ;
	    RECT 41.4000 55.1000 41.8000 55.2000 ;
	    RECT 42.2000 55.1000 42.6000 55.2000 ;
	    RECT 41.4000 54.8000 42.6000 55.1000 ;
	    RECT 57.4000 55.1000 57.8000 55.2000 ;
	    RECT 58.2000 55.1000 58.6000 55.2000 ;
	    RECT 57.4000 54.8000 58.6000 55.1000 ;
	    RECT 63.8000 54.8000 64.2000 55.2000 ;
	    RECT 72.6000 55.1000 72.9000 55.8000 ;
	    RECT 83.0000 55.8000 83.4000 56.2000 ;
	    RECT 136.6000 56.1000 137.0000 56.2000 ;
	    RECT 137.4000 56.1000 137.8000 56.2000 ;
	    RECT 136.6000 55.8000 137.8000 56.1000 ;
	    RECT 140.6000 55.8000 141.0000 56.2000 ;
	    RECT 143.0000 56.1000 143.4000 56.2000 ;
	    RECT 149.4000 56.1000 149.8000 56.2000 ;
	    RECT 143.0000 55.8000 149.8000 56.1000 ;
	    RECT 155.0000 56.1000 155.4000 56.2000 ;
	    RECT 159.8000 56.1000 160.2000 56.2000 ;
	    RECT 155.0000 55.8000 160.9000 56.1000 ;
	    RECT 83.0000 55.1000 83.3000 55.8000 ;
	    RECT 72.6000 54.8000 83.3000 55.1000 ;
	    RECT 140.6000 55.1000 140.9000 55.8000 ;
	    RECT 146.2000 55.1000 146.6000 55.2000 ;
	    RECT 140.6000 54.8000 146.6000 55.1000 ;
	    RECT 163.0000 54.8000 163.4000 55.2000 ;
	    RECT 164.6000 55.1000 165.0000 55.2000 ;
	    RECT 165.4000 55.1000 165.8000 55.2000 ;
	    RECT 164.6000 54.8000 165.8000 55.1000 ;
	    RECT 63.8000 54.2000 64.1000 54.8000 ;
	    RECT 163.0000 54.2000 163.3000 54.8000 ;
	    RECT 2.2000 54.1000 2.6000 54.2000 ;
	    RECT 5.4000 54.1000 5.8000 54.2000 ;
	    RECT 2.2000 53.8000 5.8000 54.1000 ;
	    RECT 15.0000 54.1000 15.4000 54.2000 ;
	    RECT 17.4000 54.1000 17.8000 54.2000 ;
	    RECT 15.0000 53.8000 17.8000 54.1000 ;
	    RECT 18.2000 54.1000 18.6000 54.2000 ;
	    RECT 19.0000 54.1000 19.4000 54.2000 ;
	    RECT 18.2000 53.8000 19.4000 54.1000 ;
	    RECT 26.2000 54.1000 26.6000 54.2000 ;
	    RECT 39.0000 54.1000 39.4000 54.2000 ;
	    RECT 26.2000 53.8000 39.4000 54.1000 ;
	    RECT 40.6000 54.1000 41.0000 54.2000 ;
	    RECT 49.4000 54.1000 49.8000 54.2000 ;
	    RECT 40.6000 53.8000 49.8000 54.1000 ;
	    RECT 63.8000 53.8000 64.2000 54.2000 ;
	    RECT 70.2000 54.1000 70.6000 54.2000 ;
	    RECT 75.8000 54.1000 76.2000 54.2000 ;
	    RECT 70.2000 53.8000 76.2000 54.1000 ;
	    RECT 78.2000 54.1000 78.6000 54.2000 ;
	    RECT 79.0000 54.1000 79.4000 54.2000 ;
	    RECT 78.2000 53.8000 79.4000 54.1000 ;
	    RECT 108.6000 54.1000 109.0000 54.2000 ;
	    RECT 111.8000 54.1000 112.2000 54.2000 ;
	    RECT 108.6000 53.8000 112.2000 54.1000 ;
	    RECT 121.4000 54.1000 121.8000 54.2000 ;
	    RECT 123.0000 54.1000 123.4000 54.2000 ;
	    RECT 125.4000 54.1000 125.8000 54.2000 ;
	    RECT 128.6000 54.1000 129.0000 54.2000 ;
	    RECT 135.0000 54.1000 135.4000 54.2000 ;
	    RECT 121.4000 53.8000 135.4000 54.1000 ;
	    RECT 163.0000 53.8000 163.4000 54.2000 ;
	    RECT 168.6000 54.1000 169.0000 54.2000 ;
	    RECT 170.2000 54.1000 170.6000 54.2000 ;
	    RECT 168.6000 53.8000 170.6000 54.1000 ;
	    RECT 21.4000 53.1000 21.8000 53.2000 ;
	    RECT 32.6000 53.1000 33.0000 53.2000 ;
	    RECT 21.4000 52.8000 33.0000 53.1000 ;
	    RECT 35.8000 53.1000 36.2000 53.2000 ;
	    RECT 39.0000 53.1000 39.4000 53.2000 ;
	    RECT 41.4000 53.1000 41.8000 53.2000 ;
	    RECT 43.8000 53.1000 44.2000 53.2000 ;
	    RECT 35.8000 52.8000 44.2000 53.1000 ;
	    RECT 71.8000 53.1000 72.2000 53.2000 ;
	    RECT 72.6000 53.1000 73.0000 53.2000 ;
	    RECT 71.8000 52.8000 73.0000 53.1000 ;
	    RECT 143.8000 53.1000 144.2000 53.2000 ;
	    RECT 148.6000 53.1000 149.0000 53.2000 ;
	    RECT 143.8000 52.8000 149.0000 53.1000 ;
	    RECT 159.8000 53.1000 160.2000 53.2000 ;
	    RECT 169.4000 53.1000 169.8000 53.2000 ;
	    RECT 159.8000 52.8000 169.8000 53.1000 ;
	    RECT 15.0000 52.1000 15.4000 52.2000 ;
	    RECT 31.8000 52.1000 32.2000 52.2000 ;
	    RECT 15.0000 51.8000 32.2000 52.1000 ;
	    RECT 24.6000 51.1000 25.0000 51.2000 ;
	    RECT 33.4000 51.1000 33.8000 51.2000 ;
	    RECT 24.6000 50.8000 33.8000 51.1000 ;
	    RECT 116.6000 51.1000 117.0000 51.2000 ;
	    RECT 123.0000 51.1000 123.4000 51.2000 ;
	    RECT 116.6000 50.8000 123.4000 51.1000 ;
	    RECT 126.2000 51.1000 126.6000 51.2000 ;
	    RECT 127.0000 51.1000 127.4000 51.2000 ;
	    RECT 126.2000 50.8000 127.4000 51.1000 ;
	    RECT 9.4000 50.1000 9.8000 50.2000 ;
	    RECT 43.0000 50.1000 43.4000 50.2000 ;
	    RECT 9.4000 49.8000 43.4000 50.1000 ;
	    RECT 64.6000 50.1000 65.0000 50.2000 ;
	    RECT 79.0000 50.1000 79.4000 50.2000 ;
	    RECT 64.6000 49.8000 79.4000 50.1000 ;
	    RECT 118.2000 50.1000 118.6000 50.2000 ;
	    RECT 120.6000 50.1000 121.0000 50.2000 ;
	    RECT 118.2000 49.8000 121.0000 50.1000 ;
	    RECT 15.8000 49.1000 16.2000 49.2000 ;
	    RECT 27.8000 49.1000 28.2000 49.2000 ;
	    RECT 15.8000 48.8000 28.2000 49.1000 ;
	    RECT 171.0000 48.8000 171.4000 49.2000 ;
	    RECT 7.0000 48.1000 7.4000 48.2000 ;
	    RECT 10.2000 48.1000 10.6000 48.2000 ;
	    RECT 7.0000 47.8000 10.6000 48.1000 ;
	    RECT 19.8000 48.1000 20.2000 48.2000 ;
	    RECT 28.6000 48.1000 29.0000 48.2000 ;
	    RECT 19.8000 47.8000 29.0000 48.1000 ;
	    RECT 38.2000 48.1000 38.6000 48.2000 ;
	    RECT 41.4000 48.1000 41.8000 48.2000 ;
	    RECT 43.8000 48.1000 44.2000 48.2000 ;
	    RECT 38.2000 47.8000 44.2000 48.1000 ;
	    RECT 63.8000 47.8000 64.2000 48.2000 ;
	    RECT 72.6000 48.1000 73.0000 48.2000 ;
	    RECT 79.0000 48.1000 79.4000 48.2000 ;
	    RECT 72.6000 47.8000 79.4000 48.1000 ;
	    RECT 139.0000 48.1000 139.4000 48.2000 ;
	    RECT 146.2000 48.1000 146.6000 48.2000 ;
	    RECT 139.0000 47.8000 146.6000 48.1000 ;
	    RECT 169.4000 48.1000 169.8000 48.2000 ;
	    RECT 171.0000 48.1000 171.3000 48.8000 ;
	    RECT 169.4000 47.8000 171.3000 48.1000 ;
	    RECT 3.8000 46.8000 4.2000 47.2000 ;
	    RECT 23.0000 47.1000 23.4000 47.2000 ;
	    RECT 27.0000 47.1000 27.4000 47.2000 ;
	    RECT 38.2000 47.1000 38.6000 47.2000 ;
	    RECT 23.0000 46.8000 38.6000 47.1000 ;
	    RECT 40.6000 47.1000 41.0000 47.2000 ;
	    RECT 45.4000 47.1000 45.8000 47.2000 ;
	    RECT 40.6000 46.8000 45.8000 47.1000 ;
	    RECT 53.4000 47.1000 53.8000 47.2000 ;
	    RECT 61.4000 47.1000 61.8000 47.2000 ;
	    RECT 53.4000 46.8000 61.8000 47.1000 ;
	    RECT 63.8000 47.1000 64.1000 47.8000 ;
	    RECT 66.2000 47.1000 66.6000 47.2000 ;
	    RECT 63.8000 46.8000 66.6000 47.1000 ;
	    RECT 71.8000 47.1000 72.2000 47.2000 ;
	    RECT 75.0000 47.1000 75.4000 47.2000 ;
	    RECT 71.8000 46.8000 75.4000 47.1000 ;
	    RECT 77.4000 47.1000 77.8000 47.2000 ;
	    RECT 82.2000 47.1000 82.6000 47.2000 ;
	    RECT 89.4000 47.1000 89.8000 47.2000 ;
	    RECT 77.4000 46.8000 89.8000 47.1000 ;
	    RECT 91.0000 47.1000 91.4000 47.2000 ;
	    RECT 91.8000 47.1000 92.2000 47.2000 ;
	    RECT 91.0000 46.8000 92.2000 47.1000 ;
	    RECT 96.6000 47.1000 97.0000 47.2000 ;
	    RECT 102.2000 47.1000 102.6000 47.2000 ;
	    RECT 96.6000 46.8000 102.6000 47.1000 ;
	    RECT 119.0000 46.8000 119.4000 47.2000 ;
	    RECT 142.2000 47.1000 142.6000 47.2000 ;
	    RECT 140.6000 46.8000 142.6000 47.1000 ;
	    RECT 147.0000 47.1000 147.4000 47.2000 ;
	    RECT 147.8000 47.1000 148.2000 47.2000 ;
	    RECT 154.2000 47.1000 154.6000 47.2000 ;
	    RECT 147.0000 46.8000 154.6000 47.1000 ;
	    RECT 155.8000 46.8000 156.2000 47.2000 ;
	    RECT 158.2000 47.1000 158.6000 47.2000 ;
	    RECT 163.0000 47.1000 163.4000 47.2000 ;
	    RECT 158.2000 46.8000 163.4000 47.1000 ;
	    RECT 2.2000 46.1000 2.6000 46.2000 ;
	    RECT 3.8000 46.1000 4.1000 46.8000 ;
	    RECT 2.2000 45.8000 4.1000 46.1000 ;
	    RECT 10.2000 46.1000 10.6000 46.2000 ;
	    RECT 15.0000 46.1000 15.4000 46.2000 ;
	    RECT 10.2000 45.8000 15.4000 46.1000 ;
	    RECT 19.0000 46.1000 19.4000 46.2000 ;
	    RECT 21.4000 46.1000 21.8000 46.2000 ;
	    RECT 19.0000 45.8000 21.8000 46.1000 ;
	    RECT 28.6000 46.1000 29.0000 46.2000 ;
	    RECT 29.4000 46.1000 29.8000 46.2000 ;
	    RECT 28.6000 45.8000 29.8000 46.1000 ;
	    RECT 100.6000 46.1000 101.0000 46.2000 ;
	    RECT 101.4000 46.1000 101.8000 46.2000 ;
	    RECT 100.6000 45.8000 101.8000 46.1000 ;
	    RECT 104.6000 46.1000 105.0000 46.2000 ;
	    RECT 108.6000 46.1000 109.0000 46.2000 ;
	    RECT 112.6000 46.1000 113.0000 46.2000 ;
	    RECT 104.6000 45.8000 113.0000 46.1000 ;
	    RECT 117.4000 46.1000 117.8000 46.2000 ;
	    RECT 119.0000 46.1000 119.3000 46.8000 ;
	    RECT 140.6000 46.2000 140.9000 46.8000 ;
	    RECT 117.4000 45.8000 119.3000 46.1000 ;
	    RECT 123.8000 46.1000 124.2000 46.2000 ;
	    RECT 125.4000 46.1000 125.8000 46.2000 ;
	    RECT 123.8000 45.8000 125.8000 46.1000 ;
	    RECT 127.0000 46.1000 127.4000 46.2000 ;
	    RECT 130.2000 46.1000 130.6000 46.2000 ;
	    RECT 136.6000 46.1000 137.0000 46.2000 ;
	    RECT 127.0000 45.8000 128.1000 46.1000 ;
	    RECT 130.2000 45.8000 137.7000 46.1000 ;
	    RECT 140.6000 45.8000 141.0000 46.2000 ;
	    RECT 155.8000 46.1000 156.1000 46.8000 ;
	    RECT 157.4000 46.1000 157.8000 46.2000 ;
	    RECT 155.8000 45.8000 157.8000 46.1000 ;
	    RECT 166.2000 46.1000 166.6000 46.2000 ;
	    RECT 167.8000 46.1000 168.2000 46.2000 ;
	    RECT 166.2000 45.8000 168.2000 46.1000 ;
	    RECT 168.6000 45.8000 169.0000 46.2000 ;
	    RECT 15.0000 45.1000 15.4000 45.2000 ;
	    RECT 15.8000 45.1000 16.2000 45.2000 ;
	    RECT 15.0000 44.8000 16.2000 45.1000 ;
	    RECT 46.2000 45.1000 46.6000 45.2000 ;
	    RECT 47.0000 45.1000 47.4000 45.2000 ;
	    RECT 58.2000 45.1000 58.6000 45.2000 ;
	    RECT 46.2000 44.8000 47.4000 45.1000 ;
	    RECT 55.8000 44.8000 58.6000 45.1000 ;
	    RECT 60.6000 45.1000 61.0000 45.2000 ;
	    RECT 67.8000 45.1000 68.2000 45.2000 ;
	    RECT 60.6000 44.8000 68.2000 45.1000 ;
	    RECT 92.6000 45.1000 93.0000 45.2000 ;
	    RECT 93.4000 45.1000 93.8000 45.2000 ;
	    RECT 92.6000 44.8000 93.8000 45.1000 ;
	    RECT 108.6000 44.8000 109.0000 45.2000 ;
	    RECT 127.0000 44.8000 127.4000 45.2000 ;
	    RECT 127.8000 45.1000 128.1000 45.8000 ;
	    RECT 136.6000 45.1000 137.0000 45.2000 ;
	    RECT 137.4000 45.1000 137.8000 45.2000 ;
	    RECT 127.8000 44.8000 132.1000 45.1000 ;
	    RECT 136.6000 44.8000 137.8000 45.1000 ;
	    RECT 143.8000 45.1000 144.2000 45.2000 ;
	    RECT 144.6000 45.1000 145.0000 45.2000 ;
	    RECT 143.8000 44.8000 145.0000 45.1000 ;
	    RECT 149.4000 45.1000 149.8000 45.2000 ;
	    RECT 150.2000 45.1000 150.6000 45.2000 ;
	    RECT 149.4000 44.8000 150.6000 45.1000 ;
	    RECT 151.0000 45.1000 151.4000 45.2000 ;
	    RECT 163.8000 45.1000 164.2000 45.2000 ;
	    RECT 167.0000 45.1000 167.4000 45.2000 ;
	    RECT 168.6000 45.1000 168.9000 45.8000 ;
	    RECT 151.0000 44.8000 152.9000 45.1000 ;
	    RECT 163.8000 44.8000 165.7000 45.1000 ;
	    RECT 167.0000 44.8000 168.9000 45.1000 ;
	    RECT 55.8000 44.2000 56.1000 44.8000 ;
	    RECT 3.0000 44.1000 3.4000 44.2000 ;
	    RECT 7.8000 44.1000 8.2000 44.2000 ;
	    RECT 3.0000 43.8000 8.2000 44.1000 ;
	    RECT 11.8000 44.1000 12.2000 44.2000 ;
	    RECT 24.6000 44.1000 25.0000 44.2000 ;
	    RECT 11.8000 43.8000 25.0000 44.1000 ;
	    RECT 25.4000 43.8000 25.8000 44.2000 ;
	    RECT 31.8000 44.1000 32.2000 44.2000 ;
	    RECT 33.4000 44.1000 33.8000 44.2000 ;
	    RECT 31.8000 43.8000 33.8000 44.1000 ;
	    RECT 35.0000 44.1000 35.4000 44.2000 ;
	    RECT 44.6000 44.1000 45.0000 44.2000 ;
	    RECT 35.0000 43.8000 45.0000 44.1000 ;
	    RECT 51.8000 43.8000 52.2000 44.2000 ;
	    RECT 55.8000 43.8000 56.2000 44.2000 ;
	    RECT 59.0000 44.1000 59.4000 44.2000 ;
	    RECT 67.0000 44.1000 67.4000 44.2000 ;
	    RECT 59.0000 43.8000 67.4000 44.1000 ;
	    RECT 70.2000 44.1000 70.6000 44.2000 ;
	    RECT 84.6000 44.1000 85.0000 44.2000 ;
	    RECT 70.2000 43.8000 85.0000 44.1000 ;
	    RECT 86.2000 44.1000 86.6000 44.2000 ;
	    RECT 90.2000 44.1000 90.6000 44.2000 ;
	    RECT 86.2000 43.8000 90.6000 44.1000 ;
	    RECT 95.8000 44.1000 96.2000 44.2000 ;
	    RECT 97.4000 44.1000 97.8000 44.2000 ;
	    RECT 95.8000 43.8000 97.8000 44.1000 ;
	    RECT 102.2000 44.1000 102.6000 44.2000 ;
	    RECT 108.6000 44.1000 108.9000 44.8000 ;
	    RECT 127.0000 44.2000 127.3000 44.8000 ;
	    RECT 131.8000 44.2000 132.1000 44.8000 ;
	    RECT 102.2000 43.8000 108.9000 44.1000 ;
	    RECT 124.6000 44.1000 125.0000 44.2000 ;
	    RECT 126.2000 44.1000 126.6000 44.2000 ;
	    RECT 124.6000 43.8000 126.6000 44.1000 ;
	    RECT 127.0000 43.8000 127.4000 44.2000 ;
	    RECT 131.8000 43.8000 132.2000 44.2000 ;
	    RECT 152.6000 44.1000 152.9000 44.8000 ;
	    RECT 165.4000 44.2000 165.7000 44.8000 ;
	    RECT 162.2000 44.1000 162.6000 44.2000 ;
	    RECT 152.6000 43.8000 162.6000 44.1000 ;
	    RECT 165.4000 43.8000 165.8000 44.2000 ;
	    RECT 25.4000 43.2000 25.7000 43.8000 ;
	    RECT 18.2000 42.8000 18.6000 43.2000 ;
	    RECT 25.4000 42.8000 25.8000 43.2000 ;
	    RECT 51.8000 42.8000 52.1000 43.8000 ;
	    RECT 52.6000 43.1000 53.0000 43.2000 ;
	    RECT 57.4000 43.1000 57.8000 43.2000 ;
	    RECT 52.6000 42.8000 57.8000 43.1000 ;
	    RECT 61.4000 43.1000 61.8000 43.2000 ;
	    RECT 65.4000 43.1000 65.8000 43.2000 ;
	    RECT 61.4000 42.8000 65.8000 43.1000 ;
	    RECT 67.8000 43.1000 68.2000 43.2000 ;
	    RECT 71.0000 43.1000 71.4000 43.2000 ;
	    RECT 67.8000 42.8000 71.4000 43.1000 ;
	    RECT 74.2000 43.1000 74.6000 43.2000 ;
	    RECT 75.0000 43.1000 75.4000 43.2000 ;
	    RECT 74.2000 42.8000 75.4000 43.1000 ;
	    RECT 159.0000 43.1000 159.4000 43.2000 ;
	    RECT 164.6000 43.1000 165.0000 43.2000 ;
	    RECT 159.0000 42.8000 165.0000 43.1000 ;
	    RECT 4.6000 42.1000 5.0000 42.2000 ;
	    RECT 18.2000 42.1000 18.5000 42.8000 ;
	    RECT 4.6000 41.8000 18.5000 42.1000 ;
	    RECT 24.6000 42.1000 25.0000 42.2000 ;
	    RECT 117.4000 42.1000 117.8000 42.2000 ;
	    RECT 125.4000 42.1000 125.8000 42.2000 ;
	    RECT 24.6000 41.8000 30.5000 42.1000 ;
	    RECT 117.4000 41.8000 125.8000 42.1000 ;
	    RECT 126.2000 42.1000 126.6000 42.2000 ;
	    RECT 130.2000 42.1000 130.6000 42.2000 ;
	    RECT 126.2000 41.8000 130.6000 42.1000 ;
	    RECT 141.4000 42.1000 141.8000 42.2000 ;
	    RECT 144.6000 42.1000 145.0000 42.2000 ;
	    RECT 141.4000 41.8000 145.0000 42.1000 ;
	    RECT 148.6000 42.1000 149.0000 42.2000 ;
	    RECT 150.2000 42.1000 150.6000 42.2000 ;
	    RECT 148.6000 41.8000 150.6000 42.1000 ;
	    RECT 154.2000 42.1000 154.6000 42.2000 ;
	    RECT 156.6000 42.1000 157.0000 42.2000 ;
	    RECT 154.2000 41.8000 157.0000 42.1000 ;
	    RECT 30.2000 41.2000 30.5000 41.8000 ;
	    RECT 30.2000 40.8000 30.6000 41.2000 ;
	    RECT 67.0000 41.1000 67.4000 41.2000 ;
	    RECT 81.4000 41.1000 81.8000 41.2000 ;
	    RECT 67.0000 40.8000 81.8000 41.1000 ;
	    RECT 89.4000 41.1000 89.8000 41.2000 ;
	    RECT 95.0000 41.1000 95.4000 41.2000 ;
	    RECT 89.4000 40.8000 95.4000 41.1000 ;
	    RECT 106.2000 41.1000 106.6000 41.2000 ;
	    RECT 120.6000 41.1000 121.0000 41.2000 ;
	    RECT 106.2000 40.8000 121.0000 41.1000 ;
	    RECT 128.6000 41.1000 129.0000 41.2000 ;
	    RECT 144.6000 41.1000 145.0000 41.2000 ;
	    RECT 128.6000 40.8000 145.0000 41.1000 ;
	    RECT 147.8000 41.1000 148.2000 41.2000 ;
	    RECT 148.6000 41.1000 149.0000 41.2000 ;
	    RECT 147.8000 40.8000 149.0000 41.1000 ;
	    RECT 152.6000 41.1000 153.0000 41.2000 ;
	    RECT 163.8000 41.1000 164.2000 41.2000 ;
	    RECT 152.6000 40.8000 164.2000 41.1000 ;
	    RECT 15.0000 40.1000 15.4000 40.2000 ;
	    RECT 36.6000 40.1000 37.0000 40.2000 ;
	    RECT 15.0000 39.8000 37.0000 40.1000 ;
	    RECT 91.0000 40.1000 91.4000 40.2000 ;
	    RECT 104.6000 40.1000 105.0000 40.2000 ;
	    RECT 91.0000 39.8000 105.0000 40.1000 ;
	    RECT 110.2000 40.1000 110.6000 40.2000 ;
	    RECT 116.6000 40.1000 117.0000 40.2000 ;
	    RECT 110.2000 39.8000 117.0000 40.1000 ;
	    RECT 142.2000 40.1000 142.6000 40.2000 ;
	    RECT 147.8000 40.1000 148.2000 40.2000 ;
	    RECT 142.2000 39.8000 148.2000 40.1000 ;
	    RECT 162.2000 40.1000 162.6000 40.2000 ;
	    RECT 165.4000 40.1000 165.8000 40.2000 ;
	    RECT 162.2000 39.8000 165.8000 40.1000 ;
	    RECT 162.2000 39.1000 162.6000 39.2000 ;
	    RECT 163.0000 39.1000 163.4000 39.2000 ;
	    RECT 162.2000 38.8000 163.4000 39.1000 ;
	    RECT 17.4000 38.1000 17.8000 38.2000 ;
	    RECT 23.0000 38.1000 23.4000 38.2000 ;
	    RECT 17.4000 37.8000 23.4000 38.1000 ;
	    RECT 30.2000 38.1000 30.6000 38.2000 ;
	    RECT 39.8000 38.1000 40.2000 38.2000 ;
	    RECT 30.2000 37.8000 40.2000 38.1000 ;
	    RECT 49.4000 38.1000 49.8000 38.2000 ;
	    RECT 51.0000 38.1000 51.4000 38.2000 ;
	    RECT 59.0000 38.1000 59.4000 38.2000 ;
	    RECT 49.4000 37.8000 59.4000 38.1000 ;
	    RECT 65.4000 38.1000 65.8000 38.2000 ;
	    RECT 68.6000 38.1000 69.0000 38.2000 ;
	    RECT 72.6000 38.1000 73.0000 38.2000 ;
	    RECT 86.2000 38.1000 86.6000 38.2000 ;
	    RECT 97.4000 38.1000 97.8000 38.2000 ;
	    RECT 65.4000 37.8000 69.0000 38.1000 ;
	    RECT 71.8000 37.8000 73.0000 38.1000 ;
	    RECT 85.4000 37.8000 97.8000 38.1000 ;
	    RECT 98.2000 38.1000 98.6000 38.2000 ;
	    RECT 109.4000 38.1000 109.8000 38.2000 ;
	    RECT 119.8000 38.1000 120.2000 38.2000 ;
	    RECT 124.6000 38.1000 125.0000 38.2000 ;
	    RECT 98.2000 37.8000 125.0000 38.1000 ;
	    RECT 1.4000 37.1000 1.8000 37.2000 ;
	    RECT 2.2000 37.1000 2.6000 37.2000 ;
	    RECT 1.4000 36.8000 2.6000 37.1000 ;
	    RECT 133.4000 37.1000 133.8000 37.2000 ;
	    RECT 139.8000 37.1000 140.2000 37.2000 ;
	    RECT 133.4000 36.8000 140.2000 37.1000 ;
	    RECT 141.4000 37.1000 141.8000 37.2000 ;
	    RECT 142.2000 37.1000 142.6000 37.2000 ;
	    RECT 148.6000 37.1000 149.0000 37.2000 ;
	    RECT 156.6000 37.1000 157.0000 37.2000 ;
	    RECT 161.4000 37.1000 161.8000 37.2000 ;
	    RECT 141.4000 36.8000 142.6000 37.1000 ;
	    RECT 147.8000 36.8000 149.0000 37.1000 ;
	    RECT 155.8000 36.8000 161.8000 37.1000 ;
	    RECT 5.4000 36.1000 5.8000 36.2000 ;
	    RECT 16.6000 36.1000 17.0000 36.2000 ;
	    RECT 17.4000 36.1000 17.8000 36.2000 ;
	    RECT 5.4000 35.8000 17.8000 36.1000 ;
	    RECT 18.2000 36.1000 18.6000 36.2000 ;
	    RECT 19.8000 36.1000 20.2000 36.2000 ;
	    RECT 18.2000 35.8000 20.2000 36.1000 ;
	    RECT 21.4000 35.8000 21.8000 36.2000 ;
	    RECT 23.0000 36.1000 23.4000 36.2000 ;
	    RECT 28.6000 36.1000 29.0000 36.2000 ;
	    RECT 23.0000 35.8000 29.0000 36.1000 ;
	    RECT 31.8000 35.8000 32.2000 36.2000 ;
	    RECT 39.8000 36.1000 40.2000 36.2000 ;
	    RECT 42.2000 36.1000 42.6000 36.2000 ;
	    RECT 39.8000 35.8000 42.6000 36.1000 ;
	    RECT 43.8000 36.1000 44.2000 36.2000 ;
	    RECT 53.4000 36.1000 53.8000 36.2000 ;
	    RECT 43.8000 35.8000 53.8000 36.1000 ;
	    RECT 55.8000 36.1000 56.2000 36.2000 ;
	    RECT 63.0000 36.1000 63.4000 36.2000 ;
	    RECT 64.6000 36.1000 65.0000 36.2000 ;
	    RECT 55.8000 35.8000 65.0000 36.1000 ;
	    RECT 66.2000 36.1000 66.6000 36.2000 ;
	    RECT 70.2000 36.1000 70.6000 36.2000 ;
	    RECT 66.2000 35.8000 70.6000 36.1000 ;
	    RECT 76.6000 36.1000 77.0000 36.2000 ;
	    RECT 82.2000 36.1000 82.6000 36.2000 ;
	    RECT 76.6000 35.8000 82.6000 36.1000 ;
	    RECT 88.6000 36.1000 89.0000 36.2000 ;
	    RECT 89.4000 36.1000 89.8000 36.2000 ;
	    RECT 88.6000 35.8000 89.8000 36.1000 ;
	    RECT 93.4000 35.8000 93.8000 36.2000 ;
	    RECT 97.4000 36.1000 97.8000 36.2000 ;
	    RECT 99.8000 36.1000 100.2000 36.2000 ;
	    RECT 97.4000 35.8000 100.2000 36.1000 ;
	    RECT 100.6000 35.8000 101.0000 36.2000 ;
	    RECT 102.2000 36.1000 102.6000 36.2000 ;
	    RECT 104.6000 36.1000 105.0000 36.2000 ;
	    RECT 102.2000 35.8000 105.0000 36.1000 ;
	    RECT 114.2000 36.1000 114.6000 36.2000 ;
	    RECT 118.2000 36.1000 118.6000 36.2000 ;
	    RECT 127.8000 36.1000 128.2000 36.2000 ;
	    RECT 114.2000 35.8000 128.2000 36.1000 ;
	    RECT 163.0000 36.1000 163.4000 36.2000 ;
	    RECT 163.8000 36.1000 164.2000 36.2000 ;
	    RECT 163.0000 35.8000 164.2000 36.1000 ;
	    RECT 166.2000 36.1000 166.6000 36.2000 ;
	    RECT 170.2000 36.1000 170.6000 36.2000 ;
	    RECT 166.2000 35.8000 170.6000 36.1000 ;
	    RECT 21.4000 35.2000 21.7000 35.8000 ;
	    RECT 4.6000 35.1000 5.0000 35.2000 ;
	    RECT 7.0000 35.1000 7.4000 35.2000 ;
	    RECT 4.6000 34.8000 7.4000 35.1000 ;
	    RECT 11.0000 34.8000 11.4000 35.2000 ;
	    RECT 12.6000 35.1000 13.0000 35.2000 ;
	    RECT 18.2000 35.1000 18.6000 35.2000 ;
	    RECT 12.6000 34.8000 18.6000 35.1000 ;
	    RECT 21.4000 34.8000 21.8000 35.2000 ;
	    RECT 23.0000 35.1000 23.4000 35.2000 ;
	    RECT 23.8000 35.1000 24.2000 35.2000 ;
	    RECT 28.6000 35.1000 29.0000 35.2000 ;
	    RECT 23.0000 34.8000 24.2000 35.1000 ;
	    RECT 25.4000 34.8000 29.0000 35.1000 ;
	    RECT 30.2000 35.1000 30.6000 35.2000 ;
	    RECT 31.8000 35.1000 32.1000 35.8000 ;
	    RECT 47.8000 35.1000 48.2000 35.2000 ;
	    RECT 30.2000 34.8000 32.1000 35.1000 ;
	    RECT 46.2000 34.8000 48.2000 35.1000 ;
	    RECT 56.6000 35.1000 57.0000 35.2000 ;
	    RECT 58.2000 35.1000 58.6000 35.2000 ;
	    RECT 56.6000 34.8000 58.6000 35.1000 ;
	    RECT 75.8000 35.1000 76.2000 35.2000 ;
	    RECT 76.6000 35.1000 77.0000 35.2000 ;
	    RECT 75.8000 34.8000 77.0000 35.1000 ;
	    RECT 78.2000 35.1000 78.6000 35.2000 ;
	    RECT 82.2000 35.1000 82.6000 35.2000 ;
	    RECT 78.2000 34.8000 82.6000 35.1000 ;
	    RECT 93.4000 35.1000 93.7000 35.8000 ;
	    RECT 95.0000 35.1000 95.4000 35.2000 ;
	    RECT 100.6000 35.1000 100.9000 35.8000 ;
	    RECT 93.4000 34.8000 95.4000 35.1000 ;
	    RECT 99.0000 34.8000 100.9000 35.1000 ;
	    RECT 104.6000 35.1000 105.0000 35.2000 ;
	    RECT 134.2000 35.1000 134.6000 35.2000 ;
	    RECT 104.6000 34.8000 134.6000 35.1000 ;
	    RECT 139.0000 35.1000 139.4000 35.2000 ;
	    RECT 141.4000 35.1000 141.8000 35.2000 ;
	    RECT 139.0000 34.8000 141.8000 35.1000 ;
	    RECT 145.4000 35.1000 145.8000 35.2000 ;
	    RECT 150.2000 35.1000 150.6000 35.2000 ;
	    RECT 151.0000 35.1000 151.4000 35.2000 ;
	    RECT 162.2000 35.1000 162.6000 35.2000 ;
	    RECT 163.0000 35.1000 163.4000 35.2000 ;
	    RECT 145.4000 34.8000 152.1000 35.1000 ;
	    RECT 162.2000 34.8000 163.4000 35.1000 ;
	    RECT 166.2000 35.1000 166.6000 35.2000 ;
	    RECT 171.8000 35.1000 172.2000 35.2000 ;
	    RECT 166.2000 34.8000 172.2000 35.1000 ;
	    RECT 11.0000 34.2000 11.3000 34.8000 ;
	    RECT 25.4000 34.2000 25.7000 34.8000 ;
	    RECT 46.2000 34.2000 46.5000 34.8000 ;
	    RECT 99.0000 34.2000 99.3000 34.8000 ;
	    RECT 0.6000 34.1000 1.0000 34.2000 ;
	    RECT 5.4000 34.1000 5.8000 34.2000 ;
	    RECT 0.6000 33.8000 5.8000 34.1000 ;
	    RECT 11.0000 33.8000 11.4000 34.2000 ;
	    RECT 25.4000 33.8000 25.8000 34.2000 ;
	    RECT 26.2000 34.1000 26.6000 34.2000 ;
	    RECT 39.0000 34.1000 39.4000 34.2000 ;
	    RECT 26.2000 33.8000 39.4000 34.1000 ;
	    RECT 46.2000 33.8000 46.6000 34.2000 ;
	    RECT 48.6000 34.1000 49.0000 34.2000 ;
	    RECT 55.8000 34.1000 56.2000 34.2000 ;
	    RECT 48.6000 33.8000 56.2000 34.1000 ;
	    RECT 57.4000 34.1000 57.8000 34.2000 ;
	    RECT 58.2000 34.1000 58.6000 34.2000 ;
	    RECT 57.4000 33.8000 58.6000 34.1000 ;
	    RECT 64.6000 34.1000 65.0000 34.2000 ;
	    RECT 65.4000 34.1000 65.8000 34.2000 ;
	    RECT 64.6000 33.8000 65.8000 34.1000 ;
	    RECT 73.4000 34.1000 73.8000 34.2000 ;
	    RECT 76.6000 34.1000 77.0000 34.2000 ;
	    RECT 73.4000 33.8000 77.0000 34.1000 ;
	    RECT 87.0000 34.1000 87.4000 34.2000 ;
	    RECT 89.4000 34.1000 89.8000 34.2000 ;
	    RECT 91.0000 34.1000 91.4000 34.2000 ;
	    RECT 87.0000 33.8000 91.4000 34.1000 ;
	    RECT 97.4000 34.1000 97.8000 34.2000 ;
	    RECT 97.4000 33.8000 98.5000 34.1000 ;
	    RECT 99.0000 33.8000 99.4000 34.2000 ;
	    RECT 104.6000 34.1000 105.0000 34.2000 ;
	    RECT 109.4000 34.1000 109.8000 34.2000 ;
	    RECT 116.6000 34.1000 117.0000 34.2000 ;
	    RECT 118.2000 34.1000 118.6000 34.2000 ;
	    RECT 104.6000 33.8000 109.8000 34.1000 ;
	    RECT 115.8000 33.8000 118.6000 34.1000 ;
	    RECT 119.0000 34.1000 119.4000 34.2000 ;
	    RECT 120.6000 34.1000 121.0000 34.2000 ;
	    RECT 119.0000 33.8000 121.0000 34.1000 ;
	    RECT 125.4000 33.8000 125.8000 34.2000 ;
	    RECT 132.6000 34.1000 133.0000 34.2000 ;
	    RECT 143.0000 34.1000 143.4000 34.2000 ;
	    RECT 132.6000 33.8000 143.4000 34.1000 ;
	    RECT 143.8000 34.1000 144.2000 34.2000 ;
	    RECT 154.2000 34.1000 154.6000 34.2000 ;
	    RECT 143.8000 33.8000 154.6000 34.1000 ;
	    RECT 159.0000 34.1000 159.4000 34.2000 ;
	    RECT 161.4000 34.1000 161.8000 34.2000 ;
	    RECT 159.0000 33.8000 161.8000 34.1000 ;
	    RECT 125.4000 33.2000 125.7000 33.8000 ;
	    RECT 1.4000 33.1000 1.8000 33.2000 ;
	    RECT 3.0000 33.1000 3.4000 33.2000 ;
	    RECT 22.2000 33.1000 22.6000 33.2000 ;
	    RECT 1.4000 32.8000 22.6000 33.1000 ;
	    RECT 24.6000 33.1000 25.0000 33.2000 ;
	    RECT 36.6000 33.1000 37.0000 33.2000 ;
	    RECT 24.6000 32.8000 37.0000 33.1000 ;
	    RECT 55.0000 33.1000 55.4000 33.2000 ;
	    RECT 58.2000 33.1000 58.6000 33.2000 ;
	    RECT 55.0000 32.8000 58.6000 33.1000 ;
	    RECT 67.8000 33.1000 68.2000 33.2000 ;
	    RECT 75.0000 33.1000 75.4000 33.2000 ;
	    RECT 67.8000 32.8000 75.4000 33.1000 ;
	    RECT 125.4000 32.8000 125.8000 33.2000 ;
	    RECT 137.4000 33.1000 137.8000 33.2000 ;
	    RECT 146.2000 33.1000 146.6000 33.2000 ;
	    RECT 137.4000 32.8000 146.6000 33.1000 ;
	    RECT 2.2000 32.1000 2.6000 32.2000 ;
	    RECT 4.6000 32.1000 5.0000 32.2000 ;
	    RECT 2.2000 31.8000 5.0000 32.1000 ;
	    RECT 21.4000 32.1000 21.8000 32.2000 ;
	    RECT 27.0000 32.1000 27.4000 32.2000 ;
	    RECT 21.4000 31.8000 27.4000 32.1000 ;
	    RECT 53.4000 32.1000 53.8000 32.2000 ;
	    RECT 59.0000 32.1000 59.4000 32.2000 ;
	    RECT 53.4000 31.8000 59.4000 32.1000 ;
	    RECT 74.2000 32.1000 74.6000 32.2000 ;
	    RECT 91.0000 32.1000 91.4000 32.2000 ;
	    RECT 74.2000 31.8000 91.4000 32.1000 ;
	    RECT 136.6000 32.1000 137.0000 32.2000 ;
	    RECT 142.2000 32.1000 142.6000 32.2000 ;
	    RECT 136.6000 31.8000 142.6000 32.1000 ;
	    RECT 144.6000 32.1000 145.0000 32.2000 ;
	    RECT 147.0000 32.1000 147.4000 32.2000 ;
	    RECT 144.6000 31.8000 147.4000 32.1000 ;
	    RECT 147.8000 32.1000 148.2000 32.2000 ;
	    RECT 149.4000 32.1000 149.8000 32.2000 ;
	    RECT 147.8000 31.8000 149.8000 32.1000 ;
	    RECT 150.2000 32.1000 150.6000 32.2000 ;
	    RECT 151.8000 32.1000 152.2000 32.2000 ;
	    RECT 150.2000 31.8000 152.2000 32.1000 ;
	    RECT 1.4000 31.1000 1.8000 31.2000 ;
	    RECT 2.2000 31.1000 2.6000 31.2000 ;
	    RECT 1.4000 30.8000 2.6000 31.1000 ;
	    RECT 98.2000 31.1000 98.6000 31.2000 ;
	    RECT 109.4000 31.1000 109.8000 31.2000 ;
	    RECT 98.2000 30.8000 109.8000 31.1000 ;
	    RECT 116.6000 31.1000 117.0000 31.2000 ;
	    RECT 117.4000 31.1000 117.8000 31.2000 ;
	    RECT 116.6000 30.8000 117.8000 31.1000 ;
	    RECT 105.4000 30.1000 105.8000 30.2000 ;
	    RECT 110.2000 30.1000 110.6000 30.2000 ;
	    RECT 105.4000 29.8000 110.6000 30.1000 ;
	    RECT 117.4000 30.1000 117.8000 30.2000 ;
	    RECT 121.4000 30.1000 121.8000 30.2000 ;
	    RECT 117.4000 29.8000 121.8000 30.1000 ;
	    RECT 127.8000 30.1000 128.2000 30.2000 ;
	    RECT 129.4000 30.1000 129.8000 30.2000 ;
	    RECT 135.8000 30.1000 136.2000 30.2000 ;
	    RECT 139.8000 30.1000 140.2000 30.2000 ;
	    RECT 159.0000 30.1000 159.4000 30.2000 ;
	    RECT 127.8000 29.8000 159.4000 30.1000 ;
	    RECT 11.0000 28.8000 11.4000 29.2000 ;
	    RECT 30.2000 29.1000 30.6000 29.2000 ;
	    RECT 34.2000 29.1000 34.6000 29.2000 ;
	    RECT 39.0000 29.1000 39.4000 29.2000 ;
	    RECT 40.6000 29.1000 41.0000 29.2000 ;
	    RECT 30.2000 28.8000 41.0000 29.1000 ;
	    RECT 67.8000 29.1000 68.2000 29.2000 ;
	    RECT 75.8000 29.1000 76.2000 29.2000 ;
	    RECT 67.8000 28.8000 76.2000 29.1000 ;
	    RECT 95.8000 29.1000 96.2000 29.2000 ;
	    RECT 99.8000 29.1000 100.2000 29.2000 ;
	    RECT 111.0000 29.1000 111.4000 29.2000 ;
	    RECT 114.2000 29.1000 114.6000 29.2000 ;
	    RECT 95.8000 28.8000 114.6000 29.1000 ;
	    RECT 156.6000 28.8000 157.0000 29.2000 ;
	    RECT 168.6000 29.1000 169.0000 29.2000 ;
	    RECT 169.4000 29.1000 169.8000 29.2000 ;
	    RECT 168.6000 28.8000 169.8000 29.1000 ;
	    RECT 3.8000 28.1000 4.2000 28.2000 ;
	    RECT 6.2000 28.1000 6.6000 28.2000 ;
	    RECT 11.0000 28.1000 11.3000 28.8000 ;
	    RECT 3.8000 27.8000 11.3000 28.1000 ;
	    RECT 28.6000 28.1000 29.0000 28.2000 ;
	    RECT 30.2000 28.1000 30.5000 28.8000 ;
	    RECT 28.6000 27.8000 30.5000 28.1000 ;
	    RECT 32.6000 28.1000 33.0000 28.2000 ;
	    RECT 50.2000 28.1000 50.6000 28.2000 ;
	    RECT 63.8000 28.1000 64.2000 28.2000 ;
	    RECT 67.8000 28.1000 68.1000 28.8000 ;
	    RECT 69.4000 28.1000 69.8000 28.2000 ;
	    RECT 32.6000 27.8000 40.1000 28.1000 ;
	    RECT 50.2000 27.8000 69.8000 28.1000 ;
	    RECT 73.4000 28.1000 73.8000 28.2000 ;
	    RECT 81.4000 28.1000 81.8000 28.2000 ;
	    RECT 73.4000 27.8000 81.8000 28.1000 ;
	    RECT 85.4000 28.1000 85.8000 28.2000 ;
	    RECT 89.4000 28.1000 89.8000 28.2000 ;
	    RECT 110.2000 28.1000 110.6000 28.2000 ;
	    RECT 85.4000 27.8000 110.6000 28.1000 ;
	    RECT 115.8000 28.1000 116.2000 28.2000 ;
	    RECT 119.8000 28.1000 120.2000 28.2000 ;
	    RECT 127.8000 28.1000 128.2000 28.2000 ;
	    RECT 115.8000 27.8000 128.2000 28.1000 ;
	    RECT 156.6000 28.1000 156.9000 28.8000 ;
	    RECT 159.8000 28.1000 160.2000 28.2000 ;
	    RECT 167.8000 28.1000 168.2000 28.2000 ;
	    RECT 171.0000 28.1000 171.4000 28.2000 ;
	    RECT 156.6000 27.8000 171.4000 28.1000 ;
	    RECT 39.8000 27.2000 40.1000 27.8000 ;
	    RECT 11.0000 26.8000 11.4000 27.2000 ;
	    RECT 23.0000 27.1000 23.4000 27.2000 ;
	    RECT 26.2000 27.1000 26.6000 27.2000 ;
	    RECT 23.0000 26.8000 26.6000 27.1000 ;
	    RECT 36.6000 26.8000 37.0000 27.2000 ;
	    RECT 39.8000 26.8000 40.2000 27.2000 ;
	    RECT 88.6000 26.8000 89.0000 27.2000 ;
	    RECT 95.0000 27.1000 95.4000 27.2000 ;
	    RECT 98.2000 27.1000 98.6000 27.2000 ;
	    RECT 95.0000 26.8000 98.6000 27.1000 ;
	    RECT 100.6000 27.1000 101.0000 27.2000 ;
	    RECT 101.4000 27.1000 101.8000 27.2000 ;
	    RECT 100.6000 26.8000 101.8000 27.1000 ;
	    RECT 107.0000 27.1000 107.4000 27.2000 ;
	    RECT 108.6000 27.1000 109.0000 27.2000 ;
	    RECT 110.2000 27.1000 110.5000 27.8000 ;
	    RECT 107.0000 26.8000 110.5000 27.1000 ;
	    RECT 130.2000 26.8000 130.6000 27.2000 ;
	    RECT 142.2000 26.8000 142.6000 27.2000 ;
	    RECT 11.0000 26.2000 11.3000 26.8000 ;
	    RECT 11.0000 25.8000 11.4000 26.2000 ;
	    RECT 35.0000 26.1000 35.4000 26.2000 ;
	    RECT 36.6000 26.1000 36.9000 26.8000 ;
	    RECT 52.6000 26.1000 53.0000 26.2000 ;
	    RECT 53.4000 26.1000 53.8000 26.2000 ;
	    RECT 35.0000 25.8000 36.9000 26.1000 ;
	    RECT 51.8000 25.8000 53.8000 26.1000 ;
	    RECT 55.0000 26.1000 55.4000 26.2000 ;
	    RECT 56.6000 26.1000 57.0000 26.2000 ;
	    RECT 55.0000 25.8000 57.0000 26.1000 ;
	    RECT 87.0000 25.8000 87.4000 26.2000 ;
	    RECT 88.6000 26.1000 88.9000 26.8000 ;
	    RECT 122.2000 26.1000 122.6000 26.2000 ;
	    RECT 123.0000 26.1000 123.4000 26.2000 ;
	    RECT 88.6000 25.8000 112.1000 26.1000 ;
	    RECT 121.4000 25.8000 123.4000 26.1000 ;
	    RECT 125.4000 25.8000 125.8000 26.2000 ;
	    RECT 130.2000 26.1000 130.5000 26.8000 ;
	    RECT 131.8000 26.1000 132.2000 26.2000 ;
	    RECT 130.2000 25.8000 132.2000 26.1000 ;
	    RECT 142.2000 26.1000 142.5000 26.8000 ;
	    RECT 143.8000 26.1000 144.2000 26.2000 ;
	    RECT 142.2000 25.8000 144.2000 26.1000 ;
	    RECT 163.0000 26.1000 163.4000 26.2000 ;
	    RECT 171.8000 26.1000 172.2000 26.2000 ;
	    RECT 163.0000 25.8000 172.2000 26.1000 ;
	    RECT 22.2000 25.1000 22.6000 25.2000 ;
	    RECT 26.2000 25.1000 26.6000 25.2000 ;
	    RECT 31.8000 25.1000 32.2000 25.2000 ;
	    RECT 34.2000 25.1000 34.6000 25.2000 ;
	    RECT 22.2000 24.8000 34.6000 25.1000 ;
	    RECT 45.4000 25.1000 45.8000 25.2000 ;
	    RECT 53.4000 25.1000 53.8000 25.2000 ;
	    RECT 45.4000 24.8000 53.8000 25.1000 ;
	    RECT 57.4000 25.1000 57.8000 25.2000 ;
	    RECT 60.6000 25.1000 61.0000 25.2000 ;
	    RECT 57.4000 24.8000 61.0000 25.1000 ;
	    RECT 64.6000 25.1000 65.0000 25.2000 ;
	    RECT 67.0000 25.1000 67.4000 25.2000 ;
	    RECT 64.6000 24.8000 67.4000 25.1000 ;
	    RECT 87.0000 25.1000 87.3000 25.8000 ;
	    RECT 95.0000 25.1000 95.4000 25.2000 ;
	    RECT 87.0000 24.8000 95.4000 25.1000 ;
	    RECT 111.8000 25.1000 112.1000 25.8000 ;
	    RECT 125.4000 25.2000 125.7000 25.8000 ;
	    RECT 115.0000 25.1000 115.4000 25.2000 ;
	    RECT 111.8000 24.8000 115.4000 25.1000 ;
	    RECT 115.8000 25.1000 116.2000 25.2000 ;
	    RECT 123.0000 25.1000 123.4000 25.2000 ;
	    RECT 115.8000 24.8000 123.4000 25.1000 ;
	    RECT 125.4000 24.8000 125.8000 25.2000 ;
	    RECT 132.6000 25.1000 133.0000 25.2000 ;
	    RECT 135.0000 25.1000 135.4000 25.2000 ;
	    RECT 132.6000 24.8000 135.4000 25.1000 ;
	    RECT 135.8000 25.1000 136.2000 25.2000 ;
	    RECT 147.8000 25.1000 148.2000 25.2000 ;
	    RECT 151.0000 25.1000 151.4000 25.2000 ;
	    RECT 135.8000 24.8000 148.2000 25.1000 ;
	    RECT 150.2000 24.8000 151.4000 25.1000 ;
	    RECT 151.8000 25.1000 152.2000 25.2000 ;
	    RECT 162.2000 25.1000 162.6000 25.2000 ;
	    RECT 151.8000 24.8000 162.6000 25.1000 ;
	    RECT 150.2000 24.2000 150.5000 24.8000 ;
	    RECT 7.0000 24.1000 7.4000 24.2000 ;
	    RECT 7.8000 24.1000 8.2000 24.2000 ;
	    RECT 7.0000 23.8000 8.2000 24.1000 ;
	    RECT 14.2000 24.1000 14.6000 24.2000 ;
	    RECT 15.0000 24.1000 15.4000 24.2000 ;
	    RECT 14.2000 23.8000 15.4000 24.1000 ;
	    RECT 19.8000 24.1000 20.2000 24.2000 ;
	    RECT 25.4000 24.1000 25.8000 24.2000 ;
	    RECT 19.8000 23.8000 25.8000 24.1000 ;
	    RECT 26.2000 24.1000 26.6000 24.2000 ;
	    RECT 31.0000 24.1000 31.4000 24.2000 ;
	    RECT 26.2000 23.8000 31.4000 24.1000 ;
	    RECT 123.8000 24.1000 124.2000 24.2000 ;
	    RECT 135.0000 24.1000 135.4000 24.2000 ;
	    RECT 123.8000 23.8000 135.4000 24.1000 ;
	    RECT 139.0000 24.1000 139.4000 24.2000 ;
	    RECT 140.6000 24.1000 141.0000 24.2000 ;
	    RECT 139.0000 23.8000 141.0000 24.1000 ;
	    RECT 150.2000 23.8000 150.6000 24.2000 ;
	    RECT 153.4000 24.1000 153.8000 24.2000 ;
	    RECT 159.0000 24.1000 159.4000 24.2000 ;
	    RECT 153.4000 23.8000 159.4000 24.1000 ;
	    RECT 9.4000 23.1000 9.8000 23.2000 ;
	    RECT 23.8000 23.1000 24.2000 23.2000 ;
	    RECT 9.4000 22.8000 24.2000 23.1000 ;
	    RECT 24.6000 23.1000 25.0000 23.2000 ;
	    RECT 34.2000 23.1000 34.6000 23.2000 ;
	    RECT 24.6000 22.8000 34.6000 23.1000 ;
	    RECT 54.2000 23.1000 54.6000 23.2000 ;
	    RECT 56.6000 23.1000 57.0000 23.2000 ;
	    RECT 54.2000 22.8000 57.0000 23.1000 ;
	    RECT 17.4000 22.1000 17.8000 22.2000 ;
	    RECT 27.0000 22.1000 27.4000 22.2000 ;
	    RECT 17.4000 21.8000 27.4000 22.1000 ;
	    RECT 49.4000 22.1000 49.8000 22.2000 ;
	    RECT 55.0000 22.1000 55.4000 22.2000 ;
	    RECT 49.4000 21.8000 55.4000 22.1000 ;
	    RECT 75.0000 22.1000 75.4000 22.2000 ;
	    RECT 76.6000 22.1000 77.0000 22.2000 ;
	    RECT 75.0000 21.8000 77.0000 22.1000 ;
	    RECT 83.0000 22.1000 83.4000 22.2000 ;
	    RECT 85.4000 22.1000 85.8000 22.2000 ;
	    RECT 91.0000 22.1000 91.4000 22.2000 ;
	    RECT 94.2000 22.1000 94.6000 22.2000 ;
	    RECT 83.0000 21.8000 85.8000 22.1000 ;
	    RECT 90.2000 21.8000 94.6000 22.1000 ;
	    RECT 100.6000 22.1000 101.0000 22.2000 ;
	    RECT 107.8000 22.1000 108.2000 22.2000 ;
	    RECT 100.6000 21.8000 108.2000 22.1000 ;
	    RECT 108.6000 22.1000 109.0000 22.2000 ;
	    RECT 111.8000 22.1000 112.2000 22.2000 ;
	    RECT 108.6000 21.8000 112.2000 22.1000 ;
	    RECT 115.8000 22.1000 116.2000 22.2000 ;
	    RECT 116.6000 22.1000 117.0000 22.2000 ;
	    RECT 115.8000 21.8000 117.0000 22.1000 ;
	    RECT 18.2000 21.1000 18.6000 21.2000 ;
	    RECT 23.8000 21.1000 24.2000 21.2000 ;
	    RECT 18.2000 20.8000 24.2000 21.1000 ;
	    RECT 69.4000 21.1000 69.8000 21.2000 ;
	    RECT 73.4000 21.1000 73.8000 21.2000 ;
	    RECT 69.4000 20.8000 73.8000 21.1000 ;
	    RECT 111.0000 21.1000 111.4000 21.2000 ;
	    RECT 124.6000 21.1000 125.0000 21.2000 ;
	    RECT 111.0000 20.8000 125.0000 21.1000 ;
	    RECT 133.4000 21.1000 133.8000 21.2000 ;
	    RECT 147.0000 21.1000 147.4000 21.2000 ;
	    RECT 149.4000 21.1000 149.8000 21.2000 ;
	    RECT 161.4000 21.1000 161.8000 21.2000 ;
	    RECT 164.6000 21.1000 165.0000 21.2000 ;
	    RECT 133.4000 20.8000 165.0000 21.1000 ;
	    RECT 155.8000 20.1000 156.2000 20.2000 ;
	    RECT 165.4000 20.1000 165.8000 20.2000 ;
	    RECT 155.8000 19.8000 165.8000 20.1000 ;
	    RECT 1.4000 19.1000 1.8000 19.2000 ;
	    RECT 5.4000 19.1000 5.8000 19.2000 ;
	    RECT 1.4000 18.8000 5.8000 19.1000 ;
	    RECT 18.2000 19.1000 18.6000 19.2000 ;
	    RECT 109.4000 19.1000 109.8000 19.2000 ;
	    RECT 123.0000 19.1000 123.4000 19.2000 ;
	    RECT 18.2000 18.8000 32.9000 19.1000 ;
	    RECT 109.4000 18.8000 123.4000 19.1000 ;
	    RECT 131.0000 18.8000 131.4000 19.2000 ;
	    RECT 32.6000 18.2000 32.9000 18.8000 ;
	    RECT 21.4000 17.8000 21.8000 18.2000 ;
	    RECT 32.6000 17.8000 33.0000 18.2000 ;
	    RECT 106.2000 18.1000 106.6000 18.2000 ;
	    RECT 113.4000 18.1000 113.8000 18.2000 ;
	    RECT 106.2000 17.8000 113.8000 18.1000 ;
	    RECT 123.8000 18.1000 124.2000 18.2000 ;
	    RECT 131.0000 18.1000 131.3000 18.8000 ;
	    RECT 123.8000 17.8000 131.3000 18.1000 ;
	    RECT 143.8000 17.8000 144.2000 18.2000 ;
	    RECT 1.4000 17.1000 1.8000 17.2000 ;
	    RECT 3.0000 17.1000 3.4000 17.2000 ;
	    RECT 1.4000 16.8000 3.4000 17.1000 ;
	    RECT 6.2000 17.1000 6.6000 17.2000 ;
	    RECT 8.6000 17.1000 9.0000 17.2000 ;
	    RECT 6.2000 16.8000 9.0000 17.1000 ;
	    RECT 19.8000 17.1000 20.2000 17.2000 ;
	    RECT 21.4000 17.1000 21.7000 17.8000 ;
	    RECT 19.8000 16.8000 21.7000 17.1000 ;
	    RECT 22.2000 17.1000 22.6000 17.2000 ;
	    RECT 23.0000 17.1000 23.4000 17.2000 ;
	    RECT 22.2000 16.8000 23.4000 17.1000 ;
	    RECT 28.6000 17.1000 29.0000 17.2000 ;
	    RECT 30.2000 17.1000 30.6000 17.2000 ;
	    RECT 28.6000 16.8000 30.6000 17.1000 ;
	    RECT 31.8000 17.1000 32.2000 17.2000 ;
	    RECT 46.2000 17.1000 46.6000 17.2000 ;
	    RECT 31.8000 16.8000 46.6000 17.1000 ;
	    RECT 58.2000 17.1000 58.6000 17.2000 ;
	    RECT 63.8000 17.1000 64.2000 17.2000 ;
	    RECT 58.2000 16.8000 64.2000 17.1000 ;
	    RECT 64.6000 17.1000 65.0000 17.2000 ;
	    RECT 67.0000 17.1000 67.4000 17.2000 ;
	    RECT 64.6000 16.8000 67.4000 17.1000 ;
	    RECT 68.6000 17.1000 69.0000 17.2000 ;
	    RECT 73.4000 17.1000 73.8000 17.2000 ;
	    RECT 81.4000 17.1000 81.8000 17.2000 ;
	    RECT 68.6000 16.8000 72.9000 17.1000 ;
	    RECT 73.4000 16.8000 81.8000 17.1000 ;
	    RECT 83.8000 17.1000 84.2000 17.2000 ;
	    RECT 85.4000 17.1000 85.8000 17.2000 ;
	    RECT 83.8000 16.8000 85.8000 17.1000 ;
	    RECT 87.8000 16.8000 88.2000 17.2000 ;
	    RECT 93.4000 17.1000 93.8000 17.2000 ;
	    RECT 97.4000 17.1000 97.8000 17.2000 ;
	    RECT 93.4000 16.8000 97.8000 17.1000 ;
	    RECT 100.6000 17.1000 101.0000 17.2000 ;
	    RECT 101.4000 17.1000 101.8000 17.2000 ;
	    RECT 100.6000 16.8000 101.8000 17.1000 ;
	    RECT 112.6000 17.1000 113.0000 17.2000 ;
	    RECT 122.2000 17.1000 122.6000 17.2000 ;
	    RECT 112.6000 16.8000 122.6000 17.1000 ;
	    RECT 127.0000 17.1000 127.4000 17.2000 ;
	    RECT 143.8000 17.1000 144.1000 17.8000 ;
	    RECT 127.0000 16.8000 144.1000 17.1000 ;
	    RECT 151.0000 17.1000 151.4000 17.2000 ;
	    RECT 159.0000 17.1000 159.4000 17.2000 ;
	    RECT 151.0000 16.8000 159.4000 17.1000 ;
	    RECT 72.6000 16.2000 72.9000 16.8000 ;
	    RECT 6.2000 15.8000 6.6000 16.2000 ;
	    RECT 16.6000 16.1000 17.0000 16.2000 ;
	    RECT 17.4000 16.1000 17.8000 16.2000 ;
	    RECT 12.6000 15.8000 17.8000 16.1000 ;
	    RECT 35.0000 15.8000 35.4000 16.2000 ;
	    RECT 38.2000 15.8000 38.6000 16.2000 ;
	    RECT 72.6000 15.8000 73.0000 16.2000 ;
	    RECT 82.2000 16.1000 82.6000 16.2000 ;
	    RECT 80.6000 15.8000 82.6000 16.1000 ;
	    RECT 85.4000 16.1000 85.8000 16.2000 ;
	    RECT 87.8000 16.1000 88.1000 16.8000 ;
	    RECT 85.4000 15.8000 88.1000 16.1000 ;
	    RECT 94.2000 15.8000 94.6000 16.2000 ;
	    RECT 115.8000 15.8000 116.2000 16.2000 ;
	    RECT 116.6000 16.1000 117.0000 16.2000 ;
	    RECT 124.6000 16.1000 125.0000 16.2000 ;
	    RECT 127.0000 16.1000 127.4000 16.2000 ;
	    RECT 116.6000 15.8000 119.3000 16.1000 ;
	    RECT 124.6000 15.8000 127.4000 16.1000 ;
	    RECT 134.2000 15.8000 134.6000 16.2000 ;
	    RECT 136.6000 16.1000 137.0000 16.2000 ;
	    RECT 141.4000 16.1000 141.8000 16.2000 ;
	    RECT 136.6000 15.8000 141.8000 16.1000 ;
	    RECT 150.2000 15.8000 150.6000 16.2000 ;
	    RECT 152.6000 16.1000 153.0000 16.2000 ;
	    RECT 153.4000 16.1000 153.8000 16.2000 ;
	    RECT 152.6000 15.8000 153.8000 16.1000 ;
	    RECT 159.8000 16.1000 160.2000 16.2000 ;
	    RECT 163.8000 16.1000 164.2000 16.2000 ;
	    RECT 159.8000 15.8000 164.2000 16.1000 ;
	    RECT 5.4000 15.1000 5.8000 15.2000 ;
	    RECT 6.2000 15.1000 6.5000 15.8000 ;
	    RECT 5.4000 14.8000 6.5000 15.1000 ;
	    RECT 12.6000 15.2000 12.9000 15.8000 ;
	    RECT 12.6000 14.8000 13.0000 15.2000 ;
	    RECT 18.2000 15.1000 18.6000 15.2000 ;
	    RECT 19.0000 15.1000 19.4000 15.2000 ;
	    RECT 18.2000 14.8000 19.4000 15.1000 ;
	    RECT 23.8000 14.8000 24.2000 15.2000 ;
	    RECT 27.8000 15.1000 28.2000 15.2000 ;
	    RECT 33.4000 15.1000 33.8000 15.2000 ;
	    RECT 35.0000 15.1000 35.3000 15.8000 ;
	    RECT 27.8000 14.8000 32.1000 15.1000 ;
	    RECT 33.4000 14.8000 35.3000 15.1000 ;
	    RECT 36.6000 15.1000 37.0000 15.2000 ;
	    RECT 38.2000 15.1000 38.5000 15.8000 ;
	    RECT 80.6000 15.2000 80.9000 15.8000 ;
	    RECT 36.6000 14.8000 38.5000 15.1000 ;
	    RECT 39.0000 14.8000 41.7000 15.1000 ;
	    RECT 23.8000 14.2000 24.1000 14.8000 ;
	    RECT 4.6000 14.1000 5.0000 14.2000 ;
	    RECT 11.0000 14.1000 11.4000 14.2000 ;
	    RECT 4.6000 13.8000 11.4000 14.1000 ;
	    RECT 15.8000 14.1000 16.2000 14.2000 ;
	    RECT 23.0000 14.1000 23.4000 14.2000 ;
	    RECT 15.8000 13.8000 23.4000 14.1000 ;
	    RECT 23.8000 13.8000 24.2000 14.2000 ;
	    RECT 24.6000 14.1000 25.0000 14.2000 ;
	    RECT 27.0000 14.1000 27.4000 14.2000 ;
	    RECT 24.6000 13.8000 27.4000 14.1000 ;
	    RECT 31.0000 13.8000 31.4000 14.2000 ;
	    RECT 31.8000 14.1000 32.1000 14.8000 ;
	    RECT 39.0000 14.1000 39.3000 14.8000 ;
	    RECT 31.8000 13.8000 39.3000 14.1000 ;
	    RECT 41.4000 14.2000 41.7000 14.8000 ;
	    RECT 44.6000 14.8000 45.0000 15.2000 ;
	    RECT 47.8000 14.8000 48.2000 15.2000 ;
	    RECT 51.8000 15.1000 52.2000 15.2000 ;
	    RECT 57.4000 15.1000 57.8000 15.2000 ;
	    RECT 66.2000 15.1000 66.6000 15.2000 ;
	    RECT 51.8000 14.8000 52.9000 15.1000 ;
	    RECT 57.4000 14.8000 66.6000 15.1000 ;
	    RECT 69.4000 15.1000 69.8000 15.2000 ;
	    RECT 73.4000 15.1000 73.8000 15.2000 ;
	    RECT 69.4000 14.8000 73.8000 15.1000 ;
	    RECT 75.8000 15.1000 76.2000 15.2000 ;
	    RECT 78.2000 15.1000 78.6000 15.2000 ;
	    RECT 75.8000 14.8000 78.6000 15.1000 ;
	    RECT 80.6000 14.8000 81.0000 15.2000 ;
	    RECT 81.4000 15.1000 81.8000 15.2000 ;
	    RECT 91.0000 15.1000 91.4000 15.2000 ;
	    RECT 81.4000 14.8000 91.4000 15.1000 ;
	    RECT 92.6000 15.1000 93.0000 15.2000 ;
	    RECT 94.2000 15.1000 94.5000 15.8000 ;
	    RECT 92.6000 14.8000 94.5000 15.1000 ;
	    RECT 103.8000 15.1000 104.2000 15.2000 ;
	    RECT 107.8000 15.1000 108.2000 15.2000 ;
	    RECT 103.8000 14.8000 108.2000 15.1000 ;
	    RECT 110.2000 15.1000 110.6000 15.2000 ;
	    RECT 115.8000 15.1000 116.1000 15.8000 ;
	    RECT 110.2000 14.8000 116.1000 15.1000 ;
	    RECT 119.0000 15.2000 119.3000 15.8000 ;
	    RECT 119.0000 14.8000 119.4000 15.2000 ;
	    RECT 129.4000 15.1000 129.8000 15.2000 ;
	    RECT 134.2000 15.1000 134.5000 15.8000 ;
	    RECT 129.4000 14.8000 134.5000 15.1000 ;
	    RECT 149.4000 15.1000 149.8000 15.2000 ;
	    RECT 150.2000 15.1000 150.5000 15.8000 ;
	    RECT 149.4000 14.8000 150.5000 15.1000 ;
	    RECT 151.0000 15.1000 151.4000 15.2000 ;
	    RECT 154.2000 15.1000 154.6000 15.2000 ;
	    RECT 151.0000 14.8000 154.6000 15.1000 ;
	    RECT 157.4000 15.1000 157.8000 15.2000 ;
	    RECT 158.2000 15.1000 158.6000 15.2000 ;
	    RECT 157.4000 14.8000 158.6000 15.1000 ;
	    RECT 162.2000 15.1000 162.6000 15.2000 ;
	    RECT 163.0000 15.1000 163.4000 15.2000 ;
	    RECT 162.2000 14.8000 163.4000 15.1000 ;
	    RECT 41.4000 13.8000 41.8000 14.2000 ;
	    RECT 44.6000 14.1000 44.9000 14.8000 ;
	    RECT 47.8000 14.1000 48.1000 14.8000 ;
	    RECT 52.6000 14.2000 52.9000 14.8000 ;
	    RECT 44.6000 13.8000 48.1000 14.1000 ;
	    RECT 50.2000 14.1000 50.6000 14.2000 ;
	    RECT 51.8000 14.1000 52.2000 14.2000 ;
	    RECT 50.2000 13.8000 52.2000 14.1000 ;
	    RECT 52.6000 13.8000 53.0000 14.2000 ;
	    RECT 138.2000 14.1000 138.6000 14.2000 ;
	    RECT 140.6000 14.1000 141.0000 14.2000 ;
	    RECT 138.2000 13.8000 141.0000 14.1000 ;
	    RECT 147.8000 14.1000 148.2000 14.2000 ;
	    RECT 159.8000 14.1000 160.2000 14.2000 ;
	    RECT 147.8000 13.8000 160.2000 14.1000 ;
	    RECT 166.2000 14.1000 166.6000 14.2000 ;
	    RECT 166.2000 13.8000 169.7000 14.1000 ;
	    RECT 10.2000 13.1000 10.6000 13.2000 ;
	    RECT 17.4000 13.1000 17.8000 13.2000 ;
	    RECT 10.2000 12.8000 17.8000 13.1000 ;
	    RECT 31.0000 13.1000 31.3000 13.8000 ;
	    RECT 169.4000 13.2000 169.7000 13.8000 ;
	    RECT 36.6000 13.1000 37.0000 13.2000 ;
	    RECT 39.8000 13.1000 40.2000 13.2000 ;
	    RECT 41.4000 13.1000 41.8000 13.2000 ;
	    RECT 43.0000 13.1000 43.4000 13.2000 ;
	    RECT 45.4000 13.1000 45.8000 13.2000 ;
	    RECT 31.0000 12.8000 45.8000 13.1000 ;
	    RECT 74.2000 13.1000 74.6000 13.2000 ;
	    RECT 75.8000 13.1000 76.2000 13.2000 ;
	    RECT 74.2000 12.8000 76.2000 13.1000 ;
	    RECT 91.0000 13.1000 91.4000 13.2000 ;
	    RECT 108.6000 13.1000 109.0000 13.2000 ;
	    RECT 91.0000 12.8000 109.0000 13.1000 ;
	    RECT 109.4000 13.1000 109.8000 13.2000 ;
	    RECT 112.6000 13.1000 113.0000 13.2000 ;
	    RECT 109.4000 12.8000 113.0000 13.1000 ;
	    RECT 115.0000 13.1000 115.4000 13.2000 ;
	    RECT 115.8000 13.1000 116.2000 13.2000 ;
	    RECT 115.0000 12.8000 116.2000 13.1000 ;
	    RECT 130.2000 12.8000 130.6000 13.2000 ;
	    RECT 169.4000 12.8000 169.8000 13.2000 ;
	    RECT 72.6000 12.1000 73.0000 12.2000 ;
	    RECT 83.0000 12.1000 83.4000 12.2000 ;
	    RECT 72.6000 11.8000 83.4000 12.1000 ;
	    RECT 87.8000 12.1000 88.2000 12.2000 ;
	    RECT 100.6000 12.1000 101.0000 12.2000 ;
	    RECT 87.8000 11.8000 101.0000 12.1000 ;
	    RECT 103.8000 12.1000 104.2000 12.2000 ;
	    RECT 106.2000 12.1000 106.6000 12.2000 ;
	    RECT 103.8000 11.8000 106.6000 12.1000 ;
	    RECT 124.6000 12.1000 125.0000 12.2000 ;
	    RECT 130.2000 12.1000 130.5000 12.8000 ;
	    RECT 133.4000 12.1000 133.8000 12.2000 ;
	    RECT 136.6000 12.1000 137.0000 12.2000 ;
	    RECT 143.8000 12.1000 144.2000 12.2000 ;
	    RECT 124.6000 11.8000 144.2000 12.1000 ;
	    RECT 159.0000 12.1000 159.4000 12.2000 ;
	    RECT 167.8000 12.1000 168.2000 12.2000 ;
	    RECT 159.0000 11.8000 168.2000 12.1000 ;
	    RECT 34.2000 11.1000 34.6000 11.2000 ;
	    RECT 67.0000 11.1000 67.4000 11.2000 ;
	    RECT 34.2000 10.8000 67.4000 11.1000 ;
	    RECT 84.6000 11.1000 85.0000 11.2000 ;
	    RECT 90.2000 11.1000 90.6000 11.2000 ;
	    RECT 96.6000 11.1000 97.0000 11.2000 ;
	    RECT 84.6000 10.8000 97.0000 11.1000 ;
	    RECT 118.2000 11.1000 118.6000 11.2000 ;
	    RECT 119.8000 11.1000 120.2000 11.2000 ;
	    RECT 121.4000 11.1000 121.8000 11.2000 ;
	    RECT 118.2000 10.8000 121.8000 11.1000 ;
	    RECT 123.8000 11.1000 124.2000 11.2000 ;
	    RECT 135.8000 11.1000 136.2000 11.2000 ;
	    RECT 123.8000 10.8000 136.2000 11.1000 ;
	    RECT 136.6000 11.1000 137.0000 11.2000 ;
	    RECT 140.6000 11.1000 141.0000 11.2000 ;
	    RECT 136.6000 10.8000 141.0000 11.1000 ;
	    RECT 141.4000 11.1000 141.8000 11.2000 ;
	    RECT 153.4000 11.1000 153.8000 11.2000 ;
	    RECT 141.4000 10.8000 153.8000 11.1000 ;
	    RECT 154.2000 11.1000 154.6000 11.2000 ;
	    RECT 162.2000 11.1000 162.6000 11.2000 ;
	    RECT 154.2000 10.8000 162.6000 11.1000 ;
	    RECT 138.2000 10.1000 138.6000 10.2000 ;
	    RECT 139.8000 10.1000 140.2000 10.2000 ;
	    RECT 142.2000 10.1000 142.6000 10.2000 ;
	    RECT 152.6000 10.1000 153.0000 10.2000 ;
	    RECT 155.0000 10.1000 155.4000 10.2000 ;
	    RECT 167.0000 10.1000 167.4000 10.2000 ;
	    RECT 138.2000 9.8000 167.4000 10.1000 ;
	    RECT 12.6000 8.8000 13.0000 9.2000 ;
	    RECT 80.6000 8.8000 81.0000 9.2000 ;
	    RECT 99.0000 9.1000 99.4000 9.2000 ;
	    RECT 103.0000 9.1000 103.4000 9.2000 ;
	    RECT 104.6000 9.1000 105.0000 9.2000 ;
	    RECT 110.2000 9.1000 110.6000 9.2000 ;
	    RECT 119.8000 9.1000 120.2000 9.2000 ;
	    RECT 99.0000 8.8000 120.2000 9.1000 ;
	    RECT 133.4000 9.1000 133.8000 9.2000 ;
	    RECT 138.2000 9.1000 138.6000 9.2000 ;
	    RECT 133.4000 8.8000 138.6000 9.1000 ;
	    RECT 146.2000 9.1000 146.6000 9.2000 ;
	    RECT 148.6000 9.1000 149.0000 9.2000 ;
	    RECT 151.8000 9.1000 152.2000 9.2000 ;
	    RECT 155.0000 9.1000 155.4000 9.2000 ;
	    RECT 166.2000 9.1000 166.6000 9.2000 ;
	    RECT 146.2000 8.8000 166.6000 9.1000 ;
	    RECT 8.6000 8.1000 9.0000 8.2000 ;
	    RECT 12.6000 8.1000 12.9000 8.8000 ;
	    RECT 8.6000 7.8000 12.9000 8.1000 ;
	    RECT 54.2000 8.1000 54.6000 8.2000 ;
	    RECT 55.0000 8.1000 55.4000 8.2000 ;
	    RECT 58.2000 8.1000 58.6000 8.2000 ;
	    RECT 60.6000 8.1000 61.0000 8.2000 ;
	    RECT 70.2000 8.1000 70.6000 8.2000 ;
	    RECT 54.2000 7.8000 70.6000 8.1000 ;
	    RECT 71.0000 8.1000 71.4000 8.2000 ;
	    RECT 75.0000 8.1000 75.4000 8.2000 ;
	    RECT 80.6000 8.1000 80.9000 8.8000 ;
	    RECT 84.6000 8.1000 85.0000 8.2000 ;
	    RECT 71.0000 7.8000 85.0000 8.1000 ;
	    RECT 99.8000 7.8000 100.2000 8.2000 ;
	    RECT 157.4000 8.1000 157.8000 8.2000 ;
	    RECT 160.6000 8.1000 161.0000 8.2000 ;
	    RECT 157.4000 7.8000 161.0000 8.1000 ;
	    RECT 1.4000 7.1000 1.8000 7.2000 ;
	    RECT 3.8000 7.1000 4.2000 7.2000 ;
	    RECT 8.6000 7.1000 9.0000 7.2000 ;
	    RECT 1.4000 6.8000 9.0000 7.1000 ;
	    RECT 22.2000 7.1000 22.6000 7.2000 ;
	    RECT 25.4000 7.1000 25.8000 7.2000 ;
	    RECT 27.8000 7.1000 28.2000 7.2000 ;
	    RECT 31.8000 7.1000 32.2000 7.2000 ;
	    RECT 34.2000 7.1000 34.6000 7.2000 ;
	    RECT 35.8000 7.1000 36.2000 7.2000 ;
	    RECT 22.2000 6.8000 36.2000 7.1000 ;
	    RECT 37.4000 7.1000 37.8000 7.2000 ;
	    RECT 42.2000 7.1000 42.6000 7.2000 ;
	    RECT 43.8000 7.1000 44.2000 7.2000 ;
	    RECT 47.8000 7.1000 48.2000 7.2000 ;
	    RECT 37.4000 6.8000 43.3000 7.1000 ;
	    RECT 43.8000 6.8000 48.2000 7.1000 ;
	    RECT 88.6000 7.1000 89.0000 7.2000 ;
	    RECT 92.6000 7.1000 93.0000 7.2000 ;
	    RECT 88.6000 6.8000 93.0000 7.1000 ;
	    RECT 96.6000 7.1000 97.0000 7.2000 ;
	    RECT 99.8000 7.1000 100.1000 7.8000 ;
	    RECT 96.6000 6.8000 100.1000 7.1000 ;
	    RECT 108.6000 7.1000 109.0000 7.2000 ;
	    RECT 111.8000 7.1000 112.2000 7.2000 ;
	    RECT 108.6000 6.8000 112.2000 7.1000 ;
	    RECT 116.6000 7.1000 117.0000 7.2000 ;
	    RECT 123.0000 7.1000 123.4000 7.2000 ;
	    RECT 124.6000 7.1000 125.0000 7.2000 ;
	    RECT 116.6000 6.8000 125.0000 7.1000 ;
	    RECT 135.0000 7.1000 135.4000 7.2000 ;
	    RECT 149.4000 7.1000 149.8000 7.2000 ;
	    RECT 135.0000 6.8000 149.8000 7.1000 ;
	    RECT 167.0000 7.1000 167.4000 7.2000 ;
	    RECT 168.6000 7.1000 169.0000 7.2000 ;
	    RECT 167.0000 6.8000 169.0000 7.1000 ;
	    RECT 170.2000 7.1000 170.6000 7.2000 ;
	    RECT 170.2000 7.0000 171.3000 7.1000 ;
	    RECT 170.2000 6.8000 171.4000 7.0000 ;
	    RECT 171.0000 6.6000 171.4000 6.8000 ;
	    RECT 2.2000 6.1000 2.6000 6.2000 ;
	    RECT 15.8000 6.1000 16.2000 6.2000 ;
	    RECT 2.2000 5.8000 16.2000 6.1000 ;
	    RECT 98.2000 6.1000 98.6000 6.2000 ;
	    RECT 100.6000 6.1000 101.0000 6.2000 ;
	    RECT 98.2000 5.8000 101.0000 6.1000 ;
	    RECT 129.4000 6.1000 129.8000 6.2000 ;
	    RECT 135.8000 6.1000 136.2000 6.2000 ;
	    RECT 129.4000 5.8000 136.2000 6.1000 ;
	    RECT 3.8000 5.1000 4.2000 5.2000 ;
	    RECT 7.0000 5.1000 7.4000 5.2000 ;
	    RECT 3.8000 4.8000 7.4000 5.1000 ;
	    RECT 34.2000 5.1000 34.6000 5.2000 ;
	    RECT 35.0000 5.1000 35.4000 5.2000 ;
	    RECT 34.2000 4.8000 35.4000 5.1000 ;
	    RECT 41.4000 4.8000 41.8000 5.2000 ;
	    RECT 42.2000 5.1000 42.6000 5.2000 ;
	    RECT 43.8000 5.1000 44.2000 5.2000 ;
	    RECT 42.2000 4.8000 44.2000 5.1000 ;
	    RECT 17.4000 4.1000 17.8000 4.2000 ;
	    RECT 41.4000 4.1000 41.7000 4.8000 ;
	    RECT 17.4000 3.8000 41.7000 4.1000 ;
	    RECT 27.8000 2.1000 28.2000 2.2000 ;
	    RECT 45.4000 2.1000 45.8000 2.2000 ;
	    RECT 27.8000 1.8000 45.8000 2.1000 ;
         LAYER metal4 ;
	    RECT 155.0000 155.8000 155.4000 156.2000 ;
	    RECT 123.0000 154.8000 123.4000 155.2000 ;
	    RECT 131.8000 154.8000 132.2000 155.2000 ;
	    RECT 18.2000 153.8000 18.6000 154.2000 ;
	    RECT 36.6000 154.1000 37.0000 154.2000 ;
	    RECT 37.4000 154.1000 37.8000 154.2000 ;
	    RECT 36.6000 153.8000 37.8000 154.1000 ;
	    RECT 47.0000 154.1000 47.4000 154.2000 ;
	    RECT 47.8000 154.1000 48.2000 154.2000 ;
	    RECT 47.0000 153.8000 48.2000 154.1000 ;
	    RECT 109.4000 153.8000 109.8000 154.2000 ;
	    RECT 7.0000 148.8000 7.4000 149.2000 ;
	    RECT 5.4000 146.8000 5.8000 147.2000 ;
	    RECT 5.4000 137.2000 5.7000 146.8000 ;
	    RECT 6.2000 144.1000 6.6000 144.2000 ;
	    RECT 7.0000 144.1000 7.3000 148.8000 ;
	    RECT 6.2000 143.8000 7.3000 144.1000 ;
	    RECT 5.4000 136.8000 5.8000 137.2000 ;
	    RECT 18.2000 134.2000 18.5000 153.8000 ;
	    RECT 98.2000 152.8000 98.6000 153.2000 ;
	    RECT 55.0000 151.8000 55.4000 152.2000 ;
	    RECT 87.0000 151.8000 87.4000 152.2000 ;
	    RECT 96.6000 152.1000 97.0000 152.2000 ;
	    RECT 97.4000 152.1000 97.8000 152.2000 ;
	    RECT 96.6000 151.8000 97.8000 152.1000 ;
	    RECT 47.8000 144.8000 48.2000 145.2000 ;
	    RECT 18.2000 133.8000 18.6000 134.2000 ;
	    RECT 27.8000 127.1000 28.2000 127.2000 ;
	    RECT 27.8000 126.8000 28.9000 127.1000 ;
	    RECT 28.6000 124.2000 28.9000 126.8000 ;
	    RECT 28.6000 123.8000 29.0000 124.2000 ;
	    RECT 2.2000 121.8000 2.6000 122.2000 ;
	    RECT 2.2000 103.2000 2.5000 121.8000 ;
	    RECT 32.6000 118.8000 33.0000 119.2000 ;
	    RECT 21.4000 117.8000 21.8000 118.2000 ;
	    RECT 15.8000 115.8000 16.2000 116.2000 ;
	    RECT 2.2000 102.8000 2.6000 103.2000 ;
	    RECT 3.0000 101.8000 3.4000 102.2000 ;
	    RECT 3.0000 65.2000 3.3000 101.8000 ;
	    RECT 3.8000 76.8000 4.2000 77.2000 ;
	    RECT 3.0000 64.8000 3.4000 65.2000 ;
	    RECT 3.8000 58.2000 4.1000 76.8000 ;
	    RECT 15.0000 66.1000 15.4000 66.2000 ;
	    RECT 15.8000 66.1000 16.1000 115.8000 ;
	    RECT 19.8000 106.8000 20.2000 107.2000 ;
	    RECT 19.8000 106.2000 20.1000 106.8000 ;
	    RECT 19.8000 105.8000 20.2000 106.2000 ;
	    RECT 19.0000 87.1000 19.4000 87.2000 ;
	    RECT 19.8000 87.1000 20.2000 87.2000 ;
	    RECT 19.0000 86.8000 20.2000 87.1000 ;
	    RECT 15.0000 65.8000 16.1000 66.1000 ;
	    RECT 18.2000 60.8000 18.6000 61.2000 ;
	    RECT 3.8000 57.8000 4.2000 58.2000 ;
	    RECT 12.6000 57.1000 13.0000 57.2000 ;
	    RECT 13.4000 57.1000 13.8000 57.2000 ;
	    RECT 12.6000 56.8000 13.8000 57.1000 ;
	    RECT 15.8000 56.8000 16.2000 57.2000 ;
	    RECT 15.8000 55.2000 16.1000 56.8000 ;
	    RECT 15.8000 54.8000 16.2000 55.2000 ;
	    RECT 18.2000 54.1000 18.5000 60.8000 ;
	    RECT 21.4000 58.1000 21.7000 117.8000 ;
	    RECT 32.6000 104.2000 32.9000 118.8000 ;
	    RECT 47.8000 116.2000 48.1000 144.8000 ;
	    RECT 55.0000 136.2000 55.3000 151.8000 ;
	    RECT 81.4000 137.8000 81.8000 138.2000 ;
	    RECT 53.4000 136.1000 53.8000 136.2000 ;
	    RECT 54.2000 136.1000 54.6000 136.2000 ;
	    RECT 53.4000 135.8000 54.6000 136.1000 ;
	    RECT 55.0000 135.8000 55.4000 136.2000 ;
	    RECT 56.6000 136.1000 57.0000 136.2000 ;
	    RECT 57.4000 136.1000 57.8000 136.2000 ;
	    RECT 56.6000 135.8000 57.8000 136.1000 ;
	    RECT 76.6000 134.8000 77.0000 135.2000 ;
	    RECT 69.4000 127.8000 69.8000 128.2000 ;
	    RECT 69.4000 117.2000 69.7000 127.8000 ;
	    RECT 68.6000 116.8000 69.0000 117.2000 ;
	    RECT 69.4000 116.8000 69.8000 117.2000 ;
	    RECT 47.8000 115.8000 48.2000 116.2000 ;
	    RECT 39.0000 106.1000 39.4000 106.2000 ;
	    RECT 39.8000 106.1000 40.2000 106.2000 ;
	    RECT 39.0000 105.8000 40.2000 106.1000 ;
	    RECT 32.6000 103.8000 33.0000 104.2000 ;
	    RECT 47.8000 97.2000 48.1000 115.8000 ;
	    RECT 67.8000 106.8000 68.2000 107.2000 ;
	    RECT 67.8000 105.2000 68.1000 106.8000 ;
	    RECT 67.8000 104.8000 68.2000 105.2000 ;
	    RECT 58.2000 103.8000 58.6000 104.2000 ;
	    RECT 57.4000 100.8000 57.8000 101.2000 ;
	    RECT 47.8000 96.8000 48.2000 97.2000 ;
	    RECT 23.8000 95.8000 24.2000 96.2000 ;
	    RECT 22.2000 86.8000 22.6000 87.2000 ;
	    RECT 22.2000 86.2000 22.5000 86.8000 ;
	    RECT 22.2000 85.8000 22.6000 86.2000 ;
	    RECT 23.8000 85.2000 24.1000 95.8000 ;
	    RECT 57.4000 95.2000 57.7000 100.8000 ;
	    RECT 58.2000 100.2000 58.5000 103.8000 ;
	    RECT 58.2000 99.8000 58.6000 100.2000 ;
	    RECT 68.6000 95.2000 68.9000 116.8000 ;
	    RECT 75.8000 109.8000 76.2000 110.2000 ;
	    RECT 29.4000 95.1000 29.8000 95.2000 ;
	    RECT 30.2000 95.1000 30.6000 95.2000 ;
	    RECT 29.4000 94.8000 30.6000 95.1000 ;
	    RECT 36.6000 95.1000 37.0000 95.2000 ;
	    RECT 37.4000 95.1000 37.8000 95.2000 ;
	    RECT 36.6000 94.8000 37.8000 95.1000 ;
	    RECT 57.4000 94.8000 57.8000 95.2000 ;
	    RECT 68.6000 94.8000 69.0000 95.2000 ;
	    RECT 42.2000 94.1000 42.6000 94.2000 ;
	    RECT 43.0000 94.1000 43.4000 94.2000 ;
	    RECT 42.2000 93.8000 43.4000 94.1000 ;
	    RECT 44.6000 93.8000 45.0000 94.2000 ;
	    RECT 32.6000 87.8000 33.0000 88.2000 ;
	    RECT 30.2000 86.8000 30.6000 87.2000 ;
	    RECT 24.6000 85.8000 25.0000 86.2000 ;
	    RECT 25.4000 86.1000 25.8000 86.2000 ;
	    RECT 26.2000 86.1000 26.6000 86.2000 ;
	    RECT 25.4000 85.8000 26.6000 86.1000 ;
	    RECT 29.4000 86.1000 29.8000 86.2000 ;
	    RECT 30.2000 86.1000 30.5000 86.8000 ;
	    RECT 29.4000 85.8000 30.5000 86.1000 ;
	    RECT 32.6000 86.2000 32.9000 87.8000 ;
	    RECT 32.6000 85.8000 33.0000 86.2000 ;
	    RECT 34.2000 86.1000 34.6000 86.2000 ;
	    RECT 35.0000 86.1000 35.4000 86.2000 ;
	    RECT 34.2000 85.8000 35.4000 86.1000 ;
	    RECT 43.8000 85.8000 44.2000 86.2000 ;
	    RECT 24.6000 85.2000 24.9000 85.8000 ;
	    RECT 43.8000 85.2000 44.1000 85.8000 ;
	    RECT 23.8000 84.8000 24.2000 85.2000 ;
	    RECT 24.6000 84.8000 25.0000 85.2000 ;
	    RECT 43.8000 84.8000 44.2000 85.2000 ;
	    RECT 44.6000 66.2000 44.9000 93.8000 ;
	    RECT 75.0000 93.1000 75.4000 93.2000 ;
	    RECT 75.8000 93.1000 76.1000 109.8000 ;
	    RECT 76.6000 104.2000 76.9000 134.8000 ;
	    RECT 77.4000 130.8000 77.8000 131.2000 ;
	    RECT 76.6000 103.8000 77.0000 104.2000 ;
	    RECT 77.4000 97.2000 77.7000 130.8000 ;
	    RECT 78.2000 114.8000 78.6000 115.2000 ;
	    RECT 77.4000 96.8000 77.8000 97.2000 ;
	    RECT 75.0000 92.8000 76.1000 93.1000 ;
	    RECT 76.6000 95.8000 77.0000 96.2000 ;
	    RECT 67.0000 86.8000 67.4000 87.2000 ;
	    RECT 64.6000 84.8000 65.0000 85.2000 ;
	    RECT 64.6000 82.2000 64.9000 84.8000 ;
	    RECT 64.6000 81.8000 65.0000 82.2000 ;
	    RECT 59.0000 79.8000 59.4000 80.2000 ;
	    RECT 59.0000 66.2000 59.3000 79.8000 ;
	    RECT 44.6000 65.8000 45.0000 66.2000 ;
	    RECT 59.0000 65.8000 59.4000 66.2000 ;
	    RECT 67.0000 64.2000 67.3000 86.8000 ;
	    RECT 75.0000 86.1000 75.4000 86.2000 ;
	    RECT 75.8000 86.1000 76.2000 86.2000 ;
	    RECT 75.0000 85.8000 76.2000 86.1000 ;
	    RECT 76.6000 85.2000 76.9000 95.8000 ;
	    RECT 76.6000 84.8000 77.0000 85.2000 ;
	    RECT 67.8000 81.8000 68.2000 82.2000 ;
	    RECT 67.8000 71.2000 68.1000 81.8000 ;
	    RECT 69.4000 78.8000 69.8000 79.2000 ;
	    RECT 69.4000 77.2000 69.7000 78.8000 ;
	    RECT 69.4000 76.8000 69.8000 77.2000 ;
	    RECT 78.2000 73.2000 78.5000 114.8000 ;
	    RECT 80.6000 110.1000 81.0000 110.2000 ;
	    RECT 81.4000 110.1000 81.7000 137.8000 ;
	    RECT 80.6000 109.8000 81.7000 110.1000 ;
	    RECT 83.8000 114.8000 84.2000 115.2000 ;
	    RECT 80.6000 107.1000 81.0000 107.2000 ;
	    RECT 81.4000 107.1000 81.8000 107.2000 ;
	    RECT 80.6000 106.8000 81.8000 107.1000 ;
	    RECT 83.0000 98.8000 83.4000 99.2000 ;
	    RECT 79.0000 85.8000 79.4000 86.2000 ;
	    RECT 81.4000 85.8000 81.8000 86.2000 ;
	    RECT 79.0000 85.2000 79.3000 85.8000 ;
	    RECT 79.0000 84.8000 79.4000 85.2000 ;
	    RECT 81.4000 82.2000 81.7000 85.8000 ;
	    RECT 81.4000 81.8000 81.8000 82.2000 ;
	    RECT 83.0000 76.2000 83.3000 98.8000 ;
	    RECT 83.8000 86.2000 84.1000 114.8000 ;
	    RECT 84.6000 104.1000 85.0000 104.2000 ;
	    RECT 85.4000 104.1000 85.8000 104.2000 ;
	    RECT 84.6000 103.8000 85.8000 104.1000 ;
	    RECT 87.0000 86.2000 87.3000 151.8000 ;
	    RECT 95.8000 135.1000 96.2000 135.2000 ;
	    RECT 96.6000 135.1000 97.0000 135.2000 ;
	    RECT 95.8000 134.8000 97.0000 135.1000 ;
	    RECT 98.2000 128.2000 98.5000 152.8000 ;
	    RECT 103.8000 152.1000 104.2000 152.2000 ;
	    RECT 104.6000 152.1000 105.0000 152.2000 ;
	    RECT 103.8000 151.8000 105.0000 152.1000 ;
	    RECT 106.2000 150.8000 106.6000 151.2000 ;
	    RECT 106.2000 144.2000 106.5000 150.8000 ;
	    RECT 106.2000 143.8000 106.6000 144.2000 ;
	    RECT 104.6000 130.1000 105.0000 130.2000 ;
	    RECT 103.8000 129.8000 105.0000 130.1000 ;
	    RECT 98.2000 127.8000 98.6000 128.2000 ;
	    RECT 91.8000 125.8000 92.2000 126.2000 ;
	    RECT 90.2000 111.8000 90.6000 112.2000 ;
	    RECT 90.2000 104.2000 90.5000 111.8000 ;
	    RECT 91.0000 108.8000 91.4000 109.2000 ;
	    RECT 90.2000 103.8000 90.6000 104.2000 ;
	    RECT 83.8000 85.8000 84.2000 86.2000 ;
	    RECT 87.0000 85.8000 87.4000 86.2000 ;
	    RECT 91.0000 85.2000 91.3000 108.8000 ;
	    RECT 91.0000 84.8000 91.4000 85.2000 ;
	    RECT 91.8000 83.2000 92.1000 125.8000 ;
	    RECT 98.2000 124.2000 98.5000 127.8000 ;
	    RECT 103.8000 125.2000 104.1000 129.8000 ;
	    RECT 103.8000 124.8000 104.2000 125.2000 ;
	    RECT 98.2000 123.8000 98.6000 124.2000 ;
	    RECT 96.6000 110.8000 97.0000 111.2000 ;
	    RECT 92.6000 107.8000 93.0000 108.2000 ;
	    RECT 92.6000 84.2000 92.9000 107.8000 ;
	    RECT 96.6000 88.2000 96.9000 110.8000 ;
	    RECT 101.4000 105.8000 101.8000 106.2000 ;
	    RECT 99.0000 95.1000 99.4000 95.2000 ;
	    RECT 99.8000 95.1000 100.2000 95.2000 ;
	    RECT 99.0000 94.8000 100.2000 95.1000 ;
	    RECT 99.8000 92.1000 100.2000 92.2000 ;
	    RECT 99.0000 91.8000 100.2000 92.1000 ;
	    RECT 96.6000 87.8000 97.0000 88.2000 ;
	    RECT 95.8000 86.1000 96.2000 86.2000 ;
	    RECT 96.6000 86.1000 97.0000 86.2000 ;
	    RECT 95.8000 85.8000 97.0000 86.1000 ;
	    RECT 92.6000 83.8000 93.0000 84.2000 ;
	    RECT 91.8000 82.8000 92.2000 83.2000 ;
	    RECT 93.4000 77.1000 93.8000 77.2000 ;
	    RECT 94.2000 77.1000 94.6000 77.2000 ;
	    RECT 93.4000 76.8000 94.6000 77.1000 ;
	    RECT 83.0000 75.8000 83.4000 76.2000 ;
	    RECT 78.2000 72.8000 78.6000 73.2000 ;
	    RECT 67.8000 70.8000 68.2000 71.2000 ;
	    RECT 96.6000 71.1000 97.0000 71.2000 ;
	    RECT 96.6000 70.8000 97.7000 71.1000 ;
	    RECT 67.0000 63.8000 67.4000 64.2000 ;
	    RECT 97.4000 63.2000 97.7000 70.8000 ;
	    RECT 99.0000 64.2000 99.3000 91.8000 ;
	    RECT 101.4000 88.2000 101.7000 105.8000 ;
	    RECT 104.6000 94.1000 105.0000 94.2000 ;
	    RECT 105.4000 94.1000 105.8000 94.2000 ;
	    RECT 104.6000 93.8000 105.8000 94.1000 ;
	    RECT 103.8000 93.1000 104.2000 93.2000 ;
	    RECT 103.8000 92.8000 104.9000 93.1000 ;
	    RECT 101.4000 87.8000 101.8000 88.2000 ;
	    RECT 100.6000 86.8000 101.0000 87.2000 ;
	    RECT 100.6000 86.2000 100.9000 86.8000 ;
	    RECT 100.6000 85.8000 101.0000 86.2000 ;
	    RECT 103.0000 76.8000 103.4000 77.2000 ;
	    RECT 99.0000 63.8000 99.4000 64.2000 ;
	    RECT 26.2000 62.8000 26.6000 63.2000 ;
	    RECT 97.4000 62.8000 97.8000 63.2000 ;
	    RECT 22.2000 58.1000 22.6000 58.2000 ;
	    RECT 21.4000 57.8000 22.6000 58.1000 ;
	    RECT 26.2000 55.2000 26.5000 62.8000 ;
	    RECT 62.2000 59.8000 62.6000 60.2000 ;
	    RECT 62.2000 59.2000 62.5000 59.8000 ;
	    RECT 103.0000 59.2000 103.3000 76.8000 ;
	    RECT 104.6000 62.2000 104.9000 92.8000 ;
	    RECT 109.4000 69.2000 109.7000 153.8000 ;
	    RECT 119.0000 149.8000 119.4000 150.2000 ;
	    RECT 119.0000 145.2000 119.3000 149.8000 ;
	    RECT 119.0000 144.8000 119.4000 145.2000 ;
	    RECT 123.0000 144.2000 123.3000 154.8000 ;
	    RECT 131.0000 153.8000 131.4000 154.2000 ;
	    RECT 131.0000 153.2000 131.3000 153.8000 ;
	    RECT 131.0000 152.8000 131.4000 153.2000 ;
	    RECT 131.8000 147.2000 132.1000 154.8000 ;
	    RECT 141.4000 154.1000 141.8000 154.2000 ;
	    RECT 142.2000 154.1000 142.6000 154.2000 ;
	    RECT 141.4000 153.8000 142.6000 154.1000 ;
	    RECT 131.8000 146.8000 132.2000 147.2000 ;
	    RECT 123.0000 143.8000 123.4000 144.2000 ;
	    RECT 126.2000 136.8000 126.6000 137.2000 ;
	    RECT 130.2000 136.8000 130.6000 137.2000 ;
	    RECT 114.2000 135.1000 114.6000 135.2000 ;
	    RECT 115.0000 135.1000 115.4000 135.2000 ;
	    RECT 114.2000 134.8000 115.4000 135.1000 ;
	    RECT 115.8000 134.8000 116.2000 135.2000 ;
	    RECT 115.8000 131.2000 116.1000 134.8000 ;
	    RECT 121.4000 133.8000 121.8000 134.2000 ;
	    RECT 121.4000 133.2000 121.7000 133.8000 ;
	    RECT 121.4000 132.8000 121.8000 133.2000 ;
	    RECT 115.8000 130.8000 116.2000 131.2000 ;
	    RECT 112.6000 127.8000 113.0000 128.2000 ;
	    RECT 110.2000 127.1000 110.6000 127.2000 ;
	    RECT 111.0000 127.1000 111.4000 127.2000 ;
	    RECT 110.2000 126.8000 111.4000 127.1000 ;
	    RECT 112.6000 126.2000 112.9000 127.8000 ;
	    RECT 113.4000 126.8000 113.8000 127.2000 ;
	    RECT 113.4000 126.2000 113.7000 126.8000 ;
	    RECT 126.2000 126.2000 126.5000 136.8000 ;
	    RECT 130.2000 129.2000 130.5000 136.8000 ;
	    RECT 151.8000 135.8000 152.2000 136.2000 ;
	    RECT 132.6000 134.1000 133.0000 134.2000 ;
	    RECT 133.4000 134.1000 133.8000 134.2000 ;
	    RECT 132.6000 133.8000 133.8000 134.1000 ;
	    RECT 130.2000 128.8000 130.6000 129.2000 ;
	    RECT 135.8000 127.8000 136.2000 128.2000 ;
	    RECT 112.6000 125.8000 113.0000 126.2000 ;
	    RECT 113.4000 125.8000 113.8000 126.2000 ;
	    RECT 122.2000 125.8000 122.6000 126.2000 ;
	    RECT 126.2000 125.8000 126.6000 126.2000 ;
	    RECT 115.0000 106.1000 115.4000 106.2000 ;
	    RECT 115.8000 106.1000 116.2000 106.2000 ;
	    RECT 115.0000 105.8000 116.2000 106.1000 ;
	    RECT 116.6000 105.8000 117.0000 106.2000 ;
	    RECT 110.2000 93.8000 110.6000 94.2000 ;
	    RECT 109.4000 68.8000 109.8000 69.2000 ;
	    RECT 110.2000 63.2000 110.5000 93.8000 ;
	    RECT 116.6000 92.2000 116.9000 105.8000 ;
	    RECT 122.2000 99.2000 122.5000 125.8000 ;
	    RECT 135.8000 102.2000 136.1000 127.8000 ;
	    RECT 146.2000 111.8000 146.6000 112.2000 ;
	    RECT 139.0000 106.8000 139.4000 107.2000 ;
	    RECT 135.8000 101.8000 136.2000 102.2000 ;
	    RECT 122.2000 98.8000 122.6000 99.2000 ;
	    RECT 139.0000 93.2000 139.3000 106.8000 ;
	    RECT 139.0000 92.8000 139.4000 93.2000 ;
	    RECT 115.8000 91.8000 116.2000 92.2000 ;
	    RECT 116.6000 91.8000 117.0000 92.2000 ;
	    RECT 115.8000 90.2000 116.1000 91.8000 ;
	    RECT 146.2000 90.2000 146.5000 111.8000 ;
	    RECT 151.8000 93.2000 152.1000 135.8000 ;
	    RECT 151.8000 92.8000 152.2000 93.2000 ;
	    RECT 155.0000 90.2000 155.3000 155.8000 ;
	    RECT 165.4000 146.8000 165.8000 147.2000 ;
	    RECT 164.6000 142.8000 165.0000 143.2000 ;
	    RECT 158.2000 136.8000 158.6000 137.2000 ;
	    RECT 155.8000 132.8000 156.2000 133.2000 ;
	    RECT 155.8000 129.2000 156.1000 132.8000 ;
	    RECT 155.8000 128.8000 156.2000 129.2000 ;
	    RECT 115.8000 89.8000 116.2000 90.2000 ;
	    RECT 146.2000 89.8000 146.6000 90.2000 ;
	    RECT 155.0000 89.8000 155.4000 90.2000 ;
	    RECT 158.2000 88.2000 158.5000 136.8000 ;
	    RECT 161.4000 133.8000 161.8000 134.2000 ;
	    RECT 161.4000 125.2000 161.7000 133.8000 ;
	    RECT 161.4000 124.8000 161.8000 125.2000 ;
	    RECT 160.6000 113.8000 161.0000 114.2000 ;
	    RECT 158.2000 87.8000 158.6000 88.2000 ;
	    RECT 158.2000 86.8000 158.6000 87.2000 ;
	    RECT 139.0000 77.8000 139.4000 78.2000 ;
	    RECT 139.0000 75.2000 139.3000 77.8000 ;
	    RECT 139.0000 74.8000 139.4000 75.2000 ;
	    RECT 153.4000 74.1000 153.8000 74.2000 ;
	    RECT 152.6000 73.8000 153.8000 74.1000 ;
	    RECT 148.6000 73.1000 149.0000 73.2000 ;
	    RECT 147.8000 72.8000 149.0000 73.1000 ;
	    RECT 110.2000 62.8000 110.6000 63.2000 ;
	    RECT 104.6000 61.8000 105.0000 62.2000 ;
	    RECT 44.6000 59.1000 45.0000 59.2000 ;
	    RECT 45.4000 59.1000 45.8000 59.2000 ;
	    RECT 44.6000 58.8000 45.8000 59.1000 ;
	    RECT 62.2000 58.8000 62.6000 59.2000 ;
	    RECT 103.0000 58.8000 103.4000 59.2000 ;
	    RECT 27.8000 56.8000 28.2000 57.2000 ;
	    RECT 42.2000 56.8000 42.6000 57.2000 ;
	    RECT 70.2000 57.1000 70.6000 57.2000 ;
	    RECT 70.2000 56.8000 71.3000 57.1000 ;
	    RECT 26.2000 54.8000 26.6000 55.2000 ;
	    RECT 19.0000 54.1000 19.4000 54.2000 ;
	    RECT 18.2000 53.8000 19.4000 54.1000 ;
	    RECT 24.6000 50.8000 25.0000 51.2000 ;
	    RECT 24.6000 44.2000 24.9000 50.8000 ;
	    RECT 27.8000 49.2000 28.1000 56.8000 ;
	    RECT 36.6000 56.1000 37.0000 56.2000 ;
	    RECT 37.4000 56.1000 37.8000 56.2000 ;
	    RECT 36.6000 55.8000 37.8000 56.1000 ;
	    RECT 40.6000 55.8000 41.0000 56.2000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 39.0000 55.1000 39.4000 55.2000 ;
	    RECT 38.2000 54.8000 39.4000 55.1000 ;
	    RECT 40.6000 54.2000 40.9000 55.8000 ;
	    RECT 42.2000 55.2000 42.5000 56.8000 ;
	    RECT 63.8000 55.8000 64.2000 56.2000 ;
	    RECT 63.8000 55.2000 64.1000 55.8000 ;
	    RECT 42.2000 54.8000 42.6000 55.2000 ;
	    RECT 58.2000 54.8000 58.6000 55.2000 ;
	    RECT 63.8000 54.8000 64.2000 55.2000 ;
	    RECT 40.6000 53.8000 41.0000 54.2000 ;
	    RECT 27.8000 48.8000 28.2000 49.2000 ;
	    RECT 28.6000 46.8000 29.0000 47.2000 ;
	    RECT 28.6000 46.1000 28.9000 46.8000 ;
	    RECT 29.4000 46.1000 29.8000 46.2000 ;
	    RECT 28.6000 45.8000 29.8000 46.1000 ;
	    RECT 24.6000 43.8000 25.0000 44.2000 ;
	    RECT 25.4000 43.8000 25.8000 44.2000 ;
	    RECT 51.8000 43.8000 52.2000 44.2000 ;
	    RECT 1.4000 36.8000 1.8000 37.2000 ;
	    RECT 1.4000 31.2000 1.7000 36.8000 ;
	    RECT 17.4000 36.1000 17.8000 36.2000 ;
	    RECT 16.6000 35.8000 17.8000 36.1000 ;
	    RECT 21.4000 36.1000 21.8000 36.2000 ;
	    RECT 22.2000 36.1000 22.6000 36.2000 ;
	    RECT 21.4000 35.8000 22.6000 36.1000 ;
	    RECT 11.0000 33.8000 11.4000 34.2000 ;
	    RECT 1.4000 30.8000 1.8000 31.2000 ;
	    RECT 11.0000 27.2000 11.3000 33.8000 ;
	    RECT 11.0000 26.8000 11.4000 27.2000 ;
	    RECT 14.2000 24.1000 14.6000 24.2000 ;
	    RECT 15.0000 24.1000 15.4000 24.2000 ;
	    RECT 14.2000 23.8000 15.4000 24.1000 ;
	    RECT 16.6000 16.2000 16.9000 35.8000 ;
	    RECT 23.0000 35.1000 23.4000 35.2000 ;
	    RECT 23.8000 35.1000 24.2000 35.2000 ;
	    RECT 23.0000 34.8000 24.2000 35.1000 ;
	    RECT 25.4000 24.2000 25.7000 43.8000 ;
	    RECT 51.8000 43.2000 52.1000 43.8000 ;
	    RECT 51.8000 42.8000 52.2000 43.2000 ;
	    RECT 26.2000 35.8000 26.6000 36.2000 ;
	    RECT 26.2000 34.2000 26.5000 35.8000 ;
	    RECT 58.2000 35.2000 58.5000 54.8000 ;
	    RECT 71.0000 43.2000 71.3000 56.8000 ;
	    RECT 75.0000 56.8000 75.4000 57.2000 ;
	    RECT 109.4000 56.8000 109.8000 57.2000 ;
	    RECT 117.4000 56.8000 117.8000 57.2000 ;
	    RECT 71.8000 53.1000 72.2000 53.2000 ;
	    RECT 71.8000 52.8000 72.9000 53.1000 ;
	    RECT 60.6000 43.1000 61.0000 43.2000 ;
	    RECT 61.4000 43.1000 61.8000 43.2000 ;
	    RECT 60.6000 42.8000 61.8000 43.1000 ;
	    RECT 71.0000 42.8000 71.4000 43.2000 ;
	    RECT 72.6000 38.2000 72.9000 52.8000 ;
	    RECT 75.0000 43.2000 75.3000 56.8000 ;
	    RECT 79.0000 54.1000 79.4000 54.2000 ;
	    RECT 78.2000 53.8000 79.4000 54.1000 ;
	    RECT 75.0000 42.8000 75.4000 43.2000 ;
	    RECT 72.6000 37.8000 73.0000 38.2000 ;
	    RECT 78.2000 35.2000 78.5000 53.8000 ;
	    RECT 90.2000 47.1000 90.6000 47.2000 ;
	    RECT 91.0000 47.1000 91.4000 47.2000 ;
	    RECT 90.2000 46.8000 91.4000 47.1000 ;
	    RECT 29.4000 35.1000 29.8000 35.2000 ;
	    RECT 30.2000 35.1000 30.6000 35.2000 ;
	    RECT 29.4000 34.8000 30.6000 35.1000 ;
	    RECT 58.2000 34.8000 58.6000 35.2000 ;
	    RECT 75.8000 34.8000 76.2000 35.2000 ;
	    RECT 78.2000 34.8000 78.6000 35.2000 ;
	    RECT 75.8000 34.2000 76.1000 34.8000 ;
	    RECT 26.2000 33.8000 26.6000 34.2000 ;
	    RECT 57.4000 34.1000 57.8000 34.2000 ;
	    RECT 58.2000 34.1000 58.6000 34.2000 ;
	    RECT 65.4000 34.1000 65.8000 34.2000 ;
	    RECT 57.4000 33.8000 58.6000 34.1000 ;
	    RECT 64.6000 33.8000 65.8000 34.1000 ;
	    RECT 75.8000 33.8000 76.2000 34.2000 ;
	    RECT 97.4000 34.1000 97.8000 34.2000 ;
	    RECT 98.2000 34.1000 98.6000 34.2000 ;
	    RECT 97.4000 33.8000 98.6000 34.1000 ;
	    RECT 103.8000 34.1000 104.2000 34.2000 ;
	    RECT 104.6000 34.1000 105.0000 34.2000 ;
	    RECT 103.8000 33.8000 105.0000 34.1000 ;
	    RECT 26.2000 26.8000 26.6000 27.2000 ;
	    RECT 26.2000 24.2000 26.5000 26.8000 ;
	    RECT 55.0000 25.8000 55.4000 26.2000 ;
	    RECT 24.6000 23.8000 25.0000 24.2000 ;
	    RECT 25.4000 23.8000 25.8000 24.2000 ;
	    RECT 26.2000 23.8000 26.6000 24.2000 ;
	    RECT 24.6000 23.2000 24.9000 23.8000 ;
	    RECT 24.6000 22.8000 25.0000 23.2000 ;
	    RECT 55.0000 22.2000 55.3000 25.8000 ;
	    RECT 64.6000 25.2000 64.9000 33.8000 ;
	    RECT 109.4000 31.2000 109.7000 56.8000 ;
	    RECT 117.4000 42.2000 117.7000 56.8000 ;
	    RECT 137.4000 56.1000 137.8000 56.2000 ;
	    RECT 136.6000 55.8000 137.8000 56.1000 ;
	    RECT 127.0000 50.8000 127.4000 51.2000 ;
	    RECT 125.4000 45.8000 125.8000 46.2000 ;
	    RECT 125.4000 44.1000 125.7000 45.8000 ;
	    RECT 127.0000 44.2000 127.3000 50.8000 ;
	    RECT 136.6000 45.2000 136.9000 55.8000 ;
	    RECT 136.6000 44.8000 137.0000 45.2000 ;
	    RECT 144.6000 44.8000 145.0000 45.2000 ;
	    RECT 125.4000 43.8000 126.5000 44.1000 ;
	    RECT 127.0000 43.8000 127.4000 44.2000 ;
	    RECT 126.2000 42.2000 126.5000 43.8000 ;
	    RECT 117.4000 41.8000 117.8000 42.2000 ;
	    RECT 126.2000 41.8000 126.6000 42.2000 ;
	    RECT 144.6000 41.2000 144.9000 44.8000 ;
	    RECT 147.8000 41.2000 148.1000 72.8000 ;
	    RECT 150.2000 44.8000 150.6000 45.2000 ;
	    RECT 144.6000 40.8000 145.0000 41.2000 ;
	    RECT 147.8000 40.8000 148.2000 41.2000 ;
	    RECT 142.2000 39.8000 142.6000 40.2000 ;
	    RECT 125.4000 32.8000 125.8000 33.2000 ;
	    RECT 109.4000 30.8000 109.8000 31.2000 ;
	    RECT 116.6000 31.1000 117.0000 31.2000 ;
	    RECT 116.6000 30.8000 117.7000 31.1000 ;
	    RECT 110.2000 29.8000 110.6000 30.2000 ;
	    RECT 110.2000 29.2000 110.5000 29.8000 ;
	    RECT 117.4000 29.2000 117.7000 30.8000 ;
	    RECT 110.2000 28.8000 110.6000 29.2000 ;
	    RECT 117.4000 28.8000 117.8000 29.2000 ;
	    RECT 101.4000 27.1000 101.8000 27.2000 ;
	    RECT 100.6000 26.8000 101.8000 27.1000 ;
	    RECT 108.6000 26.8000 109.0000 27.2000 ;
	    RECT 64.6000 24.8000 65.0000 25.2000 ;
	    RECT 100.6000 22.2000 100.9000 26.8000 ;
	    RECT 55.0000 21.8000 55.4000 22.2000 ;
	    RECT 100.6000 21.8000 101.0000 22.2000 ;
	    RECT 18.2000 18.8000 18.6000 19.2000 ;
	    RECT 16.6000 15.8000 17.0000 16.2000 ;
	    RECT 18.2000 15.2000 18.5000 18.8000 ;
	    RECT 22.2000 17.1000 22.6000 17.2000 ;
	    RECT 23.0000 17.1000 23.4000 17.2000 ;
	    RECT 22.2000 16.8000 23.4000 17.1000 ;
	    RECT 31.0000 17.1000 31.4000 17.2000 ;
	    RECT 31.8000 17.1000 32.2000 17.2000 ;
	    RECT 31.0000 16.8000 32.2000 17.1000 ;
	    RECT 100.6000 16.8000 101.0000 17.2000 ;
	    RECT 18.2000 14.8000 18.6000 15.2000 ;
	    RECT 23.8000 15.1000 24.2000 15.2000 ;
	    RECT 24.6000 15.1000 25.0000 15.2000 ;
	    RECT 23.8000 14.8000 25.0000 15.1000 ;
	    RECT 35.8000 15.1000 36.2000 15.2000 ;
	    RECT 36.6000 15.1000 37.0000 15.2000 ;
	    RECT 35.8000 14.8000 37.0000 15.1000 ;
	    RECT 100.6000 12.2000 100.9000 16.8000 ;
	    RECT 100.6000 11.8000 101.0000 12.2000 ;
	    RECT 34.2000 10.8000 34.6000 11.2000 ;
	    RECT 34.2000 5.2000 34.5000 10.8000 ;
	    RECT 108.6000 7.2000 108.9000 26.8000 ;
	    RECT 125.4000 26.2000 125.7000 32.8000 ;
	    RECT 142.2000 32.2000 142.5000 39.8000 ;
	    RECT 150.2000 35.2000 150.5000 44.8000 ;
	    RECT 152.6000 41.2000 152.9000 73.8000 ;
	    RECT 158.2000 69.2000 158.5000 86.8000 ;
	    RECT 158.2000 68.8000 158.6000 69.2000 ;
	    RECT 159.0000 66.8000 159.4000 67.2000 ;
	    RECT 152.6000 40.8000 153.0000 41.2000 ;
	    RECT 150.2000 34.8000 150.6000 35.2000 ;
	    RECT 159.0000 34.2000 159.3000 66.8000 ;
	    RECT 159.0000 33.8000 159.4000 34.2000 ;
	    RECT 142.2000 31.8000 142.6000 32.2000 ;
	    RECT 125.4000 25.8000 125.8000 26.2000 ;
	    RECT 151.0000 24.8000 151.4000 25.2000 ;
	    RECT 115.8000 21.8000 116.2000 22.2000 ;
	    RECT 115.8000 13.2000 116.1000 21.8000 ;
	    RECT 136.6000 15.8000 137.0000 16.2000 ;
	    RECT 115.8000 12.8000 116.2000 13.2000 ;
	    RECT 136.6000 13.1000 136.9000 15.8000 ;
	    RECT 151.0000 15.2000 151.3000 24.8000 ;
	    RECT 153.4000 15.8000 153.8000 16.2000 ;
	    RECT 135.8000 12.8000 136.9000 13.1000 ;
	    RECT 140.6000 14.8000 141.0000 15.2000 ;
	    RECT 151.0000 14.8000 151.4000 15.2000 ;
	    RECT 135.8000 11.2000 136.1000 12.8000 ;
	    RECT 140.6000 11.2000 140.9000 14.8000 ;
	    RECT 153.4000 11.2000 153.7000 15.8000 ;
	    RECT 135.8000 10.8000 136.2000 11.2000 ;
	    RECT 140.6000 10.8000 141.0000 11.2000 ;
	    RECT 153.4000 10.8000 153.8000 11.2000 ;
	    RECT 160.6000 8.2000 160.9000 113.8000 ;
	    RECT 163.0000 106.1000 163.4000 106.2000 ;
	    RECT 163.8000 106.1000 164.2000 106.2000 ;
	    RECT 163.0000 105.8000 164.2000 106.1000 ;
	    RECT 163.0000 92.8000 163.4000 93.2000 ;
	    RECT 163.0000 54.2000 163.3000 92.8000 ;
	    RECT 164.6000 55.1000 164.9000 142.8000 ;
	    RECT 165.4000 132.2000 165.7000 146.8000 ;
	    RECT 166.2000 145.8000 166.6000 146.2000 ;
	    RECT 166.2000 145.2000 166.5000 145.8000 ;
	    RECT 166.2000 144.8000 166.6000 145.2000 ;
	    RECT 166.2000 137.8000 166.6000 138.2000 ;
	    RECT 165.4000 131.8000 165.8000 132.2000 ;
	    RECT 165.4000 130.8000 165.8000 131.2000 ;
	    RECT 165.4000 86.2000 165.7000 130.8000 ;
	    RECT 166.2000 126.2000 166.5000 137.8000 ;
	    RECT 171.8000 135.8000 172.2000 136.2000 ;
	    RECT 167.0000 132.8000 167.4000 133.2000 ;
	    RECT 167.0000 129.2000 167.3000 132.8000 ;
	    RECT 167.0000 128.8000 167.4000 129.2000 ;
	    RECT 166.2000 125.8000 166.6000 126.2000 ;
	    RECT 167.0000 98.2000 167.3000 128.8000 ;
	    RECT 167.0000 98.1000 167.4000 98.2000 ;
	    RECT 167.0000 97.8000 168.1000 98.1000 ;
	    RECT 165.4000 85.8000 165.8000 86.2000 ;
	    RECT 165.4000 55.1000 165.8000 55.2000 ;
	    RECT 164.6000 54.8000 165.8000 55.1000 ;
	    RECT 163.0000 53.8000 163.4000 54.2000 ;
	    RECT 162.2000 43.8000 162.6000 44.2000 ;
	    RECT 162.2000 40.2000 162.5000 43.8000 ;
	    RECT 162.2000 39.8000 162.6000 40.2000 ;
	    RECT 162.2000 38.8000 162.6000 39.2000 ;
	    RECT 161.4000 36.8000 161.8000 37.2000 ;
	    RECT 161.4000 36.2000 161.7000 36.8000 ;
	    RECT 161.4000 35.8000 161.8000 36.2000 ;
	    RECT 162.2000 35.2000 162.5000 38.8000 ;
	    RECT 163.0000 37.2000 163.3000 53.8000 ;
	    RECT 163.0000 36.8000 163.4000 37.2000 ;
	    RECT 167.0000 36.8000 167.4000 37.2000 ;
	    RECT 163.0000 36.1000 163.4000 36.2000 ;
	    RECT 163.8000 36.1000 164.2000 36.2000 ;
	    RECT 163.0000 35.8000 164.2000 36.1000 ;
	    RECT 162.2000 34.8000 162.6000 35.2000 ;
	    RECT 162.2000 15.1000 162.6000 15.2000 ;
	    RECT 163.0000 15.1000 163.4000 15.2000 ;
	    RECT 162.2000 14.8000 163.4000 15.1000 ;
	    RECT 160.6000 7.8000 161.0000 8.2000 ;
	    RECT 167.0000 7.2000 167.3000 36.8000 ;
	    RECT 167.8000 12.2000 168.1000 97.8000 ;
	    RECT 171.8000 93.2000 172.1000 135.8000 ;
	    RECT 171.8000 92.8000 172.2000 93.2000 ;
	    RECT 170.2000 88.8000 170.6000 89.2000 ;
	    RECT 168.6000 53.8000 169.0000 54.2000 ;
	    RECT 168.6000 29.1000 168.9000 53.8000 ;
	    RECT 169.4000 29.1000 169.8000 29.2000 ;
	    RECT 168.6000 28.8000 169.8000 29.1000 ;
	    RECT 167.8000 11.8000 168.2000 12.2000 ;
	    RECT 170.2000 7.2000 170.5000 88.8000 ;
	    RECT 43.8000 6.8000 44.2000 7.2000 ;
	    RECT 108.6000 6.8000 109.0000 7.2000 ;
	    RECT 167.0000 6.8000 167.4000 7.2000 ;
	    RECT 170.2000 6.8000 170.6000 7.2000 ;
	    RECT 43.8000 5.2000 44.1000 6.8000 ;
	    RECT 34.2000 4.8000 34.6000 5.2000 ;
	    RECT 43.8000 4.8000 44.2000 5.2000 ;
         LAYER metal5 ;
	    RECT 37.4000 154.1000 37.8000 154.2000 ;
	    RECT 47.0000 154.1000 47.4000 154.2000 ;
	    RECT 37.4000 153.8000 47.4000 154.1000 ;
	    RECT 131.0000 154.1000 131.4000 154.2000 ;
	    RECT 142.2000 154.1000 142.6000 154.2000 ;
	    RECT 131.0000 153.8000 142.6000 154.1000 ;
	    RECT 97.4000 152.1000 97.8000 152.2000 ;
	    RECT 104.6000 152.1000 105.0000 152.2000 ;
	    RECT 97.4000 151.8000 105.0000 152.1000 ;
	    RECT 166.2000 145.8000 166.6000 146.2000 ;
	    RECT 166.2000 145.3000 166.5000 145.8000 ;
	    RECT 166.1000 144.7000 166.7000 145.3000 ;
	    RECT 54.2000 136.1000 54.6000 136.2000 ;
	    RECT 56.6000 136.1000 57.0000 136.2000 ;
	    RECT 54.2000 135.8000 57.0000 136.1000 ;
	    RECT 96.6000 135.1000 97.0000 135.2000 ;
	    RECT 115.0000 135.1000 115.4000 135.2000 ;
	    RECT 96.6000 134.8000 115.4000 135.1000 ;
	    RECT 121.4000 134.1000 121.8000 134.2000 ;
	    RECT 132.6000 134.1000 133.0000 134.2000 ;
	    RECT 121.4000 133.8000 133.0000 134.1000 ;
	    RECT 165.4000 131.1000 165.8000 131.2000 ;
	    RECT 166.1000 131.1000 166.7000 131.3000 ;
	    RECT 165.4000 130.8000 166.7000 131.1000 ;
	    RECT 166.1000 130.7000 166.7000 130.8000 ;
	    RECT 110.2000 127.1000 110.6000 127.2000 ;
	    RECT 113.4000 127.1000 113.8000 127.2000 ;
	    RECT 110.2000 126.8000 113.8000 127.1000 ;
	    RECT 67.8000 107.1000 68.2000 107.2000 ;
	    RECT 80.6000 107.1000 81.0000 107.2000 ;
	    RECT 67.8000 106.8000 81.0000 107.1000 ;
	    RECT 19.8000 106.1000 20.2000 106.2000 ;
	    RECT 39.0000 106.1000 39.4000 106.2000 ;
	    RECT 19.8000 105.8000 39.4000 106.1000 ;
	    RECT 115.8000 106.1000 116.2000 106.2000 ;
	    RECT 163.0000 106.1000 163.4000 106.2000 ;
	    RECT 115.8000 105.8000 163.4000 106.1000 ;
	    RECT 58.2000 104.1000 58.6000 104.2000 ;
	    RECT 84.6000 104.1000 85.0000 104.2000 ;
	    RECT 58.2000 103.8000 85.0000 104.1000 ;
	    RECT 30.2000 95.1000 30.6000 95.2000 ;
	    RECT 36.6000 95.1000 37.0000 95.2000 ;
	    RECT 30.2000 94.8000 37.0000 95.1000 ;
	    RECT 57.4000 95.1000 57.8000 95.2000 ;
	    RECT 99.0000 95.1000 99.4000 95.2000 ;
	    RECT 57.4000 94.8000 99.4000 95.1000 ;
	    RECT 43.0000 94.1000 43.4000 94.2000 ;
	    RECT 105.4000 94.1000 105.8000 94.2000 ;
	    RECT 43.0000 93.8000 105.8000 94.1000 ;
	    RECT 19.8000 87.1000 20.2000 87.2000 ;
	    RECT 30.2000 87.1000 30.6000 87.2000 ;
	    RECT 19.8000 86.8000 30.6000 87.1000 ;
	    RECT 67.0000 87.1000 67.4000 87.2000 ;
	    RECT 100.6000 87.1000 101.0000 87.2000 ;
	    RECT 67.0000 86.8000 101.0000 87.1000 ;
	    RECT 22.2000 86.1000 22.6000 86.2000 ;
	    RECT 25.4000 86.1000 25.8000 86.2000 ;
	    RECT 22.2000 85.8000 25.8000 86.1000 ;
	    RECT 32.6000 86.1000 33.0000 86.2000 ;
	    RECT 34.2000 86.1000 34.6000 86.2000 ;
	    RECT 32.6000 85.8000 34.6000 86.1000 ;
	    RECT 75.8000 86.1000 76.2000 86.2000 ;
	    RECT 95.8000 86.1000 96.2000 86.2000 ;
	    RECT 75.8000 85.8000 96.2000 86.1000 ;
	    RECT 24.6000 85.1000 25.0000 85.2000 ;
	    RECT 43.8000 85.1000 44.2000 85.2000 ;
	    RECT 24.6000 84.8000 44.2000 85.1000 ;
	    RECT 64.6000 85.1000 65.0000 85.2000 ;
	    RECT 79.0000 85.1000 79.4000 85.2000 ;
	    RECT 64.6000 84.8000 79.4000 85.1000 ;
	    RECT 69.4000 77.1000 69.8000 77.2000 ;
	    RECT 93.4000 77.1000 93.8000 77.2000 ;
	    RECT 69.4000 76.8000 93.8000 77.1000 ;
	    RECT 45.4000 59.1000 45.8000 59.2000 ;
	    RECT 62.2000 59.1000 62.6000 59.2000 ;
	    RECT 45.4000 58.8000 62.6000 59.1000 ;
	    RECT 13.4000 57.1000 13.8000 57.2000 ;
	    RECT 42.2000 57.1000 42.6000 57.2000 ;
	    RECT 13.4000 56.8000 42.6000 57.1000 ;
	    RECT 37.4000 56.1000 37.8000 56.2000 ;
	    RECT 63.8000 56.1000 64.2000 56.2000 ;
	    RECT 37.4000 55.8000 64.2000 56.1000 ;
	    RECT 15.8000 55.1000 16.2000 55.2000 ;
	    RECT 38.2000 55.1000 38.6000 55.2000 ;
	    RECT 15.8000 54.8000 38.6000 55.1000 ;
	    RECT 28.6000 47.1000 29.0000 47.2000 ;
	    RECT 90.2000 47.1000 90.6000 47.2000 ;
	    RECT 28.6000 46.8000 90.6000 47.1000 ;
	    RECT 51.8000 43.1000 52.2000 43.2000 ;
	    RECT 60.6000 43.1000 61.0000 43.2000 ;
	    RECT 51.8000 42.8000 61.0000 43.1000 ;
	    RECT 163.0000 37.1000 163.4000 37.2000 ;
	    RECT 167.0000 37.1000 167.4000 37.2000 ;
	    RECT 163.0000 36.8000 167.4000 37.1000 ;
	    RECT 22.2000 36.1000 22.6000 36.2000 ;
	    RECT 26.2000 36.1000 26.6000 36.2000 ;
	    RECT 22.2000 35.8000 26.6000 36.1000 ;
	    RECT 161.4000 36.1000 161.8000 36.2000 ;
	    RECT 163.0000 36.1000 163.4000 36.2000 ;
	    RECT 161.4000 35.8000 163.4000 36.1000 ;
	    RECT 23.8000 35.1000 24.2000 35.2000 ;
	    RECT 29.4000 35.1000 29.8000 35.2000 ;
	    RECT 23.8000 34.8000 29.8000 35.1000 ;
	    RECT 57.4000 34.1000 57.8000 34.2000 ;
	    RECT 75.8000 34.1000 76.2000 34.2000 ;
	    RECT 57.4000 33.8000 76.2000 34.1000 ;
	    RECT 98.2000 34.1000 98.6000 34.2000 ;
	    RECT 103.8000 34.1000 104.2000 34.2000 ;
	    RECT 98.2000 33.8000 104.2000 34.1000 ;
	    RECT 110.2000 29.1000 110.6000 29.2000 ;
	    RECT 117.4000 29.1000 117.8000 29.2000 ;
	    RECT 110.2000 28.8000 117.8000 29.1000 ;
	    RECT 14.2000 24.1000 14.6000 24.2000 ;
	    RECT 24.6000 24.1000 25.0000 24.2000 ;
	    RECT 14.2000 23.8000 25.0000 24.1000 ;
	    RECT 22.2000 17.1000 22.6000 17.2000 ;
	    RECT 31.0000 17.1000 31.4000 17.2000 ;
	    RECT 22.2000 16.8000 31.4000 17.1000 ;
	    RECT 24.6000 15.1000 25.0000 15.2000 ;
	    RECT 35.8000 15.1000 36.2000 15.2000 ;
	    RECT 24.6000 14.8000 36.2000 15.1000 ;
	    RECT 140.6000 15.1000 141.0000 15.2000 ;
	    RECT 163.0000 15.1000 163.4000 15.2000 ;
	    RECT 140.6000 14.8000 163.4000 15.1000 ;
         LAYER metal6 ;
	    RECT 166.1000 144.7000 166.7000 145.3000 ;
	    RECT 166.1000 131.3000 166.6000 144.7000 ;
	    RECT 166.1000 130.7000 166.7000 131.3000 ;
   END
END nibble_top
