magic
tech scmos
timestamp 1559787497
<< metal1 >>
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 485 1403 488 1407
rect 362 1368 363 1372
rect 1062 1366 1066 1368
rect 1174 1366 1178 1368
rect 70 1358 89 1361
rect 94 1358 105 1361
rect 158 1358 169 1361
rect 394 1358 409 1361
rect 414 1358 422 1361
rect 490 1358 505 1361
rect 94 1352 97 1358
rect 274 1348 289 1351
rect 442 1348 457 1351
rect 466 1348 497 1351
rect 14 1338 25 1341
rect 302 1338 321 1341
rect 334 1338 342 1341
rect 382 1338 390 1341
rect 494 1338 497 1348
rect 606 1351 609 1361
rect 590 1348 609 1351
rect 622 1351 625 1358
rect 622 1348 641 1351
rect 766 1351 769 1361
rect 854 1358 865 1361
rect 766 1348 785 1351
rect 974 1351 977 1361
rect 1118 1352 1121 1361
rect 1126 1358 1145 1361
rect 1154 1358 1158 1362
rect 1190 1361 1193 1368
rect 1358 1366 1362 1368
rect 1182 1358 1193 1361
rect 1238 1358 1249 1361
rect 1266 1358 1273 1361
rect 1374 1361 1377 1368
rect 1366 1358 1377 1361
rect 974 1348 1009 1351
rect 1066 1348 1073 1351
rect 1078 1348 1094 1351
rect 1158 1348 1174 1351
rect 1190 1348 1206 1351
rect 1214 1348 1230 1351
rect 1350 1348 1361 1351
rect 510 1341 513 1348
rect 510 1338 521 1341
rect 566 1338 577 1341
rect 678 1341 681 1348
rect 670 1338 681 1341
rect 734 1338 745 1341
rect 906 1338 913 1341
rect 942 1338 953 1341
rect 1018 1338 1025 1341
rect 1078 1338 1081 1348
rect 1110 1338 1118 1341
rect 1190 1338 1193 1348
rect 1358 1342 1361 1348
rect 1374 1348 1390 1351
rect 1414 1351 1417 1361
rect 1398 1348 1417 1351
rect 1334 1338 1342 1341
rect 1374 1338 1377 1348
rect 1430 1338 1438 1341
rect 1046 1328 1049 1338
rect 130 1318 131 1322
rect 429 1318 430 1322
rect 613 1318 614 1322
rect 690 1318 691 1322
rect 805 1318 806 1322
rect 829 1318 830 1322
rect 869 1318 870 1322
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 966 1288 974 1291
rect 958 1272 961 1281
rect 206 1268 214 1271
rect 334 1268 350 1271
rect 398 1268 409 1271
rect 710 1268 721 1271
rect 758 1268 769 1271
rect 790 1268 801 1271
rect 1062 1271 1065 1278
rect 978 1268 993 1271
rect 1054 1268 1065 1271
rect 1098 1268 1105 1271
rect 1204 1268 1206 1272
rect 238 1258 249 1261
rect 314 1258 321 1261
rect 950 1258 958 1261
rect 978 1258 1001 1261
rect 238 1252 241 1258
rect 302 1248 310 1251
rect 358 1248 369 1251
rect 374 1248 382 1251
rect 462 1248 470 1251
rect 662 1248 673 1251
rect 730 1248 737 1251
rect 1238 1248 1246 1251
rect 1422 1248 1433 1251
rect 650 1238 657 1241
rect 1054 1241 1057 1248
rect 1422 1242 1425 1248
rect 898 1238 905 1241
rect 1046 1238 1057 1241
rect 1454 1241 1458 1244
rect 1454 1238 1462 1241
rect 1142 1228 1145 1238
rect 1318 1228 1321 1238
rect 418 1218 419 1222
rect 749 1218 750 1222
rect 810 1218 811 1222
rect 1002 1218 1003 1222
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 485 1203 488 1207
rect 378 1168 393 1171
rect 966 1168 974 1171
rect 1158 1168 1169 1171
rect 1250 1168 1257 1171
rect 1294 1168 1310 1171
rect 182 1158 190 1161
rect 350 1161 353 1168
rect 1158 1162 1161 1168
rect 334 1158 345 1161
rect 350 1158 361 1161
rect 494 1158 505 1161
rect 522 1158 529 1161
rect 566 1158 577 1161
rect 758 1158 777 1161
rect 878 1158 886 1161
rect 990 1158 1017 1161
rect 1062 1158 1073 1161
rect 1174 1158 1185 1161
rect 1202 1158 1209 1161
rect 1294 1158 1297 1168
rect 678 1151 681 1158
rect 670 1148 681 1151
rect 62 1138 65 1148
rect 1150 1138 1161 1141
rect 1278 1138 1289 1141
rect 1438 1141 1441 1148
rect 1430 1138 1441 1141
rect 430 1128 433 1138
rect 1150 1132 1153 1138
rect 1286 1132 1289 1138
rect 1442 1128 1446 1132
rect 38 1118 46 1121
rect 94 1118 102 1121
rect 204 1118 206 1122
rect 330 1118 331 1122
rect 509 1118 510 1122
rect 533 1118 534 1122
rect 636 1118 638 1122
rect 690 1118 691 1122
rect 781 1118 782 1122
rect 858 1118 860 1122
rect 898 1118 905 1121
rect 1077 1118 1078 1122
rect 1106 1118 1113 1121
rect 1314 1118 1321 1121
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 730 1088 731 1092
rect 966 1088 974 1091
rect 466 1078 481 1081
rect 978 1078 993 1081
rect 22 1074 26 1078
rect 198 1068 209 1071
rect 342 1071 345 1078
rect 342 1068 350 1071
rect 710 1068 721 1071
rect 1142 1071 1145 1078
rect 1190 1072 1193 1081
rect 1142 1068 1153 1071
rect 1398 1068 1406 1071
rect 198 1062 201 1068
rect 182 1058 193 1061
rect 226 1058 233 1061
rect 182 1052 185 1058
rect 126 1048 134 1051
rect 366 1048 377 1051
rect 398 1048 409 1051
rect 454 1048 470 1051
rect 734 1048 745 1051
rect 850 1048 857 1051
rect 1074 1048 1081 1051
rect 1166 1048 1185 1051
rect 1198 1048 1209 1051
rect 422 1041 425 1048
rect 414 1038 425 1041
rect 1034 1038 1041 1041
rect 1062 1038 1078 1041
rect 1150 1041 1153 1048
rect 1150 1038 1161 1041
rect 1246 1041 1249 1061
rect 1286 1056 1290 1058
rect 1246 1038 1265 1041
rect 294 1028 297 1038
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 485 1003 488 1007
rect 246 972 249 981
rect 718 971 721 981
rect 718 968 753 971
rect 1166 968 1177 971
rect 1350 971 1353 981
rect 1318 968 1353 971
rect 1430 968 1438 971
rect 234 958 241 961
rect 662 961 665 968
rect 1174 962 1177 968
rect 654 958 665 961
rect 722 958 729 961
rect 1078 958 1089 961
rect 1110 958 1121 961
rect 1142 958 1161 961
rect 1278 958 1289 961
rect 1414 958 1425 961
rect 30 951 34 953
rect 22 948 34 951
rect 174 942 177 951
rect 474 948 481 951
rect 986 948 1009 951
rect 1238 948 1246 951
rect 190 938 198 941
rect 566 938 574 941
rect 666 938 673 941
rect 1218 938 1225 941
rect 1438 938 1446 941
rect 566 928 569 938
rect 670 928 673 938
rect 958 928 969 931
rect 214 918 222 921
rect 606 918 614 921
rect 746 918 753 921
rect 882 918 889 921
rect 1042 918 1049 921
rect 1293 918 1294 922
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 290 888 297 891
rect 394 888 395 892
rect 418 888 419 892
rect 470 871 473 881
rect 526 872 529 881
rect 470 868 494 871
rect 678 871 682 872
rect 686 871 689 878
rect 678 868 689 871
rect 934 871 937 878
rect 934 868 945 871
rect 1110 868 1121 871
rect 1206 871 1209 878
rect 1206 868 1217 871
rect 1438 868 1478 871
rect 22 858 34 861
rect 62 858 70 861
rect 174 858 186 861
rect 1110 862 1113 868
rect 598 858 609 861
rect 30 857 34 858
rect 182 857 186 858
rect 358 851 361 858
rect 598 852 601 858
rect 358 848 369 851
rect 510 848 521 851
rect 614 848 625 851
rect 690 848 697 851
rect 710 848 721 851
rect 814 848 825 851
rect 942 851 945 858
rect 942 848 953 851
rect 958 848 969 851
rect 1230 848 1249 851
rect 1262 848 1273 851
rect 350 838 358 841
rect 726 838 734 841
rect 838 841 841 848
rect 838 838 849 841
rect 1214 841 1217 848
rect 1286 841 1289 848
rect 1214 838 1225 841
rect 1278 838 1289 841
rect 994 828 1001 831
rect 472 803 474 807
rect 478 803 481 807
rect 485 803 488 807
rect 74 768 77 772
rect 898 768 905 771
rect 1006 771 1009 781
rect 986 768 1009 771
rect 470 758 497 761
rect 54 752 58 753
rect 302 751 306 753
rect 294 748 306 751
rect 550 748 558 751
rect 1414 751 1418 753
rect 1414 748 1425 751
rect 636 738 638 742
rect 826 738 828 742
rect 958 738 972 741
rect 422 728 430 731
rect 614 731 617 738
rect 606 728 617 731
rect 718 731 721 738
rect 958 732 961 738
rect 718 728 729 731
rect 501 718 502 722
rect 670 718 678 721
rect 866 718 873 721
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 430 688 438 691
rect 954 688 955 692
rect 614 681 617 688
rect 606 678 617 681
rect 794 678 801 681
rect 874 678 881 681
rect 38 668 46 671
rect 226 668 233 671
rect 462 671 465 678
rect 926 672 929 681
rect 462 668 476 671
rect 882 668 889 671
rect 994 668 1002 671
rect 1254 668 1262 671
rect 870 658 873 668
rect 1182 658 1193 661
rect 1286 658 1289 668
rect 1414 658 1425 661
rect 1462 658 1470 661
rect 38 651 41 658
rect 1182 657 1186 658
rect 1414 657 1418 658
rect 6 648 25 651
rect 30 648 41 651
rect 206 648 217 651
rect 258 648 265 651
rect 382 648 401 651
rect 710 648 721 651
rect 958 648 977 651
rect 398 642 401 648
rect 194 638 201 641
rect 350 638 358 641
rect 430 638 446 641
rect 458 638 473 641
rect 518 628 521 638
rect 472 603 474 607
rect 478 603 481 607
rect 485 603 488 607
rect 298 588 299 592
rect 98 568 118 571
rect 170 568 193 571
rect 254 568 262 571
rect 582 568 609 571
rect 718 568 729 571
rect 1110 568 1118 571
rect 1206 568 1217 571
rect 718 562 721 568
rect 1214 562 1217 568
rect 14 558 25 561
rect 238 558 249 561
rect 466 558 473 561
rect 554 558 561 561
rect 734 558 745 561
rect 766 558 777 561
rect 926 558 937 561
rect 982 558 990 561
rect 1182 558 1201 561
rect 30 548 38 551
rect 1342 542 1345 551
rect 38 538 49 541
rect 278 538 289 541
rect 374 538 393 541
rect 710 538 721 541
rect 1042 538 1049 541
rect 46 532 49 538
rect 374 532 377 538
rect 710 532 713 538
rect 974 528 977 538
rect 1002 528 1009 531
rect 1342 528 1350 531
rect 146 518 148 522
rect 781 518 782 522
rect 922 518 923 522
rect 957 518 958 522
rect 1133 518 1134 522
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 85 488 86 492
rect 210 488 217 491
rect 434 488 435 492
rect 453 488 454 492
rect 525 488 526 492
rect 581 488 582 492
rect 634 488 635 492
rect 706 488 707 492
rect 810 488 812 492
rect 1306 488 1313 491
rect 994 478 1009 481
rect 14 468 25 471
rect 282 468 297 471
rect 482 468 489 471
rect 846 471 849 478
rect 854 471 858 472
rect 846 468 858 471
rect 1014 468 1025 471
rect 1022 462 1025 468
rect 38 458 46 461
rect 414 458 422 461
rect 594 458 601 461
rect 1038 461 1041 471
rect 1070 468 1078 471
rect 1114 468 1121 471
rect 1164 468 1177 471
rect 1270 471 1274 472
rect 1278 471 1281 478
rect 1270 468 1281 471
rect 1174 462 1177 468
rect 1038 458 1046 461
rect 1050 458 1057 461
rect 1334 458 1342 461
rect 46 448 65 451
rect 838 448 846 451
rect 978 448 1006 451
rect 1030 448 1041 451
rect 294 441 297 448
rect 1022 442 1026 444
rect 294 438 305 441
rect 682 438 689 441
rect 1038 442 1041 448
rect 1190 441 1193 448
rect 1182 438 1193 441
rect 1438 418 1446 421
rect 472 403 474 407
rect 478 403 481 407
rect 485 403 488 407
rect 222 368 230 371
rect 318 368 329 371
rect 814 371 817 381
rect 814 368 849 371
rect 926 371 929 381
rect 926 368 961 371
rect 1078 368 1089 371
rect 1370 368 1377 371
rect 1430 371 1433 381
rect 1410 368 1433 371
rect 94 361 97 368
rect 318 362 321 368
rect 86 358 97 361
rect 230 358 238 361
rect 350 361 353 368
rect 334 358 345 361
rect 350 358 361 361
rect 422 358 433 361
rect 510 361 513 368
rect 502 358 513 361
rect 666 358 673 361
rect 702 358 710 361
rect 790 361 793 368
rect 1078 362 1081 368
rect 782 358 793 361
rect 1010 358 1017 361
rect 1094 358 1105 361
rect 230 352 234 354
rect 694 348 702 351
rect 1122 348 1129 351
rect 726 341 729 348
rect 726 338 737 341
rect 746 338 753 341
rect 862 338 865 348
rect 950 338 962 341
rect 1066 338 1078 341
rect 1162 338 1169 341
rect 1298 338 1305 341
rect 1462 338 1470 341
rect 950 332 953 338
rect 1150 328 1161 331
rect 306 318 307 322
rect 1394 318 1396 322
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 118 288 126 291
rect 146 288 148 292
rect 186 288 193 291
rect 250 288 251 292
rect 402 288 403 292
rect 478 288 486 291
rect 597 288 598 292
rect 842 288 849 291
rect 1125 288 1126 292
rect 1354 288 1361 291
rect 270 281 273 288
rect 270 278 281 281
rect 1446 278 1470 281
rect 322 268 329 271
rect 342 268 358 271
rect 362 268 369 271
rect 410 268 417 271
rect 606 268 614 271
rect 942 268 953 271
rect 942 262 945 268
rect 430 258 438 261
rect 1046 258 1057 261
rect 14 248 25 251
rect 170 248 177 251
rect 478 248 505 251
rect 646 251 649 258
rect 1046 252 1049 258
rect 582 248 593 251
rect 638 248 649 251
rect 662 248 673 251
rect 822 248 830 251
rect 934 248 945 251
rect 962 248 969 251
rect 1022 248 1033 251
rect 1090 248 1097 251
rect 1286 248 1294 251
rect 1390 248 1401 251
rect 1430 248 1441 251
rect 38 241 41 248
rect 30 238 41 241
rect 218 238 225 241
rect 230 238 238 241
rect 1038 238 1046 241
rect 1226 238 1241 241
rect 1334 238 1342 241
rect 702 228 705 238
rect 902 228 905 238
rect 974 228 977 238
rect 472 203 474 207
rect 478 203 481 207
rect 485 203 488 207
rect 317 188 318 192
rect 365 188 366 192
rect 506 188 507 192
rect 1102 168 1113 171
rect 1214 168 1222 171
rect 1438 168 1470 171
rect 1110 162 1113 168
rect 654 158 673 161
rect 1010 158 1017 161
rect 1086 158 1097 161
rect 1230 158 1238 161
rect 366 148 374 151
rect 414 148 422 151
rect 498 148 505 151
rect 1198 151 1201 158
rect 1190 148 1201 151
rect 206 138 217 141
rect 374 138 385 141
rect 470 138 497 141
rect 582 138 593 141
rect 614 138 622 141
rect 1114 138 1121 141
rect 206 132 209 138
rect 22 128 30 131
rect 702 128 713 131
rect 822 128 833 131
rect 990 128 998 131
rect 1118 128 1121 138
rect 710 122 713 128
rect 830 122 833 128
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 138 88 139 92
rect 218 88 219 92
rect 314 88 315 92
rect 349 88 350 92
rect 478 88 486 91
rect 938 88 939 92
rect 1213 88 1214 92
rect 1238 88 1246 91
rect 622 72 625 81
rect 1458 78 1478 81
rect 62 58 81 61
rect 102 61 105 71
rect 122 68 129 71
rect 90 58 105 61
rect 242 58 257 61
rect 278 61 281 71
rect 298 68 305 71
rect 318 68 329 71
rect 358 68 366 71
rect 374 68 385 71
rect 458 68 465 71
rect 550 68 561 71
rect 590 68 598 71
rect 630 68 641 71
rect 678 68 689 71
rect 734 68 742 71
rect 758 68 766 71
rect 878 68 889 71
rect 1014 68 1025 71
rect 1070 68 1081 71
rect 266 58 281 61
rect 318 62 321 68
rect 1078 62 1081 68
rect 406 58 425 61
rect 542 58 550 61
rect 710 58 729 61
rect 846 58 865 61
rect 986 58 1001 61
rect 1086 58 1094 61
rect 14 48 25 51
rect 62 48 65 58
rect 102 48 113 51
rect 182 48 193 51
rect 222 48 233 51
rect 278 48 289 51
rect 406 48 409 58
rect 478 48 502 51
rect 510 48 529 51
rect 566 48 577 51
rect 582 48 590 51
rect 662 48 665 58
rect 710 48 713 58
rect 790 48 809 51
rect 846 48 849 58
rect 902 51 905 58
rect 902 48 913 51
rect 942 48 953 51
rect 974 48 982 51
rect 1038 48 1049 51
rect 1250 48 1257 51
rect 1354 48 1361 51
rect 102 42 105 48
rect 278 42 281 48
rect 502 41 506 44
rect 498 38 506 41
rect 566 42 569 48
rect 614 41 618 44
rect 622 41 625 48
rect 614 38 625 41
rect 1078 42 1082 44
rect 541 28 542 32
rect 472 3 474 7
rect 478 3 481 7
rect 485 3 488 7
<< m2contact >>
rect 474 1403 478 1407
rect 481 1403 485 1407
rect 358 1368 362 1372
rect 1062 1368 1066 1372
rect 1174 1368 1178 1372
rect 1190 1368 1194 1372
rect 1358 1368 1362 1372
rect 46 1358 50 1362
rect 110 1358 114 1362
rect 134 1358 138 1362
rect 206 1358 210 1362
rect 270 1358 274 1362
rect 278 1358 282 1362
rect 342 1358 346 1362
rect 374 1358 378 1362
rect 390 1358 394 1362
rect 422 1358 426 1362
rect 446 1358 450 1362
rect 486 1358 490 1362
rect 510 1358 514 1362
rect 598 1358 602 1362
rect 30 1348 34 1352
rect 94 1348 98 1352
rect 198 1348 202 1352
rect 230 1348 234 1352
rect 270 1348 274 1352
rect 294 1348 298 1352
rect 358 1348 362 1352
rect 438 1348 442 1352
rect 462 1348 466 1352
rect 54 1338 58 1342
rect 94 1338 98 1342
rect 118 1338 122 1342
rect 142 1338 146 1342
rect 182 1338 186 1342
rect 222 1338 226 1342
rect 246 1338 250 1342
rect 254 1338 258 1342
rect 326 1338 330 1342
rect 342 1338 346 1342
rect 350 1338 354 1342
rect 390 1338 394 1342
rect 398 1338 402 1342
rect 438 1338 442 1342
rect 470 1338 474 1342
rect 510 1348 514 1352
rect 550 1348 554 1352
rect 582 1348 586 1352
rect 622 1358 626 1362
rect 630 1358 634 1362
rect 694 1358 698 1362
rect 718 1358 722 1362
rect 654 1348 658 1352
rect 678 1348 682 1352
rect 750 1348 754 1352
rect 774 1358 778 1362
rect 798 1358 802 1362
rect 822 1358 826 1362
rect 902 1358 906 1362
rect 926 1348 930 1352
rect 958 1348 962 1352
rect 998 1358 1002 1362
rect 1038 1358 1042 1362
rect 1110 1358 1114 1362
rect 1158 1358 1162 1362
rect 1374 1368 1378 1372
rect 1222 1358 1226 1362
rect 1262 1358 1266 1362
rect 1294 1358 1298 1362
rect 1318 1358 1322 1362
rect 1406 1358 1410 1362
rect 1062 1348 1066 1352
rect 1094 1348 1098 1352
rect 1118 1348 1122 1352
rect 1174 1348 1178 1352
rect 1206 1348 1210 1352
rect 1230 1348 1234 1352
rect 622 1338 626 1342
rect 646 1338 650 1342
rect 702 1338 706 1342
rect 766 1338 770 1342
rect 790 1338 794 1342
rect 814 1338 818 1342
rect 838 1338 842 1342
rect 878 1338 882 1342
rect 886 1338 890 1342
rect 902 1338 906 1342
rect 966 1338 970 1342
rect 1014 1338 1018 1342
rect 1046 1338 1050 1342
rect 1086 1338 1090 1342
rect 1118 1338 1122 1342
rect 1134 1338 1138 1342
rect 1166 1338 1170 1342
rect 1390 1348 1394 1352
rect 1438 1358 1442 1362
rect 1198 1338 1202 1342
rect 1262 1338 1266 1342
rect 1286 1338 1290 1342
rect 1310 1338 1314 1342
rect 1342 1338 1346 1342
rect 1358 1338 1362 1342
rect 1382 1338 1386 1342
rect 1438 1338 1442 1342
rect 1454 1338 1458 1342
rect 6 1328 10 1332
rect 78 1328 82 1332
rect 174 1328 178 1332
rect 310 1328 314 1332
rect 390 1328 394 1332
rect 526 1328 530 1332
rect 558 1328 562 1332
rect 726 1328 730 1332
rect 846 1328 850 1332
rect 934 1328 938 1332
rect 1054 1328 1058 1332
rect 1230 1328 1234 1332
rect 1342 1328 1346 1332
rect 46 1318 50 1322
rect 70 1318 74 1322
rect 126 1318 130 1322
rect 158 1318 162 1322
rect 206 1318 210 1322
rect 270 1318 274 1322
rect 430 1318 434 1322
rect 534 1318 538 1322
rect 614 1318 618 1322
rect 686 1318 690 1322
rect 718 1318 722 1322
rect 806 1318 810 1322
rect 830 1318 834 1322
rect 870 1318 874 1322
rect 902 1318 906 1322
rect 1038 1318 1042 1322
rect 1246 1318 1250 1322
rect 1270 1318 1274 1322
rect 1294 1318 1298 1322
rect 1318 1318 1322 1322
rect 1414 1318 1418 1322
rect 1438 1318 1442 1322
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 222 1288 226 1292
rect 974 1288 978 1292
rect 1030 1288 1034 1292
rect 1158 1288 1162 1292
rect 30 1278 34 1282
rect 94 1278 98 1282
rect 214 1278 218 1282
rect 254 1278 258 1282
rect 342 1278 346 1282
rect 350 1278 354 1282
rect 390 1278 394 1282
rect 438 1278 442 1282
rect 518 1278 522 1282
rect 582 1278 586 1282
rect 678 1278 682 1282
rect 726 1278 730 1282
rect 774 1278 778 1282
rect 782 1278 786 1282
rect 830 1278 834 1282
rect 894 1278 898 1282
rect 910 1278 914 1282
rect 942 1278 946 1282
rect 1022 1278 1026 1282
rect 1062 1278 1066 1282
rect 1094 1278 1098 1282
rect 1366 1278 1370 1282
rect 6 1268 10 1272
rect 38 1268 42 1272
rect 102 1268 106 1272
rect 214 1268 218 1272
rect 238 1268 242 1272
rect 310 1268 314 1272
rect 350 1268 354 1272
rect 382 1268 386 1272
rect 446 1268 450 1272
rect 526 1268 530 1272
rect 590 1268 594 1272
rect 606 1268 610 1272
rect 646 1268 650 1272
rect 838 1268 842 1272
rect 918 1268 922 1272
rect 958 1268 962 1272
rect 974 1268 978 1272
rect 1070 1268 1074 1272
rect 1094 1268 1098 1272
rect 1206 1268 1210 1272
rect 1358 1268 1362 1272
rect 1438 1268 1442 1272
rect 54 1258 58 1262
rect 78 1258 82 1262
rect 118 1258 122 1262
rect 134 1258 138 1262
rect 174 1258 178 1262
rect 190 1258 194 1262
rect 270 1258 274 1262
rect 310 1258 314 1262
rect 414 1258 418 1262
rect 502 1258 506 1262
rect 542 1258 546 1262
rect 558 1258 562 1262
rect 622 1258 626 1262
rect 694 1258 698 1262
rect 702 1258 706 1262
rect 750 1258 754 1262
rect 806 1258 810 1262
rect 878 1258 882 1262
rect 958 1258 962 1262
rect 974 1258 978 1262
rect 1118 1258 1122 1262
rect 1142 1258 1146 1262
rect 1174 1258 1178 1262
rect 1190 1258 1194 1262
rect 1230 1258 1234 1262
rect 1254 1258 1258 1262
rect 1286 1258 1290 1262
rect 1318 1258 1322 1262
rect 1342 1258 1346 1262
rect 1382 1258 1386 1262
rect 1414 1258 1418 1262
rect 22 1248 26 1252
rect 86 1248 90 1252
rect 126 1248 130 1252
rect 182 1248 186 1252
rect 222 1248 226 1252
rect 238 1248 242 1252
rect 262 1248 266 1252
rect 294 1248 298 1252
rect 310 1248 314 1252
rect 382 1248 386 1252
rect 430 1248 434 1252
rect 470 1248 474 1252
rect 510 1248 514 1252
rect 574 1248 578 1252
rect 614 1248 618 1252
rect 686 1248 690 1252
rect 726 1248 730 1252
rect 822 1248 826 1252
rect 854 1248 858 1252
rect 886 1248 890 1252
rect 1014 1248 1018 1252
rect 1038 1248 1042 1252
rect 1054 1248 1058 1252
rect 1086 1248 1090 1252
rect 1150 1248 1154 1252
rect 1182 1248 1186 1252
rect 1246 1248 1250 1252
rect 1278 1248 1282 1252
rect 1310 1248 1314 1252
rect 1374 1248 1378 1252
rect 70 1238 74 1242
rect 142 1238 146 1242
rect 166 1238 170 1242
rect 278 1238 282 1242
rect 494 1238 498 1242
rect 558 1238 562 1242
rect 630 1238 634 1242
rect 646 1238 650 1242
rect 870 1238 874 1242
rect 894 1238 898 1242
rect 1134 1238 1138 1242
rect 1142 1238 1146 1242
rect 1198 1238 1202 1242
rect 1222 1238 1226 1242
rect 1262 1238 1266 1242
rect 1294 1238 1298 1242
rect 1318 1238 1322 1242
rect 1326 1238 1330 1242
rect 1390 1238 1394 1242
rect 1414 1238 1418 1242
rect 1422 1238 1426 1242
rect 1462 1238 1466 1242
rect 1406 1228 1410 1232
rect 1446 1228 1450 1232
rect 14 1218 18 1222
rect 78 1218 82 1222
rect 134 1218 138 1222
rect 174 1218 178 1222
rect 270 1218 274 1222
rect 414 1218 418 1222
rect 502 1218 506 1222
rect 566 1218 570 1222
rect 638 1218 642 1222
rect 750 1218 754 1222
rect 806 1218 810 1222
rect 878 1218 882 1222
rect 934 1218 938 1222
rect 998 1218 1002 1222
rect 1230 1218 1234 1222
rect 1270 1218 1274 1222
rect 1302 1218 1306 1222
rect 1382 1218 1386 1222
rect 474 1203 478 1207
rect 481 1203 485 1207
rect 70 1188 74 1192
rect 158 1188 162 1192
rect 230 1188 234 1192
rect 422 1188 426 1192
rect 558 1188 562 1192
rect 926 1188 930 1192
rect 1430 1188 1434 1192
rect 1462 1188 1466 1192
rect 710 1178 714 1182
rect 1238 1178 1242 1182
rect 1358 1178 1362 1182
rect 38 1168 42 1172
rect 94 1168 98 1172
rect 126 1168 130 1172
rect 166 1168 170 1172
rect 198 1168 202 1172
rect 270 1168 274 1172
rect 350 1168 354 1172
rect 366 1168 370 1172
rect 374 1168 378 1172
rect 630 1168 634 1172
rect 718 1168 722 1172
rect 862 1168 866 1172
rect 902 1168 906 1172
rect 934 1168 938 1172
rect 974 1168 978 1172
rect 982 1168 986 1172
rect 1110 1168 1114 1172
rect 1246 1168 1250 1172
rect 1278 1168 1282 1172
rect 1310 1168 1314 1172
rect 1318 1168 1322 1172
rect 1366 1168 1370 1172
rect 54 1158 58 1162
rect 110 1158 114 1162
rect 142 1158 146 1162
rect 150 1158 154 1162
rect 190 1158 194 1162
rect 254 1158 258 1162
rect 382 1158 386 1162
rect 518 1158 522 1162
rect 614 1158 618 1162
rect 678 1158 682 1162
rect 694 1158 698 1162
rect 702 1158 706 1162
rect 734 1158 738 1162
rect 830 1158 834 1162
rect 886 1158 890 1162
rect 918 1158 922 1162
rect 1030 1158 1034 1162
rect 1094 1158 1098 1162
rect 1126 1158 1130 1162
rect 1158 1158 1162 1162
rect 1198 1158 1202 1162
rect 1262 1158 1266 1162
rect 1302 1158 1306 1162
rect 1350 1158 1354 1162
rect 1438 1158 1442 1162
rect 22 1148 26 1152
rect 46 1148 50 1152
rect 62 1148 66 1152
rect 102 1148 106 1152
rect 134 1148 138 1152
rect 158 1148 162 1152
rect 190 1148 194 1152
rect 214 1148 218 1152
rect 262 1148 266 1152
rect 286 1148 290 1152
rect 374 1148 378 1152
rect 606 1148 610 1152
rect 622 1148 626 1152
rect 710 1148 714 1152
rect 870 1148 874 1152
rect 894 1148 898 1152
rect 926 1148 930 1152
rect 950 1148 954 1152
rect 1102 1148 1106 1152
rect 1286 1148 1290 1152
rect 1310 1148 1314 1152
rect 1358 1148 1362 1152
rect 1414 1148 1418 1152
rect 1438 1148 1442 1152
rect 6 1138 10 1142
rect 230 1138 234 1142
rect 246 1138 250 1142
rect 302 1138 306 1142
rect 318 1138 322 1142
rect 406 1138 410 1142
rect 430 1138 434 1142
rect 454 1138 458 1142
rect 518 1138 522 1142
rect 542 1138 546 1142
rect 550 1138 554 1142
rect 654 1138 658 1142
rect 678 1138 682 1142
rect 750 1138 754 1142
rect 790 1138 794 1142
rect 814 1138 818 1142
rect 846 1138 850 1142
rect 974 1138 978 1142
rect 1046 1138 1050 1142
rect 1086 1138 1090 1142
rect 1142 1138 1146 1142
rect 1222 1138 1226 1142
rect 1246 1138 1250 1142
rect 1342 1138 1346 1142
rect 1382 1138 1386 1142
rect 1398 1138 1402 1142
rect 1454 1138 1458 1142
rect 310 1128 314 1132
rect 350 1128 354 1132
rect 414 1128 418 1132
rect 462 1128 466 1132
rect 486 1128 490 1132
rect 582 1128 586 1132
rect 590 1128 594 1132
rect 646 1128 650 1132
rect 766 1128 770 1132
rect 822 1128 826 1132
rect 1022 1128 1026 1132
rect 1054 1128 1058 1132
rect 1150 1128 1154 1132
rect 1190 1128 1194 1132
rect 1198 1128 1202 1132
rect 1214 1128 1218 1132
rect 1286 1128 1290 1132
rect 1406 1128 1410 1132
rect 1438 1128 1442 1132
rect 1470 1128 1474 1132
rect 46 1118 50 1122
rect 102 1118 106 1122
rect 126 1118 130 1122
rect 206 1118 210 1122
rect 238 1118 242 1122
rect 270 1118 274 1122
rect 326 1118 330 1122
rect 438 1118 442 1122
rect 510 1118 514 1122
rect 534 1118 538 1122
rect 638 1118 642 1122
rect 686 1118 690 1122
rect 734 1118 738 1122
rect 782 1118 786 1122
rect 798 1118 802 1122
rect 830 1118 834 1122
rect 854 1118 858 1122
rect 894 1118 898 1122
rect 1030 1118 1034 1122
rect 1078 1118 1082 1122
rect 1102 1118 1106 1122
rect 1310 1118 1314 1122
rect 1334 1118 1338 1122
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 166 1088 170 1092
rect 366 1088 370 1092
rect 726 1088 730 1092
rect 766 1088 770 1092
rect 974 1088 978 1092
rect 22 1078 26 1082
rect 198 1078 202 1082
rect 246 1078 250 1082
rect 342 1078 346 1082
rect 382 1078 386 1082
rect 390 1078 394 1082
rect 462 1078 466 1082
rect 630 1078 634 1082
rect 750 1078 754 1082
rect 846 1078 850 1082
rect 942 1078 946 1082
rect 974 1078 978 1082
rect 1142 1078 1146 1082
rect 1174 1078 1178 1082
rect 62 1068 66 1072
rect 182 1068 186 1072
rect 334 1068 338 1072
rect 350 1068 354 1072
rect 422 1068 426 1072
rect 486 1068 490 1072
rect 646 1068 650 1072
rect 758 1068 762 1072
rect 790 1068 794 1072
rect 862 1068 866 1072
rect 918 1068 922 1072
rect 934 1068 938 1072
rect 998 1068 1002 1072
rect 1014 1068 1018 1072
rect 1134 1068 1138 1072
rect 1326 1078 1330 1082
rect 1406 1078 1410 1082
rect 1470 1078 1474 1082
rect 1190 1068 1194 1072
rect 1222 1068 1226 1072
rect 1382 1068 1386 1072
rect 1406 1068 1410 1072
rect 1462 1068 1466 1072
rect 70 1059 74 1063
rect 118 1058 122 1062
rect 142 1058 146 1062
rect 198 1058 202 1062
rect 222 1058 226 1062
rect 262 1058 266 1062
rect 294 1058 298 1062
rect 318 1058 322 1062
rect 438 1058 442 1062
rect 502 1058 506 1062
rect 526 1058 530 1062
rect 558 1058 562 1062
rect 590 1058 594 1062
rect 606 1058 610 1062
rect 670 1058 674 1062
rect 694 1058 698 1062
rect 798 1058 802 1062
rect 830 1058 834 1062
rect 902 1058 906 1062
rect 950 1058 954 1062
rect 1038 1058 1042 1062
rect 1070 1058 1074 1062
rect 1094 1058 1098 1062
rect 1118 1058 1122 1062
rect 134 1048 138 1052
rect 166 1048 170 1052
rect 182 1048 186 1052
rect 254 1048 258 1052
rect 286 1048 290 1052
rect 422 1048 426 1052
rect 470 1048 474 1052
rect 534 1048 538 1052
rect 566 1048 570 1052
rect 598 1048 602 1052
rect 662 1048 666 1052
rect 806 1048 810 1052
rect 838 1048 842 1052
rect 846 1048 850 1052
rect 878 1048 882 1052
rect 910 1048 914 1052
rect 1022 1048 1026 1052
rect 1070 1048 1074 1052
rect 1086 1048 1090 1052
rect 1150 1048 1154 1052
rect 110 1038 114 1042
rect 150 1038 154 1042
rect 270 1038 274 1042
rect 294 1038 298 1042
rect 302 1038 306 1042
rect 438 1038 442 1042
rect 518 1038 522 1042
rect 550 1038 554 1042
rect 614 1038 618 1042
rect 678 1038 682 1042
rect 790 1038 794 1042
rect 822 1038 826 1042
rect 870 1038 874 1042
rect 894 1038 898 1042
rect 1030 1038 1034 1042
rect 1078 1038 1082 1042
rect 1102 1038 1106 1042
rect 1238 1038 1242 1042
rect 1278 1058 1282 1062
rect 1286 1058 1290 1062
rect 1310 1058 1314 1062
rect 1342 1058 1346 1062
rect 1366 1058 1370 1062
rect 1430 1058 1434 1062
rect 1446 1058 1450 1062
rect 1254 1048 1258 1052
rect 1318 1048 1322 1052
rect 1374 1048 1378 1052
rect 1414 1048 1418 1052
rect 1270 1038 1274 1042
rect 1302 1038 1306 1042
rect 1350 1038 1354 1042
rect 1358 1038 1362 1042
rect 1430 1038 1434 1042
rect 262 1028 266 1032
rect 118 1018 122 1022
rect 142 1018 146 1022
rect 446 1018 450 1022
rect 526 1018 530 1022
rect 558 1018 562 1022
rect 574 1018 578 1022
rect 622 1018 626 1022
rect 638 1018 642 1022
rect 654 1018 658 1022
rect 670 1018 674 1022
rect 710 1018 714 1022
rect 766 1018 770 1022
rect 830 1018 834 1022
rect 886 1018 890 1022
rect 1046 1018 1050 1022
rect 1054 1018 1058 1022
rect 1094 1018 1098 1022
rect 1214 1018 1218 1022
rect 1246 1018 1250 1022
rect 1294 1018 1298 1022
rect 1326 1018 1330 1022
rect 1422 1018 1426 1022
rect 474 1003 478 1007
rect 481 1003 485 1007
rect 150 988 154 992
rect 278 988 282 992
rect 406 988 410 992
rect 438 988 442 992
rect 518 988 522 992
rect 966 988 970 992
rect 1198 988 1202 992
rect 1254 988 1258 992
rect 1454 988 1458 992
rect 342 978 346 982
rect 630 978 634 982
rect 214 968 218 972
rect 246 968 250 972
rect 254 968 258 972
rect 286 968 290 972
rect 318 968 322 972
rect 350 968 354 972
rect 414 968 418 972
rect 446 968 450 972
rect 526 968 530 972
rect 606 968 610 972
rect 662 968 666 972
rect 710 968 714 972
rect 774 978 778 982
rect 854 978 858 982
rect 782 968 786 972
rect 886 968 890 972
rect 910 968 914 972
rect 1046 968 1050 972
rect 1190 968 1194 972
rect 1358 968 1362 972
rect 1438 968 1442 972
rect 166 958 170 962
rect 230 958 234 962
rect 270 958 274 962
rect 302 958 306 962
rect 334 958 338 962
rect 398 958 402 962
rect 430 958 434 962
rect 510 958 514 962
rect 590 958 594 962
rect 622 958 626 962
rect 646 958 650 962
rect 718 958 722 962
rect 734 958 738 962
rect 766 958 770 962
rect 838 958 842 962
rect 862 958 866 962
rect 870 958 874 962
rect 926 958 930 962
rect 1030 958 1034 962
rect 1174 958 1178 962
rect 1206 958 1210 962
rect 1334 958 1338 962
rect 1342 958 1346 962
rect 1446 958 1450 962
rect 62 948 66 952
rect 94 947 98 951
rect 126 948 130 952
rect 198 948 202 952
rect 222 948 226 952
rect 246 948 250 952
rect 286 948 290 952
rect 310 948 314 952
rect 342 948 346 952
rect 366 948 370 952
rect 406 948 410 952
rect 438 948 442 952
rect 470 948 474 952
rect 518 948 522 952
rect 542 948 546 952
rect 614 948 618 952
rect 694 948 698 952
rect 710 948 714 952
rect 742 948 746 952
rect 774 948 778 952
rect 798 948 802 952
rect 878 948 882 952
rect 902 948 906 952
rect 918 948 922 952
rect 934 948 938 952
rect 982 948 986 952
rect 1038 948 1042 952
rect 1198 948 1202 952
rect 1246 948 1250 952
rect 1326 948 1330 952
rect 1350 948 1354 952
rect 1374 948 1378 952
rect 6 938 10 942
rect 134 938 138 942
rect 158 938 162 942
rect 174 938 178 942
rect 198 938 202 942
rect 318 938 322 942
rect 382 938 386 942
rect 494 938 498 942
rect 558 938 562 942
rect 574 938 578 942
rect 662 938 666 942
rect 678 938 682 942
rect 814 938 818 942
rect 846 938 850 942
rect 950 938 954 942
rect 1022 938 1026 942
rect 1062 938 1066 942
rect 1134 938 1138 942
rect 1174 938 1178 942
rect 1214 938 1218 942
rect 1262 938 1266 942
rect 1302 938 1306 942
rect 1390 938 1394 942
rect 1446 938 1450 942
rect 1462 938 1466 942
rect 150 928 154 932
rect 174 928 178 932
rect 390 928 394 932
rect 502 928 506 932
rect 582 928 586 932
rect 638 928 642 932
rect 822 928 826 932
rect 830 928 834 932
rect 1094 928 1098 932
rect 1102 928 1106 932
rect 1150 928 1154 932
rect 1214 928 1218 932
rect 1270 928 1274 932
rect 1398 928 1402 932
rect 1406 928 1410 932
rect 222 918 226 922
rect 614 918 618 922
rect 742 918 746 922
rect 878 918 882 922
rect 1038 918 1042 922
rect 1078 918 1082 922
rect 1118 918 1122 922
rect 1294 918 1298 922
rect 1318 918 1322 922
rect 986 903 990 907
rect 993 903 997 907
rect 158 888 162 892
rect 286 888 290 892
rect 390 888 394 892
rect 414 888 418 892
rect 446 888 450 892
rect 510 888 514 892
rect 822 888 826 892
rect 1022 888 1026 892
rect 150 878 154 882
rect 334 878 338 882
rect 374 878 378 882
rect 438 878 442 882
rect 6 868 10 872
rect 134 868 138 872
rect 262 868 266 872
rect 326 868 330 872
rect 358 868 362 872
rect 382 868 386 872
rect 406 868 410 872
rect 462 868 466 872
rect 534 878 538 882
rect 630 878 634 882
rect 686 878 690 882
rect 702 878 706 882
rect 798 878 802 882
rect 806 878 810 882
rect 934 878 938 882
rect 974 878 978 882
rect 1006 878 1010 882
rect 1142 878 1146 882
rect 1206 878 1210 882
rect 1238 878 1242 882
rect 1254 878 1258 882
rect 1446 878 1450 882
rect 494 868 498 872
rect 526 868 530 872
rect 542 868 546 872
rect 598 868 602 872
rect 734 868 738 872
rect 790 868 794 872
rect 838 868 842 872
rect 926 868 930 872
rect 1014 868 1018 872
rect 1094 868 1098 872
rect 1134 868 1138 872
rect 1198 868 1202 872
rect 1286 868 1290 872
rect 1422 868 1426 872
rect 1478 868 1482 872
rect 70 858 74 862
rect 94 859 98 863
rect 126 858 130 862
rect 142 858 146 862
rect 246 859 250 863
rect 286 858 290 862
rect 310 858 314 862
rect 358 858 362 862
rect 558 858 562 862
rect 574 858 578 862
rect 654 858 658 862
rect 686 858 690 862
rect 758 858 762 862
rect 774 858 778 862
rect 862 858 866 862
rect 894 858 898 862
rect 910 858 914 862
rect 942 858 946 862
rect 1038 858 1042 862
rect 1070 858 1074 862
rect 1110 858 1114 862
rect 1158 858 1162 862
rect 1182 858 1186 862
rect 1310 858 1314 862
rect 1342 858 1346 862
rect 1366 858 1370 862
rect 1406 858 1410 862
rect 278 848 282 852
rect 342 848 346 852
rect 398 848 402 852
rect 422 848 426 852
rect 430 848 434 852
rect 566 848 570 852
rect 598 848 602 852
rect 662 848 666 852
rect 686 848 690 852
rect 766 848 770 852
rect 838 848 842 852
rect 870 848 874 852
rect 878 848 882 852
rect 1030 848 1034 852
rect 1062 848 1066 852
rect 1102 848 1106 852
rect 1150 848 1154 852
rect 1214 848 1218 852
rect 1286 848 1290 852
rect 1318 848 1322 852
rect 1350 848 1354 852
rect 1358 848 1362 852
rect 1414 848 1418 852
rect 294 838 298 842
rect 358 838 362 842
rect 582 838 586 842
rect 646 838 650 842
rect 678 838 682 842
rect 734 838 738 842
rect 750 838 754 842
rect 854 838 858 842
rect 894 838 898 842
rect 1046 838 1050 842
rect 1078 838 1082 842
rect 1166 838 1170 842
rect 1302 838 1306 842
rect 1334 838 1338 842
rect 1374 838 1378 842
rect 1390 838 1394 842
rect 1398 838 1402 842
rect 990 828 994 832
rect 1070 828 1074 832
rect 1310 828 1314 832
rect 590 818 594 822
rect 638 818 642 822
rect 742 818 746 822
rect 886 818 890 822
rect 1022 818 1026 822
rect 1038 818 1042 822
rect 1158 818 1162 822
rect 1326 818 1330 822
rect 1366 818 1370 822
rect 474 803 478 807
rect 481 803 485 807
rect 6 788 10 792
rect 30 788 34 792
rect 278 788 282 792
rect 430 788 434 792
rect 694 788 698 792
rect 790 788 794 792
rect 1270 788 1274 792
rect 1286 788 1290 792
rect 1446 788 1450 792
rect 182 778 186 782
rect 894 778 898 782
rect 70 768 74 772
rect 582 768 586 772
rect 590 768 594 772
rect 606 768 610 772
rect 638 768 642 772
rect 670 768 674 772
rect 726 768 730 772
rect 782 768 786 772
rect 798 768 802 772
rect 830 768 834 772
rect 870 768 874 772
rect 894 768 898 772
rect 966 768 970 772
rect 982 768 986 772
rect 1438 778 1442 782
rect 1014 768 1018 772
rect 1150 768 1154 772
rect 1302 768 1306 772
rect 566 758 570 762
rect 622 758 626 762
rect 654 758 658 762
rect 686 758 690 762
rect 710 758 714 762
rect 814 758 818 762
rect 846 758 850 762
rect 854 758 858 762
rect 886 758 890 762
rect 950 758 954 762
rect 998 758 1002 762
rect 1318 758 1322 762
rect 22 748 26 752
rect 46 748 50 752
rect 54 748 58 752
rect 118 747 122 751
rect 174 748 178 752
rect 246 747 250 751
rect 366 747 370 751
rect 398 748 402 752
rect 414 748 418 752
rect 454 748 458 752
rect 558 748 562 752
rect 574 748 578 752
rect 614 748 618 752
rect 646 748 650 752
rect 678 748 682 752
rect 718 748 722 752
rect 758 748 762 752
rect 806 748 810 752
rect 838 748 842 752
rect 862 748 866 752
rect 902 748 906 752
rect 918 748 922 752
rect 958 748 962 752
rect 1006 748 1010 752
rect 1030 748 1034 752
rect 1086 747 1090 751
rect 1118 748 1122 752
rect 1182 747 1186 751
rect 1214 748 1218 752
rect 1254 748 1258 752
rect 1310 748 1314 752
rect 1358 748 1362 752
rect 1382 748 1386 752
rect 1462 748 1466 752
rect 134 738 138 742
rect 158 738 162 742
rect 166 738 170 742
rect 262 738 266 742
rect 382 738 386 742
rect 406 738 410 742
rect 446 738 450 742
rect 510 738 514 742
rect 526 738 530 742
rect 542 738 546 742
rect 558 738 562 742
rect 614 738 618 742
rect 638 738 642 742
rect 702 738 706 742
rect 718 738 722 742
rect 750 738 754 742
rect 766 738 770 742
rect 822 738 826 742
rect 934 738 938 742
rect 1046 738 1050 742
rect 1278 738 1282 742
rect 1334 738 1338 742
rect 1446 738 1450 742
rect 150 728 154 732
rect 430 728 434 732
rect 462 728 466 732
rect 518 728 522 732
rect 782 728 786 732
rect 942 728 946 732
rect 958 728 962 732
rect 1054 728 1058 732
rect 502 718 506 722
rect 678 718 682 722
rect 742 718 746 722
rect 862 718 866 722
rect 1246 718 1250 722
rect 1302 718 1306 722
rect 986 703 990 707
rect 993 703 997 707
rect 150 688 154 692
rect 318 688 322 692
rect 438 688 442 692
rect 614 688 618 692
rect 750 688 754 692
rect 806 688 810 692
rect 950 688 954 692
rect 1206 688 1210 692
rect 1230 688 1234 692
rect 1310 688 1314 692
rect 1446 688 1450 692
rect 14 678 18 682
rect 46 678 50 682
rect 110 678 114 682
rect 222 678 226 682
rect 462 678 466 682
rect 558 678 562 682
rect 726 678 730 682
rect 758 678 762 682
rect 790 678 794 682
rect 870 678 874 682
rect 910 678 914 682
rect 46 668 50 672
rect 54 668 58 672
rect 70 668 74 672
rect 118 668 122 672
rect 134 668 138 672
rect 142 668 146 672
rect 190 668 194 672
rect 222 668 226 672
rect 254 668 258 672
rect 374 668 378 672
rect 966 678 970 682
rect 1118 678 1122 682
rect 1286 678 1290 682
rect 1318 678 1322 682
rect 534 668 538 672
rect 550 668 554 672
rect 694 668 698 672
rect 702 668 706 672
rect 742 668 746 672
rect 774 668 778 672
rect 814 668 818 672
rect 830 668 834 672
rect 854 668 858 672
rect 870 668 874 672
rect 878 668 882 672
rect 894 668 898 672
rect 926 668 930 672
rect 942 668 946 672
rect 990 668 994 672
rect 1262 668 1266 672
rect 1270 668 1274 672
rect 1286 668 1290 672
rect 1302 668 1306 672
rect 38 658 42 662
rect 94 658 98 662
rect 166 658 170 662
rect 294 658 298 662
rect 326 658 330 662
rect 358 658 362 662
rect 398 658 402 662
rect 438 658 442 662
rect 470 658 474 662
rect 518 658 522 662
rect 582 658 586 662
rect 614 658 618 662
rect 638 658 642 662
rect 654 658 658 662
rect 678 658 682 662
rect 734 658 738 662
rect 766 658 770 662
rect 822 658 826 662
rect 846 658 850 662
rect 902 658 906 662
rect 1022 659 1026 663
rect 1054 658 1058 662
rect 1118 659 1122 663
rect 1214 658 1218 662
rect 1238 658 1242 662
rect 1262 658 1266 662
rect 1294 658 1298 662
rect 1350 659 1354 663
rect 1382 658 1386 662
rect 1470 658 1474 662
rect 102 648 106 652
rect 158 648 162 652
rect 254 648 258 652
rect 270 648 274 652
rect 302 648 306 652
rect 334 648 338 652
rect 366 648 370 652
rect 446 648 450 652
rect 454 648 458 652
rect 526 648 530 652
rect 590 648 594 652
rect 622 648 626 652
rect 630 648 634 652
rect 686 648 690 652
rect 86 638 90 642
rect 174 638 178 642
rect 190 638 194 642
rect 286 638 290 642
rect 318 638 322 642
rect 358 638 362 642
rect 398 638 402 642
rect 406 638 410 642
rect 446 638 450 642
rect 454 638 458 642
rect 510 638 514 642
rect 518 638 522 642
rect 574 638 578 642
rect 606 638 610 642
rect 646 638 650 642
rect 670 638 674 642
rect 1086 638 1090 642
rect 1438 638 1442 642
rect 278 628 282 632
rect 342 628 346 632
rect 566 628 570 632
rect 678 628 682 632
rect 94 618 98 622
rect 166 618 170 622
rect 238 618 242 622
rect 398 618 402 622
rect 790 618 794 622
rect 838 618 842 622
rect 918 618 922 622
rect 934 618 938 622
rect 474 603 478 607
rect 481 603 485 607
rect 198 588 202 592
rect 214 588 218 592
rect 294 588 298 592
rect 318 588 322 592
rect 422 588 426 592
rect 446 588 450 592
rect 526 588 530 592
rect 614 588 618 592
rect 630 588 634 592
rect 662 588 666 592
rect 798 588 802 592
rect 1302 588 1306 592
rect 1470 588 1474 592
rect 78 578 82 582
rect 502 578 506 582
rect 1166 578 1170 582
rect 1238 578 1242 582
rect 1270 578 1274 582
rect 86 568 90 572
rect 94 568 98 572
rect 118 568 122 572
rect 126 568 130 572
rect 134 568 138 572
rect 150 568 154 572
rect 166 568 170 572
rect 262 568 266 572
rect 326 568 330 572
rect 430 568 434 572
rect 454 568 458 572
rect 510 568 514 572
rect 534 568 538 572
rect 574 568 578 572
rect 638 568 642 572
rect 670 568 674 572
rect 1118 568 1122 572
rect 1158 568 1162 572
rect 1230 568 1234 572
rect 1262 568 1266 572
rect 1294 568 1298 572
rect 102 558 106 562
rect 110 558 114 562
rect 166 558 170 562
rect 174 558 178 562
rect 310 558 314 562
rect 342 558 346 562
rect 414 558 418 562
rect 462 558 466 562
rect 494 558 498 562
rect 550 558 554 562
rect 590 558 594 562
rect 622 558 626 562
rect 654 558 658 562
rect 718 558 722 562
rect 950 558 954 562
rect 990 558 994 562
rect 1102 558 1106 562
rect 1126 558 1130 562
rect 1174 558 1178 562
rect 1214 558 1218 562
rect 1246 558 1250 562
rect 1278 558 1282 562
rect 1310 558 1314 562
rect 38 548 42 552
rect 70 548 74 552
rect 94 548 98 552
rect 118 548 122 552
rect 158 548 162 552
rect 182 548 186 552
rect 294 548 298 552
rect 334 548 338 552
rect 350 548 354 552
rect 422 548 426 552
rect 462 548 466 552
rect 502 548 506 552
rect 542 548 546 552
rect 566 548 570 552
rect 598 548 602 552
rect 630 548 634 552
rect 670 548 674 552
rect 686 548 690 552
rect 838 547 842 551
rect 870 548 874 552
rect 1062 548 1066 552
rect 1158 548 1162 552
rect 1238 548 1242 552
rect 1262 548 1266 552
rect 1302 548 1306 552
rect 1318 548 1322 552
rect 1374 548 1378 552
rect 1406 547 1410 551
rect 54 538 58 542
rect 222 538 226 542
rect 262 538 266 542
rect 366 538 370 542
rect 406 538 410 542
rect 702 538 706 542
rect 790 538 794 542
rect 806 538 810 542
rect 910 538 914 542
rect 966 538 970 542
rect 974 538 978 542
rect 1014 538 1018 542
rect 1038 538 1042 542
rect 1078 538 1082 542
rect 1118 538 1122 542
rect 1142 538 1146 542
rect 1214 538 1218 542
rect 1326 538 1330 542
rect 1342 538 1346 542
rect 1366 538 1370 542
rect 1390 538 1394 542
rect 6 528 10 532
rect 46 528 50 532
rect 230 528 234 532
rect 270 528 274 532
rect 374 528 378 532
rect 382 528 386 532
rect 710 528 714 532
rect 750 528 754 532
rect 758 528 762 532
rect 942 528 946 532
rect 998 528 1002 532
rect 1038 528 1042 532
rect 1070 528 1074 532
rect 1190 528 1194 532
rect 1350 528 1354 532
rect 1406 528 1410 532
rect 142 518 146 522
rect 214 518 218 522
rect 782 518 786 522
rect 902 518 906 522
rect 918 518 922 522
rect 958 518 962 522
rect 1030 518 1034 522
rect 1094 518 1098 522
rect 1134 518 1138 522
rect 1358 518 1362 522
rect 986 503 990 507
rect 993 503 997 507
rect 86 488 90 492
rect 150 488 154 492
rect 206 488 210 492
rect 318 488 322 492
rect 358 488 362 492
rect 390 488 394 492
rect 430 488 434 492
rect 454 488 458 492
rect 502 488 506 492
rect 526 488 530 492
rect 542 488 546 492
rect 582 488 586 492
rect 630 488 634 492
rect 646 488 650 492
rect 702 488 706 492
rect 806 488 810 492
rect 1302 488 1306 492
rect 6 478 10 482
rect 190 478 194 482
rect 286 478 290 482
rect 366 478 370 482
rect 494 478 498 482
rect 510 478 514 482
rect 566 478 570 482
rect 614 478 618 482
rect 670 478 674 482
rect 678 478 682 482
rect 766 478 770 482
rect 846 478 850 482
rect 950 478 954 482
rect 990 478 994 482
rect 1078 478 1082 482
rect 1110 478 1114 482
rect 1278 478 1282 482
rect 54 468 58 472
rect 94 468 98 472
rect 182 468 186 472
rect 278 468 282 472
rect 334 468 338 472
rect 342 468 346 472
rect 374 468 378 472
rect 398 468 402 472
rect 422 468 426 472
rect 462 468 466 472
rect 478 468 482 472
rect 534 468 538 472
rect 558 468 562 472
rect 590 468 594 472
rect 622 468 626 472
rect 662 468 666 472
rect 694 468 698 472
rect 734 468 738 472
rect 742 468 746 472
rect 758 468 762 472
rect 942 468 946 472
rect 30 458 34 462
rect 46 458 50 462
rect 118 458 122 462
rect 142 458 146 462
rect 166 458 170 462
rect 206 458 210 462
rect 238 458 242 462
rect 262 458 266 462
rect 422 458 426 462
rect 590 458 594 462
rect 790 458 794 462
rect 822 458 826 462
rect 846 458 850 462
rect 878 458 882 462
rect 902 458 906 462
rect 926 458 930 462
rect 974 458 978 462
rect 1022 458 1026 462
rect 1046 468 1050 472
rect 1078 468 1082 472
rect 1086 468 1090 472
rect 1102 468 1106 472
rect 1110 468 1114 472
rect 1190 468 1194 472
rect 1326 468 1330 472
rect 1406 468 1410 472
rect 1046 458 1050 462
rect 1134 458 1138 462
rect 1150 458 1154 462
rect 1174 458 1178 462
rect 1214 458 1218 462
rect 1238 458 1242 462
rect 1278 458 1282 462
rect 1302 458 1306 462
rect 1342 458 1346 462
rect 1374 459 1378 463
rect 70 448 74 452
rect 78 448 82 452
rect 126 448 130 452
rect 134 448 138 452
rect 198 448 202 452
rect 230 448 234 452
rect 294 448 298 452
rect 310 448 314 452
rect 318 448 322 452
rect 358 448 362 452
rect 438 448 442 452
rect 446 448 450 452
rect 518 448 522 452
rect 574 448 578 452
rect 638 448 642 452
rect 710 448 714 452
rect 726 448 730 452
rect 798 448 802 452
rect 830 448 834 452
rect 846 448 850 452
rect 870 448 874 452
rect 974 448 978 452
rect 1006 448 1010 452
rect 1070 448 1074 452
rect 1142 448 1146 452
rect 1174 448 1178 452
rect 1190 448 1194 452
rect 1222 448 1226 452
rect 1230 448 1234 452
rect 1286 448 1290 452
rect 1294 448 1298 452
rect 110 438 114 442
rect 150 438 154 442
rect 214 438 218 442
rect 246 438 250 442
rect 678 438 682 442
rect 782 438 786 442
rect 814 438 818 442
rect 854 438 858 442
rect 886 438 890 442
rect 966 438 970 442
rect 1022 438 1026 442
rect 1038 438 1042 442
rect 1158 438 1162 442
rect 1206 438 1210 442
rect 1246 438 1250 442
rect 1254 438 1258 442
rect 1270 438 1274 442
rect 1310 438 1314 442
rect 118 428 122 432
rect 238 428 242 432
rect 878 428 882 432
rect 958 428 962 432
rect 790 418 794 422
rect 918 418 922 422
rect 1214 418 1218 422
rect 1446 418 1450 422
rect 474 403 478 407
rect 481 403 485 407
rect 46 388 50 392
rect 102 388 106 392
rect 142 388 146 392
rect 174 388 178 392
rect 238 388 242 392
rect 382 388 386 392
rect 454 388 458 392
rect 518 388 522 392
rect 542 388 546 392
rect 550 388 554 392
rect 598 388 602 392
rect 654 388 658 392
rect 718 388 722 392
rect 838 388 842 392
rect 974 388 978 392
rect 1150 388 1154 392
rect 1238 388 1242 392
rect 1262 388 1266 392
rect 1334 388 1338 392
rect 414 378 418 382
rect 94 368 98 372
rect 134 368 138 372
rect 182 368 186 372
rect 214 368 218 372
rect 230 368 234 372
rect 246 368 250 372
rect 350 368 354 372
rect 390 368 394 372
rect 462 368 466 372
rect 510 368 514 372
rect 558 368 562 372
rect 590 368 594 372
rect 790 368 794 372
rect 806 368 810 372
rect 918 368 922 372
rect 1022 378 1026 382
rect 1030 368 1034 372
rect 1230 368 1234 372
rect 1286 368 1290 372
rect 1342 368 1346 372
rect 1366 368 1370 372
rect 1382 368 1386 372
rect 1398 368 1402 372
rect 1406 368 1410 372
rect 1438 368 1442 372
rect 1454 368 1458 372
rect 110 358 114 362
rect 118 358 122 362
rect 150 358 154 362
rect 166 358 170 362
rect 198 358 202 362
rect 238 358 242 362
rect 310 358 314 362
rect 318 358 322 362
rect 374 358 378 362
rect 446 358 450 362
rect 526 358 530 362
rect 574 358 578 362
rect 606 358 610 362
rect 662 358 666 362
rect 710 358 714 362
rect 726 358 730 362
rect 774 358 778 362
rect 822 358 826 362
rect 830 358 834 362
rect 934 358 938 362
rect 942 358 946 362
rect 1006 358 1010 362
rect 1078 358 1082 362
rect 1214 358 1218 362
rect 1246 358 1250 362
rect 1254 358 1258 362
rect 1278 358 1282 362
rect 1326 358 1330 362
rect 1358 358 1362 362
rect 1414 358 1418 362
rect 1422 358 1426 362
rect 6 348 10 352
rect 30 348 34 352
rect 54 348 58 352
rect 126 348 130 352
rect 182 348 186 352
rect 206 348 210 352
rect 230 348 234 352
rect 238 348 242 352
rect 262 348 266 352
rect 382 348 386 352
rect 454 348 458 352
rect 566 348 570 352
rect 598 348 602 352
rect 614 348 618 352
rect 686 348 690 352
rect 702 348 706 352
rect 726 348 730 352
rect 766 348 770 352
rect 814 348 818 352
rect 838 348 842 352
rect 862 348 866 352
rect 902 348 906 352
rect 926 348 930 352
rect 950 348 954 352
rect 990 348 994 352
rect 1022 348 1026 352
rect 1046 348 1050 352
rect 1118 348 1122 352
rect 1134 348 1138 352
rect 1182 348 1186 352
rect 1238 348 1242 352
rect 1318 348 1322 352
rect 1334 348 1338 352
rect 1366 348 1370 352
rect 1406 348 1410 352
rect 1430 348 1434 352
rect 70 338 74 342
rect 94 338 98 342
rect 158 338 162 342
rect 278 338 282 342
rect 294 338 298 342
rect 318 338 322 342
rect 406 338 410 342
rect 510 338 514 342
rect 630 338 634 342
rect 678 338 682 342
rect 742 338 746 342
rect 790 338 794 342
rect 886 338 890 342
rect 1062 338 1066 342
rect 1078 338 1082 342
rect 1158 338 1162 342
rect 1198 338 1202 342
rect 1270 338 1274 342
rect 1294 338 1298 342
rect 1470 338 1474 342
rect 78 328 82 332
rect 286 328 290 332
rect 350 328 354 332
rect 366 328 370 332
rect 438 328 442 332
rect 494 328 498 332
rect 534 328 538 332
rect 638 328 642 332
rect 646 328 650 332
rect 662 328 666 332
rect 710 328 714 332
rect 878 328 882 332
rect 950 328 954 332
rect 1070 328 1074 332
rect 1110 328 1114 332
rect 1118 328 1122 332
rect 1190 328 1194 332
rect 22 318 26 322
rect 302 318 306 322
rect 870 318 874 322
rect 1390 318 1394 322
rect 986 303 990 307
rect 993 303 997 307
rect 126 288 130 292
rect 142 288 146 292
rect 182 288 186 292
rect 246 288 250 292
rect 270 288 274 292
rect 382 288 386 292
rect 398 288 402 292
rect 454 288 458 292
rect 486 288 490 292
rect 534 288 538 292
rect 566 288 570 292
rect 598 288 602 292
rect 806 288 810 292
rect 838 288 842 292
rect 1126 288 1130 292
rect 1350 288 1354 292
rect 1430 288 1434 292
rect 6 278 10 282
rect 46 278 50 282
rect 318 278 322 282
rect 350 278 354 282
rect 358 278 362 282
rect 510 278 514 282
rect 542 278 546 282
rect 574 278 578 282
rect 614 278 618 282
rect 678 278 682 282
rect 718 278 722 282
rect 734 278 738 282
rect 926 278 930 282
rect 1014 278 1018 282
rect 1078 278 1082 282
rect 1086 278 1090 282
rect 1102 278 1106 282
rect 1190 278 1194 282
rect 1254 278 1258 282
rect 1406 278 1410 282
rect 1470 278 1474 282
rect 38 268 42 272
rect 54 268 58 272
rect 238 268 242 272
rect 310 268 314 272
rect 318 268 322 272
rect 358 268 362 272
rect 390 268 394 272
rect 406 268 410 272
rect 462 268 466 272
rect 518 268 522 272
rect 550 268 554 272
rect 614 268 618 272
rect 622 268 626 272
rect 646 268 650 272
rect 742 268 746 272
rect 758 268 762 272
rect 958 268 962 272
rect 1046 268 1050 272
rect 1070 268 1074 272
rect 1134 268 1138 272
rect 1158 268 1162 272
rect 1166 268 1170 272
rect 1198 268 1202 272
rect 1262 268 1266 272
rect 1374 268 1378 272
rect 1414 268 1418 272
rect 70 258 74 262
rect 94 258 98 262
rect 126 258 130 262
rect 158 258 162 262
rect 182 258 186 262
rect 214 258 218 262
rect 270 258 274 262
rect 438 258 442 262
rect 646 258 650 262
rect 702 258 706 262
rect 782 258 786 262
rect 814 258 818 262
rect 838 258 842 262
rect 870 258 874 262
rect 902 258 906 262
rect 942 258 946 262
rect 974 258 978 262
rect 1174 258 1178 262
rect 1214 258 1218 262
rect 1230 258 1234 262
rect 1278 258 1282 262
rect 1294 258 1298 262
rect 1318 258 1322 262
rect 1350 258 1354 262
rect 38 248 42 252
rect 102 248 106 252
rect 134 248 138 252
rect 166 248 170 252
rect 206 248 210 252
rect 254 248 258 252
rect 262 248 266 252
rect 294 248 298 252
rect 406 248 410 252
rect 534 248 538 252
rect 710 248 714 252
rect 726 248 730 252
rect 790 248 794 252
rect 830 248 834 252
rect 862 248 866 252
rect 894 248 898 252
rect 958 248 962 252
rect 1046 248 1050 252
rect 1086 248 1090 252
rect 1118 248 1122 252
rect 1142 248 1146 252
rect 1182 248 1186 252
rect 1222 248 1226 252
rect 1294 248 1298 252
rect 1342 248 1346 252
rect 86 238 90 242
rect 118 238 122 242
rect 150 238 154 242
rect 190 238 194 242
rect 214 238 218 242
rect 238 238 242 242
rect 278 238 282 242
rect 694 238 698 242
rect 702 238 706 242
rect 774 238 778 242
rect 806 238 810 242
rect 846 238 850 242
rect 878 238 882 242
rect 902 238 906 242
rect 910 238 914 242
rect 974 238 978 242
rect 982 238 986 242
rect 1046 238 1050 242
rect 1110 238 1114 242
rect 1222 238 1226 242
rect 1302 238 1306 242
rect 1342 238 1346 242
rect 1358 238 1362 242
rect 94 228 98 232
rect 654 228 658 232
rect 1150 228 1154 232
rect 782 218 786 222
rect 870 218 874 222
rect 1230 218 1234 222
rect 1294 218 1298 222
rect 1382 218 1386 222
rect 474 203 478 207
rect 481 203 485 207
rect 78 188 82 192
rect 134 188 138 192
rect 166 188 170 192
rect 318 188 322 192
rect 334 188 338 192
rect 366 188 370 192
rect 406 188 410 192
rect 454 188 458 192
rect 502 188 506 192
rect 534 188 538 192
rect 566 188 570 192
rect 678 188 682 192
rect 750 188 754 192
rect 854 188 858 192
rect 886 188 890 192
rect 990 188 994 192
rect 1222 188 1226 192
rect 1246 188 1250 192
rect 1294 188 1298 192
rect 1358 188 1362 192
rect 1374 188 1378 192
rect 1382 188 1386 192
rect 1398 188 1402 192
rect 918 178 922 182
rect 1022 178 1026 182
rect 1166 178 1170 182
rect 70 168 74 172
rect 126 168 130 172
rect 158 168 162 172
rect 238 168 242 172
rect 246 168 250 172
rect 702 168 706 172
rect 742 168 746 172
rect 822 168 826 172
rect 862 168 866 172
rect 894 168 898 172
rect 926 168 930 172
rect 1030 168 1034 172
rect 1158 168 1162 172
rect 1222 168 1226 172
rect 1254 168 1258 172
rect 1286 168 1290 172
rect 1350 168 1354 172
rect 1470 168 1474 172
rect 86 158 90 162
rect 142 158 146 162
rect 174 158 178 162
rect 230 158 234 162
rect 262 158 266 162
rect 302 158 306 162
rect 350 158 354 162
rect 518 158 522 162
rect 614 158 618 162
rect 718 158 722 162
rect 726 158 730 162
rect 838 158 842 162
rect 846 158 850 162
rect 878 158 882 162
rect 910 158 914 162
rect 1006 158 1010 162
rect 1110 158 1114 162
rect 1174 158 1178 162
rect 1182 158 1186 162
rect 1198 158 1202 162
rect 1238 158 1242 162
rect 1270 158 1274 162
rect 1334 158 1338 162
rect 6 148 10 152
rect 78 148 82 152
rect 94 148 98 152
rect 134 148 138 152
rect 166 148 170 152
rect 182 148 186 152
rect 254 148 258 152
rect 270 148 274 152
rect 318 148 322 152
rect 374 148 378 152
rect 422 148 426 152
rect 494 148 498 152
rect 598 148 602 152
rect 710 148 714 152
rect 734 148 738 152
rect 774 148 778 152
rect 830 148 834 152
rect 854 148 858 152
rect 886 148 890 152
rect 918 148 922 152
rect 974 148 978 152
rect 1022 148 1026 152
rect 1046 148 1050 152
rect 1142 148 1146 152
rect 1166 148 1170 152
rect 1214 148 1218 152
rect 1246 148 1250 152
rect 1278 148 1282 152
rect 1326 148 1330 152
rect 1342 148 1346 152
rect 1414 148 1418 152
rect 1422 148 1426 152
rect 38 138 42 142
rect 54 138 58 142
rect 198 138 202 142
rect 286 138 290 142
rect 326 138 330 142
rect 438 138 442 142
rect 550 138 554 142
rect 622 138 626 142
rect 630 138 634 142
rect 646 138 650 142
rect 686 138 690 142
rect 790 138 794 142
rect 806 138 810 142
rect 942 138 946 142
rect 958 138 962 142
rect 1062 138 1066 142
rect 1110 138 1114 142
rect 1126 138 1130 142
rect 1198 138 1202 142
rect 1310 138 1314 142
rect 30 128 34 132
rect 206 128 210 132
rect 222 128 226 132
rect 294 128 298 132
rect 342 128 346 132
rect 390 128 394 132
rect 398 128 402 132
rect 422 128 426 132
rect 430 128 434 132
rect 462 128 466 132
rect 526 128 530 132
rect 542 128 546 132
rect 574 128 578 132
rect 622 128 626 132
rect 662 128 666 132
rect 758 128 762 132
rect 782 128 786 132
rect 966 128 970 132
rect 998 128 1002 132
rect 1070 128 1074 132
rect 1078 128 1082 132
rect 1302 128 1306 132
rect 1366 128 1370 132
rect 1390 128 1394 132
rect 110 118 114 122
rect 710 118 714 122
rect 830 118 834 122
rect 986 103 990 107
rect 993 103 997 107
rect 22 88 26 92
rect 62 88 66 92
rect 134 88 138 92
rect 182 88 186 92
rect 214 88 218 92
rect 310 88 314 92
rect 350 88 354 92
rect 406 88 410 92
rect 486 88 490 92
rect 614 88 618 92
rect 742 88 746 92
rect 766 88 770 92
rect 806 88 810 92
rect 846 88 850 92
rect 934 88 938 92
rect 1014 88 1018 92
rect 1038 88 1042 92
rect 1134 88 1138 92
rect 1214 88 1218 92
rect 1246 88 1250 92
rect 1294 88 1298 92
rect 1318 88 1322 92
rect 1342 88 1346 92
rect 1390 88 1394 92
rect 1398 88 1402 92
rect 1430 88 1434 92
rect 6 78 10 82
rect 150 78 154 82
rect 158 78 162 82
rect 198 78 202 82
rect 238 78 242 82
rect 334 78 338 82
rect 366 78 370 82
rect 566 78 570 82
rect 670 78 674 82
rect 798 78 802 82
rect 894 78 898 82
rect 958 78 962 82
rect 966 78 970 82
rect 1054 78 1058 82
rect 1062 78 1066 82
rect 1182 78 1186 82
rect 1286 78 1290 82
rect 1326 78 1330 82
rect 1366 78 1370 82
rect 1422 78 1426 82
rect 1454 78 1458 82
rect 1478 78 1482 82
rect 38 68 42 72
rect 46 68 50 72
rect 94 68 98 72
rect 86 58 90 62
rect 118 68 122 72
rect 166 68 170 72
rect 206 68 210 72
rect 270 68 274 72
rect 238 58 242 62
rect 262 58 266 62
rect 294 68 298 72
rect 366 68 370 72
rect 430 68 434 72
rect 454 68 458 72
rect 518 68 522 72
rect 598 68 602 72
rect 622 68 626 72
rect 662 68 666 72
rect 710 68 714 72
rect 742 68 746 72
rect 766 68 770 72
rect 782 68 786 72
rect 822 68 826 72
rect 830 68 834 72
rect 902 68 906 72
rect 926 68 930 72
rect 1094 68 1098 72
rect 1102 68 1106 72
rect 1126 68 1130 72
rect 1158 68 1162 72
rect 1222 68 1226 72
rect 1278 68 1282 72
rect 1310 68 1314 72
rect 1374 68 1378 72
rect 1414 68 1418 72
rect 1446 68 1450 72
rect 318 58 322 62
rect 390 58 394 62
rect 438 58 442 62
rect 550 58 554 62
rect 646 58 650 62
rect 662 58 666 62
rect 694 58 698 62
rect 870 58 874 62
rect 902 58 906 62
rect 982 58 986 62
rect 1078 58 1082 62
rect 1094 58 1098 62
rect 1110 58 1114 62
rect 1150 58 1154 62
rect 1198 58 1202 62
rect 1246 58 1250 62
rect 1262 58 1266 62
rect 1350 58 1354 62
rect 70 48 74 52
rect 118 48 122 52
rect 142 48 146 52
rect 246 48 250 52
rect 294 48 298 52
rect 318 48 322 52
rect 342 48 346 52
rect 414 48 418 52
rect 502 48 506 52
rect 590 48 594 52
rect 622 48 626 52
rect 718 48 722 52
rect 742 48 746 52
rect 766 48 770 52
rect 854 48 858 52
rect 918 48 922 52
rect 982 48 986 52
rect 1126 48 1130 52
rect 1174 48 1178 52
rect 1206 48 1210 52
rect 1246 48 1250 52
rect 1294 48 1298 52
rect 1350 48 1354 52
rect 102 38 106 42
rect 278 38 282 42
rect 494 38 498 42
rect 566 38 570 42
rect 1078 38 1082 42
rect 1238 38 1242 42
rect 1342 38 1346 42
rect 542 28 546 32
rect 1166 28 1170 32
rect 474 3 478 7
rect 481 3 485 7
<< metal2 >>
rect 86 1438 90 1442
rect 166 1441 170 1442
rect 166 1438 177 1441
rect 50 1358 54 1361
rect 30 1342 33 1348
rect 58 1338 62 1341
rect 6 1322 9 1328
rect 6 1272 9 1308
rect 30 1282 33 1338
rect 86 1332 89 1438
rect 114 1358 118 1361
rect 138 1358 142 1361
rect 94 1352 97 1358
rect 98 1338 102 1341
rect 146 1338 150 1341
rect 82 1328 86 1331
rect 26 1248 30 1251
rect 14 1182 17 1218
rect 38 1192 41 1268
rect 46 1252 49 1318
rect 54 1252 57 1258
rect 38 1172 41 1178
rect 50 1158 54 1161
rect 62 1152 65 1308
rect 70 1242 73 1318
rect 94 1282 97 1338
rect 118 1312 121 1338
rect 174 1332 177 1438
rect 238 1438 242 1442
rect 342 1438 346 1442
rect 422 1438 426 1442
rect 542 1438 546 1442
rect 590 1438 594 1442
rect 630 1438 634 1442
rect 654 1438 658 1442
rect 670 1438 674 1442
rect 694 1438 698 1442
rect 718 1438 722 1442
rect 742 1438 746 1442
rect 758 1438 762 1442
rect 854 1438 858 1442
rect 878 1438 882 1442
rect 894 1438 898 1442
rect 918 1441 922 1442
rect 918 1438 929 1441
rect 210 1358 214 1361
rect 238 1352 241 1438
rect 342 1412 345 1438
rect 422 1392 425 1438
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 485 1403 488 1407
rect 270 1362 273 1368
rect 342 1362 345 1378
rect 362 1368 366 1371
rect 422 1362 425 1388
rect 510 1362 513 1378
rect 378 1358 390 1361
rect 450 1358 454 1361
rect 482 1358 486 1361
rect 226 1348 230 1351
rect 262 1351 265 1358
rect 262 1348 270 1351
rect 182 1332 185 1338
rect 126 1282 129 1318
rect 106 1268 110 1271
rect 118 1262 121 1268
rect 130 1258 134 1261
rect 78 1252 81 1258
rect 122 1248 126 1251
rect 70 1192 73 1198
rect 78 1152 81 1218
rect 86 1202 89 1248
rect 142 1242 145 1298
rect 158 1241 161 1318
rect 174 1292 177 1328
rect 190 1262 193 1268
rect 178 1258 182 1261
rect 178 1248 182 1251
rect 198 1242 201 1348
rect 246 1342 249 1348
rect 278 1342 281 1358
rect 438 1352 441 1358
rect 290 1348 294 1351
rect 354 1348 358 1351
rect 458 1348 462 1351
rect 326 1342 329 1348
rect 398 1342 401 1348
rect 510 1342 513 1348
rect 338 1338 342 1341
rect 354 1338 358 1341
rect 386 1338 390 1341
rect 474 1338 478 1341
rect 158 1238 166 1241
rect 94 1172 97 1198
rect 134 1181 137 1218
rect 158 1192 161 1198
rect 134 1178 142 1181
rect 126 1172 129 1178
rect 138 1158 142 1161
rect 50 1148 54 1151
rect 98 1148 102 1151
rect 6 1142 9 1148
rect 22 1082 25 1148
rect 62 1142 65 1148
rect 110 1122 113 1158
rect 138 1148 142 1151
rect 150 1142 153 1158
rect 158 1142 161 1148
rect 46 1042 49 1118
rect 62 1052 65 1068
rect 102 1062 105 1118
rect 62 952 65 1048
rect 70 1022 73 1059
rect 114 1058 118 1061
rect 106 1038 110 1041
rect 118 972 121 1018
rect 126 972 129 1118
rect 150 1102 153 1138
rect 166 1092 169 1168
rect 174 1151 177 1218
rect 206 1171 209 1318
rect 222 1312 225 1338
rect 254 1332 257 1338
rect 394 1328 398 1331
rect 310 1322 313 1328
rect 266 1318 270 1321
rect 222 1292 225 1298
rect 254 1282 257 1308
rect 350 1282 353 1308
rect 390 1282 393 1328
rect 218 1278 222 1281
rect 338 1278 342 1281
rect 218 1268 222 1271
rect 230 1271 233 1278
rect 310 1272 313 1278
rect 382 1272 385 1278
rect 230 1268 238 1271
rect 222 1252 225 1258
rect 202 1168 209 1171
rect 194 1158 198 1161
rect 214 1152 217 1238
rect 230 1192 233 1268
rect 350 1262 353 1268
rect 414 1262 417 1278
rect 274 1258 278 1261
rect 314 1258 318 1261
rect 238 1252 241 1258
rect 430 1252 433 1318
rect 438 1282 441 1338
rect 526 1332 529 1398
rect 542 1361 545 1438
rect 542 1358 550 1361
rect 550 1352 553 1358
rect 534 1282 537 1318
rect 558 1302 561 1328
rect 582 1282 585 1348
rect 442 1278 446 1281
rect 522 1278 526 1281
rect 578 1278 582 1281
rect 590 1272 593 1438
rect 598 1352 601 1358
rect 614 1342 617 1408
rect 630 1362 633 1438
rect 654 1412 657 1438
rect 622 1352 625 1358
rect 630 1352 633 1358
rect 654 1352 657 1358
rect 646 1342 649 1348
rect 618 1338 622 1341
rect 614 1282 617 1318
rect 646 1272 649 1338
rect 610 1268 614 1271
rect 258 1248 262 1251
rect 306 1248 310 1251
rect 386 1248 390 1251
rect 262 1202 265 1248
rect 278 1242 281 1248
rect 294 1232 297 1248
rect 446 1242 449 1268
rect 526 1262 529 1268
rect 546 1258 558 1261
rect 502 1252 505 1258
rect 474 1248 478 1251
rect 514 1248 518 1251
rect 578 1248 582 1251
rect 462 1241 465 1248
rect 462 1238 494 1241
rect 270 1181 273 1218
rect 262 1178 273 1181
rect 250 1158 254 1161
rect 174 1148 190 1151
rect 190 1072 193 1128
rect 198 1082 201 1088
rect 186 1068 190 1071
rect 198 1062 201 1068
rect 134 1032 137 1048
rect 142 1042 145 1058
rect 166 1052 169 1058
rect 182 1052 185 1058
rect 206 1052 209 1118
rect 214 1061 217 1148
rect 246 1142 249 1158
rect 262 1152 265 1178
rect 270 1162 273 1168
rect 350 1162 353 1168
rect 286 1152 289 1158
rect 302 1142 305 1148
rect 234 1138 238 1141
rect 322 1138 326 1141
rect 306 1128 310 1131
rect 214 1058 222 1061
rect 238 1052 241 1118
rect 246 1072 249 1078
rect 270 1062 273 1118
rect 262 1052 265 1058
rect 286 1052 289 1098
rect 318 1062 321 1068
rect 298 1058 302 1061
rect 326 1052 329 1118
rect 350 1112 353 1128
rect 338 1078 342 1081
rect 250 1048 254 1051
rect 150 1042 153 1048
rect 94 951 97 958
rect 126 952 129 958
rect 66 948 73 951
rect 6 942 9 948
rect 6 872 9 878
rect 70 862 73 948
rect 134 932 137 938
rect 142 912 145 1018
rect 150 992 153 1018
rect 166 962 169 1028
rect 170 958 174 961
rect 198 952 201 978
rect 210 968 214 971
rect 222 952 225 988
rect 254 982 257 1048
rect 262 1032 265 1038
rect 270 1032 273 1038
rect 286 1012 289 1048
rect 302 1042 305 1048
rect 294 1032 297 1038
rect 334 1022 337 1068
rect 274 988 278 991
rect 246 972 249 978
rect 258 968 262 971
rect 270 962 273 978
rect 286 972 289 998
rect 302 962 305 978
rect 234 958 238 961
rect 310 952 313 988
rect 322 968 326 971
rect 334 962 337 1008
rect 350 982 353 1068
rect 342 972 345 978
rect 250 948 254 951
rect 174 942 177 948
rect 126 862 129 908
rect 150 882 153 928
rect 158 912 161 938
rect 170 928 174 931
rect 162 888 166 891
rect 138 868 142 871
rect 6 792 9 828
rect 30 792 33 808
rect 46 752 49 778
rect 70 772 73 858
rect 94 852 97 859
rect 142 852 145 858
rect 54 752 57 758
rect 62 752 65 768
rect 26 748 30 751
rect 14 682 17 748
rect 118 742 121 747
rect 134 742 137 758
rect 150 732 153 878
rect 178 778 182 781
rect 174 752 177 768
rect 158 732 161 738
rect 166 732 169 738
rect 106 678 110 681
rect 14 632 17 678
rect 46 672 49 678
rect 142 672 145 708
rect 150 692 153 728
rect 190 672 193 678
rect 130 668 134 671
rect 38 652 41 658
rect 34 548 38 551
rect 6 532 9 538
rect 46 532 49 668
rect 54 612 57 668
rect 70 662 73 668
rect 94 662 97 668
rect 118 662 121 668
rect 166 662 169 668
rect 106 648 110 651
rect 162 648 166 651
rect 86 642 89 648
rect 178 638 190 641
rect 78 582 81 588
rect 94 572 97 618
rect 166 582 169 618
rect 198 592 201 938
rect 222 772 225 918
rect 286 892 289 948
rect 318 942 321 948
rect 342 942 345 948
rect 350 912 353 968
rect 358 922 361 1128
rect 366 1092 369 1168
rect 374 1152 377 1168
rect 382 1162 385 1198
rect 382 1102 385 1158
rect 406 1142 409 1178
rect 414 1162 417 1218
rect 422 1192 425 1228
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 485 1203 488 1207
rect 458 1138 462 1141
rect 414 1132 417 1138
rect 430 1132 433 1138
rect 462 1122 465 1128
rect 394 1078 398 1081
rect 382 1072 385 1078
rect 422 1072 425 1118
rect 422 1042 425 1048
rect 406 992 409 998
rect 394 958 398 961
rect 366 942 369 948
rect 406 942 409 948
rect 246 832 249 859
rect 262 762 265 868
rect 278 852 281 878
rect 334 872 337 878
rect 358 872 361 918
rect 374 882 377 888
rect 382 881 385 938
rect 390 922 393 928
rect 390 892 393 908
rect 414 892 417 968
rect 430 962 433 1098
rect 438 1062 441 1118
rect 462 1082 465 1118
rect 470 1052 473 1138
rect 490 1128 494 1131
rect 502 1082 505 1218
rect 558 1192 561 1238
rect 590 1222 593 1268
rect 622 1262 625 1268
rect 618 1248 622 1251
rect 634 1238 646 1241
rect 654 1232 657 1348
rect 514 1158 518 1161
rect 538 1138 542 1141
rect 518 1132 521 1138
rect 550 1132 553 1138
rect 490 1068 494 1071
rect 502 1062 505 1068
rect 438 1042 441 1048
rect 510 1041 513 1118
rect 534 1062 537 1118
rect 558 1062 561 1078
rect 566 1062 569 1218
rect 606 1152 609 1228
rect 630 1172 633 1188
rect 582 1122 585 1128
rect 590 1122 593 1128
rect 606 1092 609 1148
rect 614 1102 617 1158
rect 622 1152 625 1168
rect 638 1152 641 1218
rect 654 1142 657 1178
rect 642 1128 646 1131
rect 630 1092 633 1108
rect 590 1062 593 1088
rect 606 1072 609 1088
rect 630 1082 633 1088
rect 522 1058 526 1061
rect 602 1058 606 1061
rect 538 1048 542 1051
rect 550 1042 553 1058
rect 570 1048 574 1051
rect 602 1048 606 1051
rect 510 1038 518 1041
rect 618 1038 622 1041
rect 638 1032 641 1118
rect 646 1072 649 1098
rect 646 1052 649 1068
rect 662 1061 665 1148
rect 670 1102 673 1438
rect 694 1372 697 1438
rect 718 1412 721 1438
rect 694 1362 697 1368
rect 718 1362 721 1378
rect 678 1342 681 1348
rect 698 1338 702 1341
rect 678 1282 681 1288
rect 686 1252 689 1318
rect 702 1262 705 1338
rect 726 1332 729 1398
rect 742 1382 745 1438
rect 758 1402 761 1438
rect 774 1362 777 1378
rect 798 1362 801 1368
rect 818 1358 822 1361
rect 754 1348 758 1351
rect 766 1342 769 1358
rect 790 1342 793 1348
rect 814 1342 817 1348
rect 694 1162 697 1258
rect 718 1251 721 1318
rect 726 1282 729 1318
rect 746 1258 750 1261
rect 718 1248 726 1251
rect 702 1162 705 1248
rect 710 1172 713 1178
rect 722 1168 729 1171
rect 678 1152 681 1158
rect 682 1138 686 1141
rect 702 1122 705 1158
rect 710 1152 713 1158
rect 662 1058 670 1061
rect 658 1048 662 1051
rect 686 1041 689 1118
rect 694 1062 697 1068
rect 682 1038 689 1041
rect 446 1002 449 1018
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 485 1003 488 1007
rect 518 992 521 1028
rect 526 1012 529 1018
rect 558 1002 561 1018
rect 574 992 577 1018
rect 442 988 446 991
rect 450 968 457 971
rect 430 882 433 958
rect 442 948 446 951
rect 454 942 457 968
rect 466 948 470 951
rect 494 942 497 978
rect 530 968 537 971
rect 506 958 510 961
rect 522 948 526 951
rect 446 892 449 938
rect 382 878 393 881
rect 322 868 326 871
rect 378 868 382 871
rect 310 862 313 868
rect 290 858 294 861
rect 358 852 361 858
rect 346 848 350 851
rect 390 842 393 878
rect 402 868 406 871
rect 422 852 425 868
rect 430 852 433 858
rect 402 848 406 851
rect 298 838 302 841
rect 354 838 358 841
rect 278 792 281 838
rect 430 792 433 828
rect 438 782 441 878
rect 494 872 497 938
rect 502 902 505 928
rect 510 892 513 938
rect 534 932 537 968
rect 542 952 545 958
rect 574 942 577 978
rect 590 962 593 978
rect 598 942 601 988
rect 622 972 625 1018
rect 630 982 633 988
rect 638 981 641 1018
rect 638 978 649 981
rect 610 968 614 971
rect 626 958 630 961
rect 610 948 614 951
rect 562 938 566 941
rect 586 928 590 931
rect 534 902 537 918
rect 534 882 537 898
rect 526 872 529 878
rect 546 868 550 871
rect 462 822 465 868
rect 472 803 474 807
rect 478 803 481 807
rect 485 803 488 807
rect 222 682 225 718
rect 230 672 233 748
rect 246 742 249 747
rect 262 742 265 758
rect 366 742 369 747
rect 382 742 385 758
rect 398 752 401 768
rect 454 752 457 788
rect 418 748 422 751
rect 406 732 409 738
rect 430 732 433 748
rect 438 738 446 741
rect 318 692 321 728
rect 334 692 337 698
rect 438 692 441 738
rect 510 732 513 738
rect 518 732 521 868
rect 558 852 561 858
rect 566 852 569 908
rect 598 872 601 938
rect 638 932 641 968
rect 646 962 649 978
rect 654 962 657 1018
rect 662 962 665 968
rect 658 938 662 941
rect 614 862 617 918
rect 630 882 633 908
rect 626 878 630 881
rect 670 871 673 1018
rect 678 942 681 1008
rect 710 982 713 1018
rect 710 962 713 968
rect 718 962 721 1138
rect 726 1092 729 1168
rect 750 1162 753 1218
rect 738 1158 742 1161
rect 754 1138 761 1141
rect 734 1042 737 1118
rect 746 1078 750 1081
rect 758 1072 761 1138
rect 766 1132 769 1288
rect 774 1282 777 1328
rect 782 1282 785 1318
rect 806 1302 809 1318
rect 830 1302 833 1318
rect 838 1301 841 1338
rect 846 1312 849 1328
rect 854 1312 857 1438
rect 878 1412 881 1438
rect 878 1342 881 1348
rect 894 1341 897 1438
rect 906 1358 913 1361
rect 890 1338 897 1341
rect 902 1342 905 1348
rect 910 1342 913 1358
rect 926 1352 929 1438
rect 942 1438 946 1442
rect 1350 1438 1354 1442
rect 1366 1438 1370 1442
rect 886 1332 889 1338
rect 838 1298 849 1301
rect 806 1252 809 1258
rect 814 1222 817 1268
rect 822 1252 825 1298
rect 830 1262 833 1278
rect 838 1262 841 1268
rect 830 1222 833 1258
rect 838 1242 841 1258
rect 822 1218 830 1221
rect 806 1162 809 1218
rect 814 1142 817 1218
rect 822 1142 825 1218
rect 830 1162 833 1168
rect 846 1142 849 1298
rect 854 1242 857 1248
rect 862 1172 865 1298
rect 870 1242 873 1318
rect 894 1282 897 1308
rect 878 1252 881 1258
rect 902 1251 905 1318
rect 898 1248 905 1251
rect 886 1232 889 1248
rect 898 1238 902 1241
rect 910 1222 913 1278
rect 918 1252 921 1268
rect 870 1152 873 1188
rect 878 1162 881 1218
rect 906 1168 910 1171
rect 886 1162 889 1168
rect 918 1162 921 1228
rect 926 1212 929 1348
rect 942 1332 945 1438
rect 998 1362 1001 1388
rect 1062 1372 1065 1388
rect 1174 1362 1177 1368
rect 1190 1362 1193 1368
rect 1294 1362 1297 1368
rect 1042 1358 1046 1361
rect 1162 1358 1166 1361
rect 1218 1358 1222 1361
rect 1314 1358 1318 1361
rect 1110 1352 1113 1358
rect 1118 1352 1121 1358
rect 1230 1352 1233 1358
rect 1262 1352 1265 1358
rect 954 1348 958 1351
rect 1066 1348 1070 1351
rect 1014 1342 1017 1348
rect 970 1338 974 1341
rect 938 1328 942 1331
rect 970 1308 977 1311
rect 974 1292 977 1308
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 997 1303 1000 1307
rect 1022 1282 1025 1318
rect 1030 1292 1033 1338
rect 1046 1332 1049 1338
rect 1086 1332 1089 1338
rect 1054 1322 1057 1328
rect 1094 1322 1097 1348
rect 1126 1341 1129 1348
rect 1122 1338 1129 1341
rect 1134 1322 1137 1338
rect 1166 1332 1169 1338
rect 1174 1322 1177 1348
rect 1194 1338 1198 1341
rect 1206 1322 1209 1348
rect 1290 1338 1294 1341
rect 1314 1338 1318 1341
rect 1038 1282 1041 1318
rect 1062 1282 1065 1318
rect 1094 1282 1097 1318
rect 1158 1292 1161 1318
rect 1230 1292 1233 1328
rect 1262 1322 1265 1338
rect 1334 1331 1337 1398
rect 1350 1342 1353 1438
rect 1358 1372 1361 1378
rect 1358 1342 1361 1348
rect 1346 1338 1350 1341
rect 1334 1328 1342 1331
rect 946 1278 950 1281
rect 958 1272 961 1278
rect 966 1268 974 1271
rect 966 1261 969 1268
rect 962 1258 969 1261
rect 974 1222 977 1258
rect 1014 1252 1017 1278
rect 1098 1268 1102 1271
rect 1202 1268 1206 1271
rect 1070 1262 1073 1268
rect 1118 1262 1121 1268
rect 1186 1258 1190 1261
rect 1086 1252 1089 1258
rect 1142 1252 1145 1258
rect 1154 1248 1158 1251
rect 1038 1242 1041 1248
rect 1054 1242 1057 1248
rect 1130 1238 1134 1241
rect 1142 1232 1145 1238
rect 926 1192 929 1198
rect 934 1181 937 1218
rect 926 1178 937 1181
rect 794 1138 798 1141
rect 850 1138 854 1141
rect 822 1132 825 1138
rect 858 1118 862 1121
rect 766 1092 769 1118
rect 782 1041 785 1118
rect 790 1062 793 1068
rect 798 1062 801 1118
rect 830 1081 833 1118
rect 822 1078 833 1081
rect 850 1078 854 1081
rect 782 1038 790 1041
rect 806 1032 809 1048
rect 822 1042 825 1078
rect 830 1062 833 1068
rect 838 1052 841 1058
rect 850 1048 854 1051
rect 834 1018 838 1021
rect 698 948 710 951
rect 702 882 705 888
rect 686 872 689 878
rect 670 868 681 871
rect 650 858 654 861
rect 574 852 577 858
rect 582 842 585 858
rect 598 852 601 858
rect 662 842 665 848
rect 678 842 681 868
rect 690 858 694 861
rect 686 842 689 848
rect 642 838 646 841
rect 654 838 662 841
rect 526 792 529 838
rect 526 742 529 788
rect 566 762 569 838
rect 590 802 593 818
rect 638 802 641 818
rect 594 768 606 771
rect 554 748 558 751
rect 574 742 577 748
rect 582 742 585 768
rect 614 752 617 798
rect 630 771 633 798
rect 630 768 638 771
rect 622 762 625 768
rect 654 762 657 838
rect 670 772 673 798
rect 686 762 689 838
rect 694 792 697 798
rect 710 772 713 878
rect 718 852 721 958
rect 726 932 729 978
rect 766 962 769 1018
rect 862 1002 865 1068
rect 886 1062 889 1158
rect 894 1152 897 1158
rect 918 1141 921 1158
rect 926 1152 929 1178
rect 938 1168 942 1171
rect 950 1152 953 1208
rect 974 1172 977 1218
rect 982 1162 985 1168
rect 998 1162 1001 1218
rect 1142 1182 1145 1198
rect 1114 1168 1118 1171
rect 1026 1158 1030 1161
rect 1130 1158 1134 1161
rect 918 1138 926 1141
rect 894 1052 897 1118
rect 902 1062 905 1068
rect 910 1052 913 1138
rect 918 1072 921 1078
rect 874 1048 878 1051
rect 914 1048 918 1051
rect 874 1038 878 1041
rect 890 1038 894 1041
rect 926 1032 929 1138
rect 942 1072 945 1078
rect 934 1032 937 1068
rect 950 1062 953 1148
rect 1094 1142 1097 1158
rect 1102 1152 1105 1158
rect 974 1092 977 1138
rect 1018 1128 1022 1131
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 997 1103 1000 1107
rect 970 1078 974 1081
rect 774 962 777 978
rect 786 968 793 971
rect 734 952 737 958
rect 742 952 745 958
rect 726 871 729 928
rect 734 882 737 948
rect 726 868 734 871
rect 742 862 745 918
rect 758 862 761 868
rect 766 852 769 958
rect 778 948 782 951
rect 790 902 793 968
rect 798 952 801 958
rect 798 882 801 928
rect 806 882 809 968
rect 818 938 822 941
rect 830 932 833 968
rect 838 952 841 958
rect 846 942 849 998
rect 862 992 865 998
rect 854 982 857 988
rect 886 972 889 1018
rect 926 982 929 1028
rect 934 1012 937 1028
rect 910 972 913 978
rect 926 962 929 978
rect 950 962 953 1058
rect 966 992 969 1078
rect 1006 1071 1009 1098
rect 1002 1068 1009 1071
rect 1014 1072 1017 1078
rect 1014 1051 1017 1058
rect 1014 1048 1022 1051
rect 858 958 862 961
rect 818 928 822 931
rect 822 892 825 898
rect 838 882 841 928
rect 846 912 849 928
rect 870 912 873 958
rect 902 952 905 958
rect 934 952 937 958
rect 982 952 985 958
rect 882 948 886 951
rect 922 948 926 951
rect 954 938 958 941
rect 838 872 841 878
rect 794 868 798 871
rect 774 862 777 868
rect 862 862 865 868
rect 870 862 873 908
rect 878 872 881 918
rect 930 878 934 881
rect 898 858 910 861
rect 838 842 841 848
rect 738 838 750 841
rect 734 771 737 778
rect 730 768 737 771
rect 742 772 745 818
rect 790 792 793 808
rect 786 768 790 771
rect 802 768 806 771
rect 710 762 713 768
rect 538 738 542 741
rect 550 738 558 741
rect 634 738 638 741
rect 462 722 465 728
rect 226 668 230 671
rect 250 668 254 671
rect 258 648 262 651
rect 214 592 217 648
rect 150 572 153 578
rect 138 568 142 571
rect 162 568 166 571
rect 86 562 89 568
rect 110 562 113 568
rect 70 552 73 558
rect 102 552 105 558
rect 118 552 121 568
rect 126 562 129 568
rect 174 562 177 568
rect 238 562 241 618
rect 270 602 273 648
rect 286 642 289 648
rect 278 622 281 628
rect 294 622 297 658
rect 302 642 305 648
rect 318 632 321 638
rect 326 622 329 658
rect 334 652 337 688
rect 358 652 361 658
rect 374 651 377 668
rect 438 662 441 668
rect 370 648 377 651
rect 390 658 398 661
rect 366 642 369 648
rect 346 628 350 631
rect 294 592 297 598
rect 318 592 321 618
rect 266 568 270 571
rect 322 568 326 571
rect 342 562 345 598
rect 314 558 321 561
rect 338 558 342 561
rect 90 548 94 551
rect 58 538 62 541
rect 46 522 49 528
rect 86 492 89 538
rect 6 482 9 488
rect 126 482 129 548
rect 94 472 97 478
rect 6 432 9 468
rect 30 462 33 468
rect 42 458 46 461
rect 54 402 57 468
rect 118 462 121 468
rect 78 452 81 458
rect 126 452 129 478
rect 134 452 137 558
rect 158 542 161 548
rect 142 462 145 518
rect 150 492 153 528
rect 166 502 169 558
rect 182 542 185 548
rect 222 542 225 548
rect 294 542 297 548
rect 266 538 270 541
rect 166 462 169 468
rect 70 422 73 448
rect 102 438 110 441
rect 46 392 49 398
rect 70 352 73 398
rect 102 392 105 438
rect 118 432 121 448
rect 134 392 137 448
rect 142 392 145 438
rect 118 382 121 388
rect 150 381 153 438
rect 174 392 177 538
rect 182 432 185 468
rect 190 412 193 478
rect 198 452 201 498
rect 206 492 209 538
rect 234 528 238 531
rect 274 528 278 531
rect 214 462 217 518
rect 286 482 289 498
rect 294 492 297 538
rect 262 462 265 468
rect 242 458 246 461
rect 142 378 153 381
rect 94 362 97 368
rect 118 362 121 378
rect 130 368 134 371
rect 106 358 110 361
rect 10 348 14 351
rect 26 348 30 351
rect 50 348 54 351
rect 6 282 9 288
rect 6 152 9 158
rect 14 152 17 348
rect 70 342 73 348
rect 94 342 97 348
rect 78 332 81 338
rect 22 322 25 328
rect 78 322 81 328
rect 22 282 25 318
rect 42 278 46 281
rect 38 272 41 278
rect 54 272 57 298
rect 126 292 129 348
rect 90 258 94 261
rect 70 252 73 258
rect 102 252 105 268
rect 38 242 41 248
rect 126 242 129 258
rect 134 252 137 358
rect 142 292 145 378
rect 150 362 153 368
rect 166 362 169 388
rect 186 368 190 371
rect 198 362 201 448
rect 206 442 209 458
rect 230 452 233 458
rect 214 442 217 448
rect 194 358 198 361
rect 206 352 209 388
rect 230 381 233 448
rect 250 438 254 441
rect 238 432 241 438
rect 278 412 281 468
rect 310 452 313 508
rect 318 492 321 558
rect 350 552 353 558
rect 338 548 342 551
rect 358 492 361 638
rect 390 632 393 658
rect 446 652 449 698
rect 462 672 465 678
rect 458 648 462 651
rect 398 642 401 648
rect 394 618 398 621
rect 406 572 409 638
rect 414 602 417 618
rect 414 562 417 598
rect 422 592 425 628
rect 446 592 449 638
rect 454 592 457 638
rect 366 532 369 538
rect 334 472 337 488
rect 366 482 369 488
rect 374 482 377 528
rect 382 502 385 528
rect 390 492 393 558
rect 422 542 425 548
rect 406 532 409 538
rect 430 492 433 568
rect 454 492 457 568
rect 462 562 465 638
rect 470 632 473 658
rect 502 641 505 718
rect 550 712 553 738
rect 614 732 617 738
rect 646 732 649 748
rect 678 732 681 748
rect 686 742 689 758
rect 718 752 721 768
rect 814 762 817 798
rect 826 768 830 771
rect 838 752 841 778
rect 846 762 849 858
rect 878 852 881 858
rect 858 838 862 841
rect 870 802 873 848
rect 894 842 897 848
rect 926 822 929 868
rect 942 852 945 858
rect 886 812 889 818
rect 854 762 857 798
rect 934 782 937 788
rect 898 778 902 781
rect 870 762 873 768
rect 886 762 889 768
rect 758 742 761 748
rect 806 742 809 748
rect 862 742 865 748
rect 770 738 774 741
rect 826 738 830 741
rect 558 682 561 728
rect 614 682 617 688
rect 534 672 537 678
rect 558 672 561 678
rect 518 662 521 668
rect 550 662 553 668
rect 502 638 510 641
rect 518 632 521 638
rect 526 622 529 648
rect 472 603 474 607
rect 478 603 481 607
rect 485 603 488 607
rect 526 602 529 618
rect 550 612 553 658
rect 562 628 566 631
rect 574 611 577 638
rect 582 622 585 658
rect 594 648 598 651
rect 574 608 585 611
rect 530 588 534 591
rect 494 562 497 578
rect 502 572 505 578
rect 514 568 518 571
rect 526 568 534 571
rect 462 542 465 548
rect 494 492 497 558
rect 502 552 505 558
rect 502 492 505 508
rect 526 492 529 568
rect 550 562 553 578
rect 542 492 545 548
rect 370 478 374 481
rect 342 472 345 478
rect 398 472 401 478
rect 418 468 422 471
rect 374 462 377 468
rect 362 448 366 451
rect 294 442 297 448
rect 318 422 321 448
rect 374 432 377 458
rect 242 388 246 391
rect 230 378 241 381
rect 226 368 230 371
rect 158 291 161 338
rect 182 292 185 348
rect 214 342 217 368
rect 238 362 241 378
rect 250 368 254 371
rect 262 352 265 358
rect 242 348 246 351
rect 158 288 169 291
rect 158 262 161 278
rect 166 252 169 288
rect 230 272 233 348
rect 294 342 297 408
rect 382 392 385 468
rect 414 382 417 388
rect 422 382 425 458
rect 438 452 441 468
rect 446 442 449 448
rect 454 392 457 478
rect 462 472 465 488
rect 498 478 502 481
rect 474 468 478 471
rect 472 403 474 407
rect 478 403 481 407
rect 485 403 488 407
rect 510 392 513 478
rect 550 472 553 558
rect 566 542 569 548
rect 574 512 577 568
rect 582 492 585 608
rect 590 562 593 638
rect 606 632 609 638
rect 534 462 537 468
rect 518 442 521 448
rect 518 392 521 428
rect 542 392 545 438
rect 558 412 561 468
rect 566 462 569 478
rect 586 468 590 471
rect 574 442 577 448
rect 550 392 553 398
rect 590 382 593 458
rect 598 392 601 548
rect 390 372 393 378
rect 318 362 321 368
rect 350 362 353 368
rect 374 362 377 368
rect 310 352 313 358
rect 282 338 286 341
rect 246 292 249 338
rect 318 332 321 338
rect 282 328 286 331
rect 370 328 374 331
rect 270 282 273 288
rect 238 262 241 268
rect 82 238 86 241
rect 134 238 142 241
rect 94 232 97 238
rect 38 182 41 228
rect 118 222 121 238
rect 22 92 25 168
rect 38 142 41 178
rect 54 132 57 138
rect 6 82 9 88
rect 30 71 33 128
rect 62 92 65 208
rect 78 192 81 218
rect 134 192 137 238
rect 70 162 73 168
rect 86 162 89 188
rect 90 148 94 151
rect 78 142 81 148
rect 46 72 49 78
rect 30 68 38 71
rect 38 62 41 68
rect 86 62 89 118
rect 110 102 113 118
rect 94 72 97 78
rect 118 72 121 188
rect 126 141 129 168
rect 134 152 137 168
rect 142 162 145 218
rect 150 212 153 238
rect 166 222 169 248
rect 182 212 185 258
rect 206 252 209 258
rect 214 252 217 258
rect 262 252 265 268
rect 270 262 273 268
rect 294 252 297 258
rect 194 238 198 241
rect 234 238 238 241
rect 166 192 169 208
rect 126 138 137 141
rect 134 92 137 138
rect 158 132 161 168
rect 178 158 182 161
rect 170 148 182 151
rect 198 142 201 148
rect 206 122 209 128
rect 150 82 153 88
rect 158 82 161 108
rect 166 72 169 98
rect 178 88 182 91
rect 198 62 201 78
rect 206 72 209 98
rect 214 92 217 238
rect 254 222 257 248
rect 230 162 233 188
rect 238 172 241 178
rect 226 128 230 131
rect 246 92 249 168
rect 262 162 265 248
rect 302 242 305 318
rect 318 282 321 328
rect 350 312 353 328
rect 382 292 385 348
rect 398 292 401 368
rect 346 278 350 281
rect 362 278 366 281
rect 322 268 326 271
rect 310 242 313 268
rect 282 238 286 241
rect 318 192 321 218
rect 334 182 337 188
rect 358 162 361 268
rect 366 192 369 268
rect 306 158 313 161
rect 270 152 273 158
rect 258 148 262 151
rect 290 138 294 141
rect 294 102 297 128
rect 242 78 246 81
rect 262 62 265 98
rect 294 72 297 98
rect 310 92 313 158
rect 318 102 321 148
rect 326 142 329 148
rect 342 92 345 128
rect 350 92 353 158
rect 374 152 377 278
rect 390 272 393 278
rect 406 272 409 338
rect 394 268 398 271
rect 422 262 425 378
rect 458 368 462 371
rect 554 368 558 371
rect 442 358 446 361
rect 454 342 457 348
rect 434 328 438 331
rect 446 262 449 298
rect 458 288 465 291
rect 462 282 465 288
rect 438 252 441 258
rect 406 192 409 248
rect 454 192 457 278
rect 470 272 473 328
rect 486 292 489 368
rect 510 362 513 368
rect 522 358 526 361
rect 578 358 582 361
rect 570 348 574 351
rect 590 351 593 368
rect 606 362 609 598
rect 614 592 617 658
rect 622 652 625 698
rect 678 682 681 718
rect 702 702 705 738
rect 718 732 721 738
rect 726 702 729 728
rect 726 682 729 698
rect 742 681 745 718
rect 750 712 753 738
rect 754 688 758 691
rect 782 682 785 728
rect 806 692 809 728
rect 742 678 758 681
rect 762 678 766 681
rect 786 678 790 681
rect 830 672 833 708
rect 690 668 694 671
rect 810 668 814 671
rect 850 668 854 671
rect 702 662 705 668
rect 734 662 737 668
rect 674 658 678 661
rect 630 652 633 658
rect 638 652 641 658
rect 654 652 657 658
rect 686 652 689 658
rect 650 638 654 641
rect 622 562 625 598
rect 630 592 633 618
rect 662 592 665 638
rect 670 632 673 638
rect 678 632 681 638
rect 630 542 633 548
rect 638 512 641 568
rect 654 562 657 578
rect 674 568 678 571
rect 718 562 721 568
rect 674 548 686 551
rect 702 542 705 548
rect 630 492 633 508
rect 646 492 649 538
rect 702 492 705 508
rect 614 482 617 488
rect 678 482 681 488
rect 710 482 713 528
rect 742 511 745 668
rect 766 662 769 668
rect 758 532 761 538
rect 750 522 753 528
rect 742 508 753 511
rect 666 478 670 481
rect 694 472 697 478
rect 742 472 745 478
rect 622 462 625 468
rect 662 462 665 468
rect 734 462 737 468
rect 614 352 617 358
rect 582 348 593 351
rect 510 332 513 338
rect 538 328 542 331
rect 494 322 497 328
rect 510 292 513 298
rect 566 292 569 328
rect 530 288 534 291
rect 510 282 513 288
rect 574 282 577 318
rect 582 292 585 348
rect 598 341 601 348
rect 590 338 601 341
rect 538 278 542 281
rect 518 272 521 278
rect 590 272 593 338
rect 598 292 601 328
rect 622 282 625 458
rect 726 452 729 458
rect 642 448 646 451
rect 714 448 721 451
rect 654 392 657 448
rect 614 272 617 278
rect 466 268 470 271
rect 472 203 474 207
rect 478 203 481 207
rect 485 203 488 207
rect 390 112 393 128
rect 362 78 366 81
rect 274 68 278 71
rect 318 62 321 68
rect 82 58 86 61
rect 238 52 241 58
rect 74 48 78 51
rect 146 48 150 51
rect 250 48 254 51
rect 298 48 302 51
rect 102 42 105 48
rect 118 42 121 48
rect 278 42 281 48
rect 318 32 321 48
rect 334 22 337 78
rect 370 68 374 71
rect 390 62 393 68
rect 398 62 401 128
rect 406 92 409 178
rect 494 152 497 268
rect 502 192 505 248
rect 534 192 537 248
rect 550 242 553 268
rect 566 192 569 268
rect 622 222 625 268
rect 630 262 633 338
rect 654 332 657 368
rect 666 358 670 361
rect 678 342 681 438
rect 718 392 721 448
rect 726 362 729 418
rect 698 348 702 351
rect 686 332 689 348
rect 710 342 713 358
rect 726 342 729 348
rect 742 332 745 338
rect 638 282 641 328
rect 646 292 649 328
rect 662 322 665 328
rect 678 312 681 318
rect 678 282 681 308
rect 686 272 689 328
rect 710 322 713 328
rect 742 281 745 328
rect 750 312 753 508
rect 766 482 769 538
rect 774 502 777 668
rect 862 662 865 718
rect 870 682 873 748
rect 894 702 897 768
rect 918 752 921 758
rect 906 748 910 751
rect 934 742 937 778
rect 942 732 945 808
rect 950 792 953 908
rect 984 903 986 907
rect 990 903 993 907
rect 997 903 1000 907
rect 978 878 982 881
rect 1002 878 1006 881
rect 1014 872 1017 1048
rect 1030 1042 1033 1118
rect 1038 1062 1041 1108
rect 1046 1082 1049 1138
rect 1054 1122 1057 1128
rect 1046 1052 1049 1078
rect 1070 1062 1073 1068
rect 1042 1018 1046 1021
rect 1046 972 1049 998
rect 1054 962 1057 1018
rect 1022 942 1025 948
rect 1030 931 1033 958
rect 1038 952 1041 958
rect 1022 928 1033 931
rect 1022 892 1025 928
rect 1038 862 1041 918
rect 986 828 990 831
rect 950 762 953 788
rect 1014 772 1017 828
rect 1022 792 1025 818
rect 1030 802 1033 848
rect 1046 842 1049 848
rect 970 768 982 771
rect 998 762 1001 768
rect 958 752 961 758
rect 1010 748 1014 751
rect 1030 742 1033 748
rect 958 732 961 738
rect 882 668 886 671
rect 870 662 873 668
rect 818 658 822 661
rect 850 658 854 661
rect 790 552 793 618
rect 798 592 801 648
rect 894 642 897 668
rect 902 662 905 688
rect 910 682 913 718
rect 914 678 918 681
rect 926 672 929 678
rect 942 672 945 728
rect 966 712 969 728
rect 950 692 953 698
rect 966 682 969 708
rect 984 703 986 707
rect 990 703 993 707
rect 997 703 1000 707
rect 1038 692 1041 818
rect 1046 742 1049 818
rect 1054 812 1057 948
rect 1062 942 1065 988
rect 1070 982 1073 1048
rect 1078 1042 1081 1118
rect 1086 1092 1089 1138
rect 1102 1112 1105 1118
rect 1086 1052 1089 1078
rect 1134 1072 1137 1148
rect 1142 1142 1145 1178
rect 1158 1162 1161 1168
rect 1150 1091 1153 1128
rect 1174 1112 1177 1258
rect 1186 1248 1190 1251
rect 1198 1242 1201 1258
rect 1222 1242 1225 1278
rect 1230 1262 1233 1268
rect 1246 1262 1249 1318
rect 1246 1242 1249 1248
rect 1254 1232 1257 1258
rect 1270 1241 1273 1318
rect 1266 1238 1273 1241
rect 1278 1242 1281 1248
rect 1286 1232 1289 1258
rect 1294 1242 1297 1318
rect 1318 1282 1321 1318
rect 1318 1262 1321 1268
rect 1314 1248 1318 1251
rect 1202 1158 1206 1161
rect 1186 1128 1190 1131
rect 1198 1122 1201 1128
rect 1146 1088 1153 1091
rect 1142 1082 1145 1088
rect 1214 1081 1217 1128
rect 1222 1102 1225 1138
rect 1214 1078 1222 1081
rect 1174 1072 1177 1078
rect 1190 1072 1193 1078
rect 1222 1072 1225 1078
rect 1118 1062 1121 1068
rect 1098 1058 1102 1061
rect 1070 931 1073 978
rect 1062 928 1073 931
rect 1062 852 1065 928
rect 1070 862 1073 868
rect 1066 848 1070 851
rect 1078 842 1081 918
rect 1086 911 1089 1048
rect 1150 1042 1153 1048
rect 1106 1038 1110 1041
rect 1094 1002 1097 1018
rect 1134 942 1137 948
rect 1094 922 1097 928
rect 1102 922 1105 928
rect 1086 908 1097 911
rect 1094 872 1097 908
rect 1102 882 1105 918
rect 1070 832 1073 838
rect 1054 732 1057 808
rect 1094 772 1097 868
rect 1110 862 1113 868
rect 1102 852 1105 858
rect 1118 832 1121 918
rect 1134 912 1137 938
rect 1134 872 1137 908
rect 1142 902 1145 998
rect 1198 992 1201 1058
rect 1230 1041 1233 1218
rect 1238 1182 1241 1188
rect 1250 1168 1254 1171
rect 1258 1158 1262 1161
rect 1246 1082 1249 1138
rect 1270 1072 1273 1218
rect 1302 1182 1305 1218
rect 1278 1162 1281 1168
rect 1286 1152 1289 1178
rect 1310 1172 1313 1248
rect 1326 1242 1329 1288
rect 1342 1262 1345 1268
rect 1318 1232 1321 1238
rect 1322 1168 1326 1171
rect 1298 1158 1302 1161
rect 1310 1142 1313 1148
rect 1286 1132 1289 1138
rect 1334 1122 1337 1158
rect 1342 1142 1345 1238
rect 1350 1162 1353 1338
rect 1366 1331 1369 1438
rect 1374 1362 1377 1368
rect 1402 1358 1406 1361
rect 1434 1358 1438 1361
rect 1382 1342 1385 1348
rect 1358 1328 1369 1331
rect 1358 1272 1361 1328
rect 1390 1322 1393 1348
rect 1434 1338 1438 1341
rect 1454 1322 1457 1338
rect 1370 1278 1374 1281
rect 1414 1272 1417 1318
rect 1438 1292 1441 1318
rect 1430 1271 1433 1278
rect 1430 1268 1438 1271
rect 1358 1202 1361 1268
rect 1374 1242 1377 1248
rect 1382 1232 1385 1258
rect 1390 1242 1393 1268
rect 1418 1258 1422 1261
rect 1422 1242 1425 1248
rect 1414 1232 1417 1238
rect 1406 1222 1409 1228
rect 1358 1172 1361 1178
rect 1274 1058 1278 1061
rect 1290 1058 1294 1061
rect 1258 1048 1262 1051
rect 1302 1042 1305 1068
rect 1310 1062 1313 1118
rect 1326 1082 1329 1088
rect 1334 1062 1337 1118
rect 1342 1072 1345 1108
rect 1350 1082 1353 1158
rect 1358 1142 1361 1148
rect 1366 1132 1369 1168
rect 1382 1162 1385 1218
rect 1430 1192 1433 1268
rect 1446 1222 1449 1228
rect 1462 1192 1465 1238
rect 1438 1162 1441 1168
rect 1398 1152 1401 1158
rect 1398 1142 1401 1148
rect 1386 1138 1390 1141
rect 1406 1132 1409 1138
rect 1402 1078 1406 1081
rect 1342 1062 1345 1068
rect 1366 1062 1369 1068
rect 1230 1038 1238 1041
rect 1274 1038 1278 1041
rect 1218 1018 1222 1021
rect 1186 968 1190 971
rect 1150 932 1153 968
rect 1174 962 1177 968
rect 1206 962 1209 1008
rect 1246 962 1249 1018
rect 1254 992 1257 1008
rect 1202 948 1206 951
rect 1242 948 1246 951
rect 1262 942 1265 948
rect 1218 938 1222 941
rect 1174 932 1177 938
rect 1294 931 1297 1018
rect 1290 928 1297 931
rect 1302 942 1305 968
rect 1142 882 1145 898
rect 1206 882 1209 908
rect 1214 872 1217 928
rect 1238 892 1241 898
rect 1254 892 1257 918
rect 1270 902 1273 928
rect 1238 882 1241 888
rect 1254 882 1257 888
rect 1294 882 1297 918
rect 1302 872 1305 938
rect 1318 932 1321 1048
rect 1326 972 1329 1018
rect 1334 962 1337 1058
rect 1374 1052 1377 1078
rect 1382 1072 1385 1078
rect 1402 1068 1406 1071
rect 1350 1042 1353 1048
rect 1358 1022 1361 1038
rect 1374 992 1377 1048
rect 1398 1032 1401 1068
rect 1414 1062 1417 1148
rect 1438 1142 1441 1148
rect 1450 1138 1454 1141
rect 1442 1128 1446 1131
rect 1462 1072 1465 1138
rect 1470 1132 1473 1138
rect 1470 1082 1473 1088
rect 1434 1058 1438 1061
rect 1446 1052 1449 1058
rect 1418 1048 1422 1051
rect 1342 962 1345 988
rect 1362 968 1366 971
rect 1326 952 1329 958
rect 1318 912 1321 918
rect 1194 868 1198 871
rect 1290 868 1294 871
rect 1182 862 1185 868
rect 1162 858 1166 861
rect 1146 848 1150 851
rect 1170 838 1174 841
rect 1158 792 1161 818
rect 1198 812 1201 868
rect 1310 862 1313 868
rect 1334 852 1337 958
rect 1342 952 1345 958
rect 1374 952 1377 958
rect 1354 948 1358 951
rect 1390 932 1393 938
rect 1398 932 1401 938
rect 1406 932 1409 988
rect 1322 848 1326 851
rect 1214 842 1217 848
rect 1286 842 1289 848
rect 1342 842 1345 858
rect 1350 852 1353 858
rect 1358 852 1361 928
rect 1406 922 1409 928
rect 1366 862 1369 908
rect 1298 838 1302 841
rect 1330 838 1334 841
rect 1310 832 1313 838
rect 1326 802 1329 818
rect 1270 792 1273 798
rect 1290 788 1294 791
rect 1154 768 1158 771
rect 1298 768 1302 771
rect 1086 751 1089 758
rect 1118 752 1121 758
rect 1214 752 1217 758
rect 1254 752 1257 768
rect 1310 752 1313 798
rect 1318 772 1321 788
rect 1358 772 1361 848
rect 1374 842 1377 848
rect 1390 842 1393 848
rect 1398 842 1401 878
rect 1406 852 1409 858
rect 1414 852 1417 1048
rect 1434 1038 1438 1041
rect 1426 1018 1430 1021
rect 1454 992 1457 1038
rect 1470 1002 1473 1078
rect 1434 968 1438 971
rect 1442 958 1446 961
rect 1458 938 1462 941
rect 1446 882 1449 938
rect 1478 932 1481 968
rect 1422 872 1425 878
rect 1318 762 1321 768
rect 1118 682 1121 748
rect 1182 722 1185 747
rect 1334 742 1337 758
rect 1358 742 1361 748
rect 1238 718 1246 721
rect 1206 692 1209 708
rect 1230 692 1233 698
rect 990 632 993 668
rect 1054 662 1057 678
rect 1118 663 1121 668
rect 1022 652 1025 659
rect 1238 662 1241 718
rect 1258 668 1262 671
rect 1270 662 1273 668
rect 1258 658 1262 661
rect 1214 642 1217 658
rect 1278 652 1281 738
rect 1302 692 1305 718
rect 1310 692 1313 738
rect 1290 678 1294 681
rect 1286 662 1289 668
rect 1294 662 1297 668
rect 1090 638 1094 641
rect 842 618 846 621
rect 838 551 841 558
rect 870 552 873 628
rect 918 562 921 618
rect 934 572 937 618
rect 946 558 950 561
rect 994 558 998 561
rect 1014 542 1017 608
rect 1302 592 1305 668
rect 1114 568 1118 571
rect 1154 568 1158 571
rect 1102 562 1105 568
rect 1166 562 1169 578
rect 1238 572 1241 578
rect 1226 568 1230 571
rect 1258 568 1262 571
rect 1214 562 1217 568
rect 1122 558 1126 561
rect 1178 558 1185 561
rect 1066 548 1070 551
rect 1154 548 1158 551
rect 794 538 798 541
rect 914 538 918 541
rect 962 538 966 541
rect 1018 538 1022 541
rect 1042 538 1046 541
rect 758 472 761 478
rect 782 442 785 518
rect 806 512 809 538
rect 942 522 945 528
rect 806 492 809 498
rect 790 462 793 468
rect 822 462 825 468
rect 830 452 833 508
rect 846 472 849 478
rect 902 462 905 518
rect 838 458 846 461
rect 882 458 886 461
rect 794 448 798 451
rect 810 438 814 441
rect 758 301 761 438
rect 790 412 793 418
rect 790 362 793 368
rect 806 362 809 368
rect 774 352 777 358
rect 814 352 817 408
rect 830 362 833 448
rect 838 432 841 458
rect 870 452 873 458
rect 838 392 841 398
rect 738 278 745 281
rect 750 298 761 301
rect 766 332 769 348
rect 790 342 793 348
rect 650 268 654 271
rect 646 252 649 258
rect 702 252 705 258
rect 694 232 697 238
rect 702 232 705 238
rect 658 228 662 231
rect 682 188 686 191
rect 518 152 521 158
rect 418 148 422 151
rect 442 138 446 141
rect 422 122 425 128
rect 430 72 433 128
rect 462 82 465 128
rect 486 92 489 148
rect 554 138 558 141
rect 530 128 534 131
rect 518 72 521 98
rect 526 92 529 128
rect 542 72 545 128
rect 574 112 577 128
rect 598 122 601 148
rect 434 68 438 71
rect 458 68 462 71
rect 550 62 553 98
rect 574 92 577 108
rect 570 78 574 81
rect 418 48 422 51
rect 342 42 345 48
rect 438 12 441 58
rect 506 48 510 51
rect 494 32 497 38
rect 546 28 550 31
rect 454 -18 457 8
rect 472 3 474 7
rect 478 3 481 7
rect 485 3 488 7
rect 494 -18 497 28
rect 558 -18 561 78
rect 598 72 601 118
rect 614 92 617 158
rect 622 142 625 148
rect 630 142 633 158
rect 622 112 625 128
rect 622 72 625 78
rect 594 48 598 51
rect 566 42 569 48
rect 622 42 625 48
rect 630 -18 633 138
rect 646 132 649 138
rect 662 132 665 178
rect 702 172 705 188
rect 710 162 713 248
rect 718 182 721 278
rect 742 262 745 268
rect 730 248 734 251
rect 726 162 729 198
rect 750 192 753 298
rect 766 281 769 328
rect 806 292 809 348
rect 822 342 825 358
rect 766 278 774 281
rect 762 268 766 271
rect 766 238 774 241
rect 714 158 718 161
rect 710 142 713 148
rect 646 62 649 118
rect 662 91 665 128
rect 686 112 689 138
rect 710 122 713 128
rect 654 88 665 91
rect 654 -18 657 88
rect 670 82 673 88
rect 686 81 689 108
rect 686 78 694 81
rect 662 72 665 78
rect 662 52 665 58
rect 670 -18 673 78
rect 694 62 697 78
rect 710 52 713 68
rect 718 42 721 48
rect 718 -18 721 38
rect 726 12 729 158
rect 734 132 737 148
rect 742 92 745 168
rect 758 132 761 138
rect 758 82 761 128
rect 766 92 769 238
rect 782 232 785 258
rect 794 248 798 251
rect 806 232 809 238
rect 790 221 793 228
rect 786 218 793 221
rect 814 212 817 258
rect 822 202 825 338
rect 830 252 833 358
rect 838 352 841 358
rect 846 312 849 448
rect 858 438 862 441
rect 870 362 873 448
rect 918 442 921 518
rect 950 482 953 538
rect 974 532 977 538
rect 998 532 1001 538
rect 1042 528 1046 531
rect 942 472 945 478
rect 926 462 929 468
rect 890 438 894 441
rect 878 432 881 438
rect 862 342 865 348
rect 878 332 881 408
rect 918 402 921 418
rect 950 412 953 478
rect 958 441 961 518
rect 984 503 986 507
rect 990 503 993 507
rect 997 503 1000 507
rect 990 482 993 488
rect 1022 462 1025 468
rect 1030 462 1033 518
rect 1042 468 1046 471
rect 1070 462 1073 528
rect 1078 492 1081 538
rect 1098 518 1102 521
rect 1118 492 1121 538
rect 1142 532 1145 538
rect 1110 482 1113 488
rect 1134 482 1137 518
rect 1082 478 1086 481
rect 1114 468 1118 471
rect 978 458 982 461
rect 970 448 974 451
rect 958 438 966 441
rect 962 428 966 431
rect 974 392 977 408
rect 886 342 889 378
rect 914 368 918 371
rect 1006 362 1009 448
rect 1038 442 1041 448
rect 1022 422 1025 438
rect 1046 412 1049 458
rect 1078 452 1081 468
rect 1066 448 1070 451
rect 1022 362 1025 378
rect 1034 368 1038 371
rect 1078 362 1081 368
rect 930 358 934 361
rect 922 348 926 351
rect 902 342 905 348
rect 870 312 873 318
rect 838 292 841 308
rect 870 271 873 308
rect 926 282 929 288
rect 862 268 873 271
rect 830 182 833 248
rect 838 232 841 258
rect 862 252 865 268
rect 902 262 905 268
rect 850 238 857 241
rect 774 152 777 178
rect 778 128 782 131
rect 774 88 782 91
rect 742 72 745 78
rect 774 71 777 88
rect 770 68 777 71
rect 782 72 785 88
rect 738 48 742 51
rect 766 32 769 48
rect 750 -18 753 8
rect 774 -18 777 68
rect 790 42 793 138
rect 806 132 809 138
rect 806 92 809 108
rect 798 62 801 78
rect 798 -18 801 58
rect 814 -18 817 178
rect 822 112 825 168
rect 838 162 841 188
rect 846 162 849 198
rect 854 192 857 238
rect 870 232 873 258
rect 878 242 881 248
rect 862 221 865 228
rect 862 218 870 221
rect 894 212 897 248
rect 910 242 913 268
rect 934 252 937 358
rect 942 312 945 358
rect 950 352 953 358
rect 950 332 953 338
rect 990 332 993 348
rect 984 303 986 307
rect 990 303 993 307
rect 997 303 1000 307
rect 962 268 966 271
rect 942 262 945 268
rect 974 252 977 258
rect 954 248 958 251
rect 902 232 905 238
rect 830 142 833 148
rect 830 122 833 128
rect 846 92 849 138
rect 854 132 857 148
rect 862 142 865 168
rect 878 162 881 198
rect 886 192 889 208
rect 894 192 897 208
rect 934 192 937 248
rect 982 242 985 248
rect 898 168 902 171
rect 910 162 913 188
rect 958 182 961 238
rect 974 232 977 238
rect 990 192 993 268
rect 1006 212 1009 358
rect 1046 352 1049 358
rect 1026 348 1030 351
rect 1014 282 1017 308
rect 1062 272 1065 338
rect 1070 302 1073 328
rect 1078 282 1081 338
rect 1086 332 1089 468
rect 1102 462 1105 468
rect 1134 462 1137 468
rect 1146 458 1150 461
rect 1142 422 1145 448
rect 1158 442 1161 478
rect 1174 462 1177 468
rect 1170 448 1174 451
rect 1182 422 1185 558
rect 1190 532 1193 538
rect 1214 492 1217 538
rect 1238 522 1241 548
rect 1190 462 1193 468
rect 1214 462 1217 468
rect 1238 462 1241 468
rect 1246 462 1249 558
rect 1262 552 1265 558
rect 1270 552 1273 578
rect 1290 568 1294 571
rect 1310 562 1313 648
rect 1318 642 1321 678
rect 1350 652 1353 659
rect 1318 622 1321 638
rect 1282 558 1289 561
rect 1278 472 1281 478
rect 1230 452 1233 458
rect 1190 442 1193 448
rect 1202 438 1206 441
rect 1222 432 1225 448
rect 1254 442 1257 448
rect 1266 438 1270 441
rect 1150 392 1153 408
rect 1214 392 1217 418
rect 1110 332 1113 388
rect 1122 348 1126 351
rect 1134 342 1137 348
rect 1158 342 1161 378
rect 1214 362 1217 368
rect 1182 352 1185 358
rect 1186 328 1190 331
rect 1110 292 1113 328
rect 1118 312 1121 328
rect 1126 292 1129 308
rect 1086 282 1089 288
rect 1198 282 1201 338
rect 1042 268 1046 271
rect 1074 268 1078 271
rect 1046 252 1049 258
rect 1090 248 1094 251
rect 1042 238 1046 241
rect 918 172 921 178
rect 930 168 937 171
rect 886 152 889 158
rect 910 92 913 158
rect 918 142 921 148
rect 934 92 937 168
rect 958 142 961 178
rect 1006 162 1009 208
rect 1022 162 1025 178
rect 1034 168 1041 171
rect 970 148 974 151
rect 1026 148 1030 151
rect 942 132 945 138
rect 822 72 825 78
rect 830 72 833 88
rect 870 62 873 68
rect 858 48 862 51
rect 894 32 897 78
rect 926 72 929 88
rect 958 82 961 98
rect 966 92 969 128
rect 958 72 961 78
rect 906 68 910 71
rect 966 62 969 78
rect 974 61 977 148
rect 1002 128 1006 131
rect 984 103 986 107
rect 990 103 993 107
rect 997 103 1000 107
rect 1006 82 1009 98
rect 1038 92 1041 168
rect 1046 152 1049 158
rect 1066 138 1070 141
rect 1066 128 1070 131
rect 1014 82 1017 88
rect 1054 82 1057 88
rect 1078 82 1081 128
rect 1094 92 1097 118
rect 1102 102 1105 278
rect 1154 268 1158 271
rect 1114 248 1118 251
rect 1114 238 1118 241
rect 1110 162 1113 168
rect 1122 138 1126 141
rect 1046 78 1054 81
rect 974 58 982 61
rect 902 52 905 58
rect 986 48 990 51
rect 886 22 889 28
rect 918 22 921 48
rect 886 -18 889 18
rect 918 -18 921 18
rect 934 -18 937 8
rect 958 -18 961 8
rect 1006 -18 1009 78
rect 1022 -18 1025 58
rect 1046 -18 1049 78
rect 1062 32 1065 78
rect 1094 72 1097 88
rect 1110 82 1113 138
rect 1134 92 1137 268
rect 1142 242 1145 248
rect 1166 242 1169 268
rect 1174 252 1177 258
rect 1182 252 1185 258
rect 1190 242 1193 278
rect 1222 272 1225 428
rect 1238 392 1241 418
rect 1246 402 1249 438
rect 1278 422 1281 458
rect 1286 452 1289 558
rect 1298 548 1302 551
rect 1294 452 1297 498
rect 1302 492 1305 538
rect 1310 502 1313 558
rect 1318 552 1321 558
rect 1342 542 1345 548
rect 1330 538 1337 541
rect 1302 462 1305 468
rect 1326 462 1329 468
rect 1286 422 1289 448
rect 1254 381 1257 408
rect 1262 392 1265 398
rect 1246 378 1257 381
rect 1230 312 1233 368
rect 1246 362 1249 378
rect 1286 372 1289 378
rect 1254 362 1257 368
rect 1294 362 1297 448
rect 1306 438 1310 441
rect 1326 382 1329 458
rect 1334 392 1337 538
rect 1350 532 1353 638
rect 1366 551 1369 818
rect 1446 792 1449 878
rect 1478 852 1481 868
rect 1478 822 1481 848
rect 1438 782 1441 788
rect 1462 752 1465 758
rect 1382 662 1385 748
rect 1446 742 1449 748
rect 1446 692 1449 728
rect 1382 621 1385 658
rect 1438 642 1441 648
rect 1382 618 1393 621
rect 1366 548 1374 551
rect 1390 542 1393 618
rect 1470 592 1473 658
rect 1406 551 1409 558
rect 1362 538 1366 541
rect 1358 462 1361 518
rect 1406 472 1409 528
rect 1342 412 1345 458
rect 1374 452 1377 459
rect 1342 392 1345 408
rect 1274 358 1278 361
rect 1238 352 1241 358
rect 1150 232 1153 238
rect 1198 202 1201 268
rect 1214 262 1217 268
rect 1226 258 1230 261
rect 1226 248 1230 251
rect 1214 241 1217 248
rect 1214 238 1222 241
rect 1222 192 1225 198
rect 1230 192 1233 218
rect 1166 172 1169 178
rect 1154 168 1158 171
rect 1170 158 1174 161
rect 1142 152 1145 158
rect 1182 152 1185 158
rect 1198 152 1201 158
rect 1214 152 1217 188
rect 1238 172 1241 268
rect 1246 252 1249 358
rect 1294 342 1297 348
rect 1254 242 1257 278
rect 1246 192 1249 208
rect 1262 182 1265 268
rect 1270 242 1273 338
rect 1278 262 1281 268
rect 1290 258 1294 261
rect 1302 252 1305 378
rect 1346 368 1353 371
rect 1330 358 1334 361
rect 1318 342 1321 348
rect 1318 262 1321 338
rect 1298 248 1302 251
rect 1302 232 1305 238
rect 1294 201 1297 218
rect 1286 198 1297 201
rect 1286 172 1289 198
rect 1294 182 1297 188
rect 1222 152 1225 168
rect 1238 162 1241 168
rect 1162 148 1166 151
rect 1202 138 1206 141
rect 1214 92 1217 128
rect 1138 88 1142 91
rect 1182 82 1185 88
rect 1102 72 1105 78
rect 1078 62 1081 68
rect 1110 62 1113 78
rect 1158 72 1161 78
rect 1222 72 1225 138
rect 1246 92 1249 148
rect 1254 132 1257 168
rect 1270 162 1273 168
rect 1274 148 1278 151
rect 1294 92 1297 168
rect 1310 142 1313 218
rect 1334 192 1337 348
rect 1350 292 1353 368
rect 1358 362 1361 378
rect 1414 372 1417 418
rect 1370 368 1374 371
rect 1394 368 1398 371
rect 1382 362 1385 368
rect 1362 348 1366 351
rect 1342 252 1345 278
rect 1354 258 1358 261
rect 1374 242 1377 268
rect 1346 238 1350 241
rect 1362 238 1369 241
rect 1302 82 1305 128
rect 1282 78 1286 81
rect 1310 81 1313 138
rect 1318 92 1321 178
rect 1350 172 1353 208
rect 1358 192 1361 228
rect 1366 222 1369 238
rect 1330 158 1334 161
rect 1338 148 1342 151
rect 1326 142 1329 148
rect 1326 82 1329 108
rect 1342 92 1345 128
rect 1310 78 1321 81
rect 1122 68 1126 71
rect 1226 68 1230 71
rect 1306 68 1310 71
rect 1198 62 1201 68
rect 1098 58 1102 61
rect 1154 58 1158 61
rect 1250 58 1254 61
rect 1126 52 1129 58
rect 1078 22 1081 38
rect 1070 -18 1073 8
rect 1142 -18 1145 58
rect 1262 52 1265 58
rect 1170 48 1174 51
rect 1202 48 1206 51
rect 1242 48 1246 51
rect 1278 42 1281 68
rect 1290 48 1294 51
rect 1238 32 1241 38
rect 1166 22 1169 28
rect 454 -22 458 -18
rect 494 -22 498 -18
rect 558 -22 562 -18
rect 630 -22 634 -18
rect 654 -22 658 -18
rect 670 -22 674 -18
rect 718 -22 722 -18
rect 750 -22 754 -18
rect 774 -22 778 -18
rect 798 -22 802 -18
rect 814 -22 818 -18
rect 886 -22 890 -18
rect 918 -22 922 -18
rect 934 -22 938 -18
rect 958 -22 962 -18
rect 1006 -22 1010 -18
rect 1022 -22 1026 -18
rect 1046 -22 1050 -18
rect 1070 -22 1074 -18
rect 1142 -22 1146 -18
rect 1270 -19 1274 -18
rect 1278 -19 1281 38
rect 1270 -22 1281 -19
rect 1302 -18 1305 68
rect 1318 -18 1321 78
rect 1350 62 1353 158
rect 1366 142 1369 198
rect 1374 192 1377 228
rect 1382 212 1385 218
rect 1382 192 1385 198
rect 1390 162 1393 318
rect 1398 192 1401 358
rect 1406 352 1409 368
rect 1414 362 1417 368
rect 1422 362 1425 388
rect 1406 322 1409 328
rect 1406 282 1409 318
rect 1414 282 1417 358
rect 1422 348 1430 351
rect 1422 281 1425 348
rect 1438 341 1441 368
rect 1430 338 1441 341
rect 1430 292 1433 338
rect 1422 278 1433 281
rect 1414 242 1417 268
rect 1422 152 1425 248
rect 1410 148 1414 151
rect 1366 132 1369 138
rect 1386 128 1390 131
rect 1370 78 1374 81
rect 1382 71 1385 98
rect 1390 92 1393 118
rect 1430 92 1433 278
rect 1446 252 1449 418
rect 1454 372 1457 378
rect 1470 342 1473 428
rect 1474 338 1478 341
rect 1402 88 1406 91
rect 1426 78 1430 81
rect 1446 72 1449 238
rect 1454 82 1457 298
rect 1470 282 1473 288
rect 1474 278 1478 281
rect 1474 168 1478 171
rect 1478 82 1481 108
rect 1378 68 1385 71
rect 1418 68 1422 71
rect 1354 48 1358 51
rect 1338 38 1342 41
rect 1302 -22 1306 -18
rect 1318 -22 1322 -18
<< m3contact >>
rect 54 1358 58 1362
rect 30 1338 34 1342
rect 62 1338 66 1342
rect 6 1328 10 1332
rect 6 1318 10 1322
rect 6 1308 10 1312
rect 94 1358 98 1362
rect 118 1358 122 1362
rect 142 1358 146 1362
rect 102 1338 106 1342
rect 150 1338 154 1342
rect 86 1328 90 1332
rect 38 1268 42 1272
rect 30 1248 34 1252
rect 62 1308 66 1312
rect 46 1248 50 1252
rect 54 1248 58 1252
rect 38 1188 42 1192
rect 14 1178 18 1182
rect 38 1178 42 1182
rect 46 1158 50 1162
rect 214 1358 218 1362
rect 342 1408 346 1412
rect 474 1403 478 1407
rect 481 1403 485 1407
rect 526 1398 530 1402
rect 422 1388 426 1392
rect 342 1378 346 1382
rect 270 1368 274 1372
rect 366 1368 370 1372
rect 510 1378 514 1382
rect 262 1358 266 1362
rect 438 1358 442 1362
rect 454 1358 458 1362
rect 478 1358 482 1362
rect 198 1348 202 1352
rect 222 1348 226 1352
rect 238 1348 242 1352
rect 246 1348 250 1352
rect 182 1328 186 1332
rect 118 1308 122 1312
rect 142 1298 146 1302
rect 126 1278 130 1282
rect 110 1268 114 1272
rect 118 1268 122 1272
rect 126 1258 130 1262
rect 78 1248 82 1252
rect 86 1248 90 1252
rect 118 1248 122 1252
rect 70 1198 74 1202
rect 174 1288 178 1292
rect 190 1268 194 1272
rect 182 1258 186 1262
rect 174 1248 178 1252
rect 286 1348 290 1352
rect 326 1348 330 1352
rect 350 1348 354 1352
rect 398 1348 402 1352
rect 454 1348 458 1352
rect 222 1338 226 1342
rect 278 1338 282 1342
rect 334 1338 338 1342
rect 358 1338 362 1342
rect 382 1338 386 1342
rect 478 1338 482 1342
rect 510 1338 514 1342
rect 198 1238 202 1242
rect 86 1198 90 1202
rect 94 1198 98 1202
rect 126 1178 130 1182
rect 158 1198 162 1202
rect 142 1178 146 1182
rect 134 1158 138 1162
rect 6 1148 10 1152
rect 54 1148 58 1152
rect 78 1148 82 1152
rect 94 1148 98 1152
rect 62 1138 66 1142
rect 142 1148 146 1152
rect 150 1138 154 1142
rect 158 1138 162 1142
rect 110 1118 114 1122
rect 62 1048 66 1052
rect 46 1038 50 1042
rect 102 1058 106 1062
rect 110 1058 114 1062
rect 102 1038 106 1042
rect 70 1018 74 1022
rect 150 1098 154 1102
rect 254 1328 258 1332
rect 398 1328 402 1332
rect 262 1318 266 1322
rect 310 1318 314 1322
rect 222 1308 226 1312
rect 254 1308 258 1312
rect 350 1308 354 1312
rect 222 1298 226 1302
rect 222 1278 226 1282
rect 230 1278 234 1282
rect 310 1278 314 1282
rect 334 1278 338 1282
rect 382 1278 386 1282
rect 414 1278 418 1282
rect 222 1268 226 1272
rect 222 1258 226 1262
rect 214 1238 218 1242
rect 198 1158 202 1162
rect 238 1258 242 1262
rect 278 1258 282 1262
rect 318 1258 322 1262
rect 350 1258 354 1262
rect 550 1358 554 1362
rect 558 1298 562 1302
rect 446 1278 450 1282
rect 526 1278 530 1282
rect 534 1278 538 1282
rect 574 1278 578 1282
rect 614 1408 618 1412
rect 598 1348 602 1352
rect 654 1408 658 1412
rect 654 1358 658 1362
rect 622 1348 626 1352
rect 630 1348 634 1352
rect 646 1348 650 1352
rect 614 1338 618 1342
rect 614 1278 618 1282
rect 590 1268 594 1272
rect 614 1268 618 1272
rect 622 1268 626 1272
rect 254 1248 258 1252
rect 278 1248 282 1252
rect 302 1248 306 1252
rect 390 1248 394 1252
rect 526 1258 530 1262
rect 462 1248 466 1252
rect 478 1248 482 1252
rect 502 1248 506 1252
rect 518 1248 522 1252
rect 582 1248 586 1252
rect 446 1238 450 1242
rect 294 1228 298 1232
rect 422 1228 426 1232
rect 262 1198 266 1202
rect 382 1198 386 1202
rect 246 1158 250 1162
rect 190 1128 194 1132
rect 198 1088 202 1092
rect 190 1068 194 1072
rect 198 1068 202 1072
rect 166 1058 170 1062
rect 182 1058 186 1062
rect 270 1158 274 1162
rect 286 1158 290 1162
rect 350 1158 354 1162
rect 302 1148 306 1152
rect 238 1138 242 1142
rect 326 1138 330 1142
rect 302 1128 306 1132
rect 358 1128 362 1132
rect 238 1118 242 1122
rect 246 1068 250 1072
rect 286 1098 290 1102
rect 270 1058 274 1062
rect 318 1068 322 1072
rect 302 1058 306 1062
rect 350 1108 354 1112
rect 334 1078 338 1082
rect 150 1048 154 1052
rect 206 1048 210 1052
rect 238 1048 242 1052
rect 246 1048 250 1052
rect 262 1048 266 1052
rect 302 1048 306 1052
rect 326 1048 330 1052
rect 142 1038 146 1042
rect 134 1028 138 1032
rect 166 1028 170 1032
rect 150 1018 154 1022
rect 118 968 122 972
rect 126 968 130 972
rect 94 958 98 962
rect 126 958 130 962
rect 6 948 10 952
rect 6 878 10 882
rect 134 928 138 932
rect 222 988 226 992
rect 198 978 202 982
rect 174 958 178 962
rect 206 968 210 972
rect 262 1038 266 1042
rect 270 1028 274 1032
rect 294 1028 298 1032
rect 334 1018 338 1022
rect 286 1008 290 1012
rect 334 1008 338 1012
rect 286 998 290 1002
rect 270 988 274 992
rect 246 978 250 982
rect 254 978 258 982
rect 270 978 274 982
rect 262 968 266 972
rect 310 988 314 992
rect 302 978 306 982
rect 238 958 242 962
rect 326 968 330 972
rect 350 978 354 982
rect 342 968 346 972
rect 334 958 338 962
rect 174 948 178 952
rect 254 948 258 952
rect 318 948 322 952
rect 150 928 154 932
rect 126 908 130 912
rect 142 908 146 912
rect 166 928 170 932
rect 158 908 162 912
rect 166 888 170 892
rect 142 868 146 872
rect 6 828 10 832
rect 30 808 34 812
rect 46 778 50 782
rect 94 848 98 852
rect 142 848 146 852
rect 62 768 66 772
rect 54 758 58 762
rect 134 758 138 762
rect 14 748 18 752
rect 30 748 34 752
rect 62 748 66 752
rect 118 738 122 742
rect 174 778 178 782
rect 174 768 178 772
rect 158 728 162 732
rect 166 728 170 732
rect 142 708 146 712
rect 46 678 50 682
rect 102 678 106 682
rect 190 678 194 682
rect 54 668 58 672
rect 94 668 98 672
rect 126 668 130 672
rect 166 668 170 672
rect 38 648 42 652
rect 14 628 18 632
rect 30 548 34 552
rect 6 538 10 542
rect 70 658 74 662
rect 118 658 122 662
rect 86 648 90 652
rect 110 648 114 652
rect 166 648 170 652
rect 54 608 58 612
rect 78 588 82 592
rect 342 938 346 942
rect 406 1178 410 1182
rect 474 1203 478 1207
rect 481 1203 485 1207
rect 414 1158 418 1162
rect 414 1138 418 1142
rect 462 1138 466 1142
rect 470 1138 474 1142
rect 430 1128 434 1132
rect 422 1118 426 1122
rect 462 1118 466 1122
rect 382 1098 386 1102
rect 398 1078 402 1082
rect 430 1098 434 1102
rect 382 1068 386 1072
rect 422 1038 426 1042
rect 406 998 410 1002
rect 390 958 394 962
rect 366 938 370 942
rect 406 938 410 942
rect 358 918 362 922
rect 350 908 354 912
rect 278 878 282 882
rect 246 828 250 832
rect 222 768 226 772
rect 374 888 378 892
rect 390 918 394 922
rect 390 908 394 912
rect 494 1128 498 1132
rect 622 1248 626 1252
rect 606 1228 610 1232
rect 654 1228 658 1232
rect 590 1218 594 1222
rect 510 1158 514 1162
rect 534 1138 538 1142
rect 518 1128 522 1132
rect 550 1128 554 1132
rect 502 1078 506 1082
rect 494 1068 498 1072
rect 502 1068 506 1072
rect 438 1048 442 1052
rect 558 1078 562 1082
rect 630 1188 634 1192
rect 622 1168 626 1172
rect 582 1118 586 1122
rect 590 1118 594 1122
rect 654 1178 658 1182
rect 638 1148 642 1152
rect 662 1148 666 1152
rect 638 1128 642 1132
rect 630 1108 634 1112
rect 614 1098 618 1102
rect 590 1088 594 1092
rect 606 1088 610 1092
rect 630 1088 634 1092
rect 606 1068 610 1072
rect 518 1058 522 1062
rect 534 1058 538 1062
rect 550 1058 554 1062
rect 566 1058 570 1062
rect 598 1058 602 1062
rect 542 1048 546 1052
rect 574 1048 578 1052
rect 606 1048 610 1052
rect 622 1038 626 1042
rect 646 1098 650 1102
rect 718 1408 722 1412
rect 726 1398 730 1402
rect 718 1378 722 1382
rect 694 1368 698 1372
rect 678 1338 682 1342
rect 694 1338 698 1342
rect 678 1288 682 1292
rect 758 1398 762 1402
rect 742 1378 746 1382
rect 774 1378 778 1382
rect 798 1368 802 1372
rect 766 1358 770 1362
rect 814 1358 818 1362
rect 758 1348 762 1352
rect 790 1348 794 1352
rect 814 1348 818 1352
rect 838 1338 842 1342
rect 726 1328 730 1332
rect 774 1328 778 1332
rect 726 1318 730 1322
rect 702 1258 706 1262
rect 702 1248 706 1252
rect 766 1288 770 1292
rect 742 1258 746 1262
rect 710 1168 714 1172
rect 710 1158 714 1162
rect 678 1148 682 1152
rect 686 1138 690 1142
rect 718 1138 722 1142
rect 702 1118 706 1122
rect 670 1098 674 1102
rect 646 1048 650 1052
rect 654 1048 658 1052
rect 694 1068 698 1072
rect 518 1028 522 1032
rect 638 1028 642 1032
rect 474 1003 478 1007
rect 481 1003 485 1007
rect 446 998 450 1002
rect 526 1008 530 1012
rect 558 998 562 1002
rect 446 988 450 992
rect 574 988 578 992
rect 598 988 602 992
rect 494 978 498 982
rect 574 978 578 982
rect 590 978 594 982
rect 430 958 434 962
rect 446 948 450 952
rect 462 948 466 952
rect 502 958 506 962
rect 526 948 530 952
rect 446 938 450 942
rect 454 938 458 942
rect 510 938 514 942
rect 430 878 434 882
rect 310 868 314 872
rect 318 868 322 872
rect 334 868 338 872
rect 358 868 362 872
rect 374 868 378 872
rect 294 858 298 862
rect 350 848 354 852
rect 358 848 362 852
rect 398 868 402 872
rect 422 868 426 872
rect 430 858 434 862
rect 406 848 410 852
rect 278 838 282 842
rect 302 838 306 842
rect 350 838 354 842
rect 390 838 394 842
rect 430 828 434 832
rect 502 898 506 902
rect 542 958 546 962
rect 630 988 634 992
rect 614 968 618 972
rect 622 968 626 972
rect 638 968 642 972
rect 630 958 634 962
rect 606 948 610 952
rect 566 938 570 942
rect 598 938 602 942
rect 534 928 538 932
rect 590 928 594 932
rect 534 918 538 922
rect 566 908 570 912
rect 534 898 538 902
rect 526 878 530 882
rect 518 868 522 872
rect 550 868 554 872
rect 462 818 466 822
rect 474 803 478 807
rect 481 803 485 807
rect 454 788 458 792
rect 438 778 442 782
rect 398 768 402 772
rect 262 758 266 762
rect 382 758 386 762
rect 230 748 234 752
rect 222 718 226 722
rect 422 748 426 752
rect 430 748 434 752
rect 246 738 250 742
rect 366 738 370 742
rect 318 728 322 732
rect 406 728 410 732
rect 334 698 338 702
rect 654 958 658 962
rect 662 958 666 962
rect 654 938 658 942
rect 598 868 602 872
rect 630 908 634 912
rect 622 878 626 882
rect 678 1008 682 1012
rect 710 978 714 982
rect 742 1158 746 1162
rect 750 1158 754 1162
rect 750 1138 754 1142
rect 742 1078 746 1082
rect 782 1318 786 1322
rect 806 1298 810 1302
rect 822 1298 826 1302
rect 830 1298 834 1302
rect 878 1408 882 1412
rect 878 1348 882 1352
rect 902 1348 906 1352
rect 910 1338 914 1342
rect 886 1328 890 1332
rect 846 1308 850 1312
rect 854 1308 858 1312
rect 814 1268 818 1272
rect 806 1248 810 1252
rect 830 1258 834 1262
rect 838 1258 842 1262
rect 838 1238 842 1242
rect 814 1218 818 1222
rect 830 1218 834 1222
rect 806 1158 810 1162
rect 830 1168 834 1172
rect 862 1298 866 1302
rect 854 1238 858 1242
rect 894 1308 898 1312
rect 878 1248 882 1252
rect 894 1248 898 1252
rect 902 1238 906 1242
rect 886 1228 890 1232
rect 918 1248 922 1252
rect 918 1228 922 1232
rect 910 1218 914 1222
rect 870 1188 874 1192
rect 886 1168 890 1172
rect 910 1168 914 1172
rect 1334 1398 1338 1402
rect 998 1388 1002 1392
rect 1062 1388 1066 1392
rect 1294 1368 1298 1372
rect 1046 1358 1050 1362
rect 1118 1358 1122 1362
rect 1166 1358 1170 1362
rect 1174 1358 1178 1362
rect 1190 1358 1194 1362
rect 1214 1358 1218 1362
rect 1230 1358 1234 1362
rect 1310 1358 1314 1362
rect 950 1348 954 1352
rect 1014 1348 1018 1352
rect 1070 1348 1074 1352
rect 1110 1348 1114 1352
rect 1126 1348 1130 1352
rect 1262 1348 1266 1352
rect 974 1338 978 1342
rect 1030 1338 1034 1342
rect 942 1328 946 1332
rect 1022 1318 1026 1322
rect 966 1308 970 1312
rect 986 1303 990 1307
rect 993 1303 997 1307
rect 1046 1328 1050 1332
rect 1086 1328 1090 1332
rect 1166 1328 1170 1332
rect 1190 1338 1194 1342
rect 1294 1338 1298 1342
rect 1318 1338 1322 1342
rect 1054 1318 1058 1322
rect 1062 1318 1066 1322
rect 1094 1318 1098 1322
rect 1134 1318 1138 1322
rect 1158 1318 1162 1322
rect 1174 1318 1178 1322
rect 1206 1318 1210 1322
rect 1358 1378 1362 1382
rect 1358 1348 1362 1352
rect 1350 1338 1354 1342
rect 1262 1318 1266 1322
rect 1230 1288 1234 1292
rect 950 1278 954 1282
rect 958 1278 962 1282
rect 1014 1278 1018 1282
rect 1038 1278 1042 1282
rect 1222 1278 1226 1282
rect 1102 1268 1106 1272
rect 1118 1268 1122 1272
rect 1198 1268 1202 1272
rect 1070 1258 1074 1262
rect 1086 1258 1090 1262
rect 1182 1258 1186 1262
rect 1198 1258 1202 1262
rect 1142 1248 1146 1252
rect 1158 1248 1162 1252
rect 1038 1238 1042 1242
rect 1054 1238 1058 1242
rect 1126 1238 1130 1242
rect 1142 1228 1146 1232
rect 974 1218 978 1222
rect 926 1208 930 1212
rect 926 1198 930 1202
rect 950 1208 954 1212
rect 878 1158 882 1162
rect 894 1158 898 1162
rect 798 1138 802 1142
rect 822 1138 826 1142
rect 854 1138 858 1142
rect 766 1118 770 1122
rect 862 1118 866 1122
rect 734 1038 738 1042
rect 854 1078 858 1082
rect 790 1058 794 1062
rect 830 1068 834 1072
rect 838 1058 842 1062
rect 854 1048 858 1052
rect 806 1028 810 1032
rect 838 1018 842 1022
rect 726 978 730 982
rect 710 958 714 962
rect 702 888 706 892
rect 710 878 714 882
rect 686 868 690 872
rect 582 858 586 862
rect 598 858 602 862
rect 614 858 618 862
rect 646 858 650 862
rect 558 848 562 852
rect 574 848 578 852
rect 694 858 698 862
rect 526 838 530 842
rect 566 838 570 842
rect 638 838 642 842
rect 662 838 666 842
rect 686 838 690 842
rect 526 788 530 792
rect 590 798 594 802
rect 614 798 618 802
rect 630 798 634 802
rect 638 798 642 802
rect 550 748 554 752
rect 622 768 626 772
rect 670 798 674 802
rect 694 798 698 802
rect 910 1138 914 1142
rect 942 1168 946 1172
rect 1142 1198 1146 1202
rect 1142 1178 1146 1182
rect 1118 1168 1122 1172
rect 982 1158 986 1162
rect 998 1158 1002 1162
rect 1022 1158 1026 1162
rect 1102 1158 1106 1162
rect 1134 1158 1138 1162
rect 926 1138 930 1142
rect 886 1058 890 1062
rect 902 1068 906 1072
rect 918 1078 922 1082
rect 870 1048 874 1052
rect 894 1048 898 1052
rect 918 1048 922 1052
rect 878 1038 882 1042
rect 886 1038 890 1042
rect 942 1068 946 1072
rect 1134 1148 1138 1152
rect 1094 1138 1098 1142
rect 1014 1128 1018 1132
rect 986 1103 990 1107
rect 993 1103 997 1107
rect 1006 1098 1010 1102
rect 974 1088 978 1092
rect 966 1078 970 1082
rect 926 1028 930 1032
rect 934 1028 938 1032
rect 846 998 850 1002
rect 862 998 866 1002
rect 742 958 746 962
rect 774 958 778 962
rect 734 948 738 952
rect 726 928 730 932
rect 734 878 738 882
rect 758 868 762 872
rect 742 858 746 862
rect 782 948 786 952
rect 806 968 810 972
rect 830 968 834 972
rect 798 958 802 962
rect 798 928 802 932
rect 790 898 794 902
rect 822 938 826 942
rect 838 948 842 952
rect 854 988 858 992
rect 862 988 866 992
rect 934 1008 938 1012
rect 910 978 914 982
rect 926 978 930 982
rect 1014 1078 1018 1082
rect 1014 1058 1018 1062
rect 966 988 970 992
rect 854 958 858 962
rect 902 958 906 962
rect 934 958 938 962
rect 950 958 954 962
rect 982 958 986 962
rect 814 928 818 932
rect 838 928 842 932
rect 846 928 850 932
rect 822 898 826 902
rect 886 948 890 952
rect 926 948 930 952
rect 958 938 962 942
rect 846 908 850 912
rect 870 908 874 912
rect 838 878 842 882
rect 774 868 778 872
rect 798 868 802 872
rect 862 868 866 872
rect 950 908 954 912
rect 926 878 930 882
rect 878 868 882 872
rect 846 858 850 862
rect 870 858 874 862
rect 878 858 882 862
rect 718 848 722 852
rect 838 838 842 842
rect 734 778 738 782
rect 710 768 714 772
rect 718 768 722 772
rect 790 808 794 812
rect 814 798 818 802
rect 742 768 746 772
rect 790 768 794 772
rect 806 768 810 772
rect 534 738 538 742
rect 574 738 578 742
rect 582 738 586 742
rect 630 738 634 742
rect 510 728 514 732
rect 462 718 466 722
rect 446 698 450 702
rect 334 688 338 692
rect 230 668 234 672
rect 246 668 250 672
rect 214 648 218 652
rect 262 648 266 652
rect 286 648 290 652
rect 150 578 154 582
rect 166 578 170 582
rect 110 568 114 572
rect 142 568 146 572
rect 158 568 162 572
rect 174 568 178 572
rect 70 558 74 562
rect 86 558 90 562
rect 302 638 306 642
rect 318 628 322 632
rect 438 668 442 672
rect 358 648 362 652
rect 366 638 370 642
rect 350 628 354 632
rect 278 618 282 622
rect 294 618 298 622
rect 318 618 322 622
rect 326 618 330 622
rect 270 598 274 602
rect 294 598 298 602
rect 342 598 346 602
rect 270 568 274 572
rect 318 568 322 572
rect 126 558 130 562
rect 134 558 138 562
rect 238 558 242 562
rect 334 558 338 562
rect 350 558 354 562
rect 86 548 90 552
rect 102 548 106 552
rect 126 548 130 552
rect 62 538 66 542
rect 86 538 90 542
rect 46 518 50 522
rect 6 488 10 492
rect 94 478 98 482
rect 126 478 130 482
rect 6 468 10 472
rect 30 468 34 472
rect 54 468 58 472
rect 118 468 122 472
rect 38 458 42 462
rect 6 428 10 432
rect 78 458 82 462
rect 158 538 162 542
rect 150 528 154 532
rect 222 548 226 552
rect 174 538 178 542
rect 182 538 186 542
rect 206 538 210 542
rect 270 538 274 542
rect 294 538 298 542
rect 166 498 170 502
rect 166 468 170 472
rect 70 448 74 452
rect 118 448 122 452
rect 70 418 74 422
rect 46 398 50 402
rect 54 398 58 402
rect 70 398 74 402
rect 142 438 146 442
rect 118 388 122 392
rect 134 388 138 392
rect 118 378 122 382
rect 198 498 202 502
rect 182 428 186 432
rect 238 528 242 532
rect 278 528 282 532
rect 286 498 290 502
rect 310 508 314 512
rect 294 488 298 492
rect 262 468 266 472
rect 214 458 218 462
rect 230 458 234 462
rect 246 458 250 462
rect 190 408 194 412
rect 166 388 170 392
rect 126 368 130 372
rect 94 358 98 362
rect 102 358 106 362
rect 134 358 138 362
rect 14 348 18 352
rect 22 348 26 352
rect 46 348 50 352
rect 70 348 74 352
rect 94 348 98 352
rect 6 288 10 292
rect 6 158 10 162
rect 78 338 82 342
rect 22 328 26 332
rect 78 318 82 322
rect 54 298 58 302
rect 22 278 26 282
rect 38 278 42 282
rect 54 268 58 272
rect 102 268 106 272
rect 86 258 90 262
rect 70 248 74 252
rect 150 368 154 372
rect 190 368 194 372
rect 214 448 218 452
rect 206 438 210 442
rect 206 388 210 392
rect 190 358 194 362
rect 238 438 242 442
rect 254 438 258 442
rect 342 548 346 552
rect 462 668 466 672
rect 398 648 402 652
rect 462 648 466 652
rect 462 638 466 642
rect 390 628 394 632
rect 390 618 394 622
rect 422 628 426 632
rect 414 618 418 622
rect 414 598 418 602
rect 406 568 410 572
rect 454 588 458 592
rect 390 558 394 562
rect 366 528 370 532
rect 334 488 338 492
rect 366 488 370 492
rect 382 498 386 502
rect 422 538 426 542
rect 406 528 410 532
rect 838 778 842 782
rect 822 768 826 772
rect 894 848 898 852
rect 862 838 866 842
rect 942 848 946 852
rect 926 818 930 822
rect 886 808 890 812
rect 942 808 946 812
rect 854 798 858 802
rect 870 798 874 802
rect 934 788 938 792
rect 902 778 906 782
rect 934 778 938 782
rect 886 768 890 772
rect 870 758 874 762
rect 870 748 874 752
rect 686 738 690 742
rect 758 738 762 742
rect 774 738 778 742
rect 806 738 810 742
rect 830 738 834 742
rect 862 738 866 742
rect 558 728 562 732
rect 614 728 618 732
rect 646 728 650 732
rect 678 728 682 732
rect 550 708 554 712
rect 622 698 626 702
rect 534 678 538 682
rect 614 678 618 682
rect 518 668 522 672
rect 558 668 562 672
rect 550 658 554 662
rect 470 628 474 632
rect 518 628 522 632
rect 526 618 530 622
rect 474 603 478 607
rect 481 603 485 607
rect 558 628 562 632
rect 550 608 554 612
rect 598 648 602 652
rect 590 638 594 642
rect 582 618 586 622
rect 526 598 530 602
rect 534 588 538 592
rect 494 578 498 582
rect 550 578 554 582
rect 502 568 506 572
rect 518 568 522 572
rect 502 558 506 562
rect 462 538 466 542
rect 502 508 506 512
rect 462 488 466 492
rect 494 488 498 492
rect 342 478 346 482
rect 374 478 378 482
rect 398 478 402 482
rect 454 478 458 482
rect 382 468 386 472
rect 414 468 418 472
rect 438 468 442 472
rect 374 458 378 462
rect 366 448 370 452
rect 294 438 298 442
rect 374 428 378 432
rect 318 418 322 422
rect 278 408 282 412
rect 294 408 298 412
rect 246 388 250 392
rect 222 368 226 372
rect 158 338 162 342
rect 254 368 258 372
rect 262 358 266 362
rect 246 348 250 352
rect 214 338 218 342
rect 158 278 162 282
rect 414 388 418 392
rect 446 438 450 442
rect 502 478 506 482
rect 510 478 514 482
rect 470 468 474 472
rect 474 403 478 407
rect 481 403 485 407
rect 566 538 570 542
rect 574 508 578 512
rect 606 628 610 632
rect 606 598 610 602
rect 550 468 554 472
rect 534 458 538 462
rect 518 438 522 442
rect 542 438 546 442
rect 518 428 522 432
rect 582 468 586 472
rect 566 458 570 462
rect 574 438 578 442
rect 558 408 562 412
rect 550 398 554 402
rect 510 388 514 392
rect 390 378 394 382
rect 422 378 426 382
rect 590 378 594 382
rect 318 368 322 372
rect 374 368 378 372
rect 398 368 402 372
rect 350 358 354 362
rect 374 358 378 362
rect 310 348 314 352
rect 246 338 250 342
rect 286 338 290 342
rect 278 328 282 332
rect 318 328 322 332
rect 374 328 378 332
rect 270 278 274 282
rect 230 268 234 272
rect 262 268 266 272
rect 270 268 274 272
rect 206 258 210 262
rect 238 258 242 262
rect 38 238 42 242
rect 78 238 82 242
rect 94 238 98 242
rect 126 238 130 242
rect 142 238 146 242
rect 38 228 42 232
rect 78 218 82 222
rect 118 218 122 222
rect 62 208 66 212
rect 38 178 42 182
rect 22 168 26 172
rect 14 148 18 152
rect 54 128 58 132
rect 6 88 10 92
rect 142 218 146 222
rect 86 188 90 192
rect 118 188 122 192
rect 70 158 74 162
rect 86 148 90 152
rect 78 138 82 142
rect 86 118 90 122
rect 46 78 50 82
rect 110 98 114 102
rect 94 78 98 82
rect 134 168 138 172
rect 166 218 170 222
rect 294 258 298 262
rect 214 248 218 252
rect 198 238 202 242
rect 230 238 234 242
rect 150 208 154 212
rect 166 208 170 212
rect 182 208 186 212
rect 182 158 186 162
rect 198 148 202 152
rect 158 128 162 132
rect 206 118 210 122
rect 158 108 162 112
rect 150 88 154 92
rect 166 98 170 102
rect 206 98 210 102
rect 174 88 178 92
rect 118 68 122 72
rect 254 218 258 222
rect 230 188 234 192
rect 238 178 242 182
rect 230 128 234 132
rect 350 308 354 312
rect 318 278 322 282
rect 342 278 346 282
rect 366 278 370 282
rect 374 278 378 282
rect 390 278 394 282
rect 326 268 330 272
rect 366 268 370 272
rect 286 238 290 242
rect 302 238 306 242
rect 310 238 314 242
rect 318 218 322 222
rect 334 178 338 182
rect 262 158 266 162
rect 270 158 274 162
rect 262 148 266 152
rect 294 138 298 142
rect 262 98 266 102
rect 294 98 298 102
rect 246 88 250 92
rect 246 78 250 82
rect 358 158 362 162
rect 326 148 330 152
rect 318 98 322 102
rect 398 268 402 272
rect 406 268 410 272
rect 454 368 458 372
rect 486 368 490 372
rect 550 368 554 372
rect 438 358 442 362
rect 454 338 458 342
rect 430 328 434 332
rect 470 328 474 332
rect 446 298 450 302
rect 454 278 458 282
rect 462 278 466 282
rect 422 258 426 262
rect 446 258 450 262
rect 438 248 442 252
rect 510 358 514 362
rect 518 358 522 362
rect 582 358 586 362
rect 574 348 578 352
rect 718 728 722 732
rect 726 728 730 732
rect 702 698 706 702
rect 726 698 730 702
rect 678 678 682 682
rect 806 728 810 732
rect 750 708 754 712
rect 758 688 762 692
rect 830 708 834 712
rect 766 678 770 682
rect 782 678 786 682
rect 686 668 690 672
rect 734 668 738 672
rect 766 668 770 672
rect 806 668 810 672
rect 846 668 850 672
rect 630 658 634 662
rect 670 658 674 662
rect 686 658 690 662
rect 702 658 706 662
rect 638 648 642 652
rect 654 648 658 652
rect 654 638 658 642
rect 662 638 666 642
rect 678 638 682 642
rect 630 618 634 622
rect 622 598 626 602
rect 670 628 674 632
rect 654 578 658 582
rect 630 538 634 542
rect 678 568 682 572
rect 718 568 722 572
rect 702 548 706 552
rect 646 538 650 542
rect 630 508 634 512
rect 638 508 642 512
rect 702 508 706 512
rect 614 488 618 492
rect 678 488 682 492
rect 758 538 762 542
rect 766 538 770 542
rect 750 518 754 522
rect 662 478 666 482
rect 694 478 698 482
rect 710 478 714 482
rect 742 478 746 482
rect 622 458 626 462
rect 662 458 666 462
rect 726 458 730 462
rect 734 458 738 462
rect 606 358 610 362
rect 614 358 618 362
rect 510 328 514 332
rect 542 328 546 332
rect 566 328 570 332
rect 494 318 498 322
rect 510 298 514 302
rect 574 318 578 322
rect 510 288 514 292
rect 526 288 530 292
rect 582 288 586 292
rect 518 278 522 282
rect 534 278 538 282
rect 598 328 602 332
rect 646 448 650 452
rect 654 448 658 452
rect 654 368 658 372
rect 622 278 626 282
rect 470 268 474 272
rect 494 268 498 272
rect 566 268 570 272
rect 590 268 594 272
rect 614 268 618 272
rect 474 203 478 207
rect 481 203 485 207
rect 406 178 410 182
rect 390 108 394 112
rect 342 88 346 92
rect 334 78 338 82
rect 358 78 362 82
rect 278 68 282 72
rect 318 68 322 72
rect 38 58 42 62
rect 78 58 82 62
rect 198 58 202 62
rect 78 48 82 52
rect 102 48 106 52
rect 150 48 154 52
rect 238 48 242 52
rect 254 48 258 52
rect 278 48 282 52
rect 302 48 306 52
rect 118 38 122 42
rect 318 28 322 32
rect 374 68 378 72
rect 390 68 394 72
rect 502 248 506 252
rect 550 238 554 242
rect 670 358 674 362
rect 726 418 730 422
rect 694 348 698 352
rect 710 338 714 342
rect 726 338 730 342
rect 654 328 658 332
rect 686 328 690 332
rect 742 328 746 332
rect 662 318 666 322
rect 678 318 682 322
rect 678 308 682 312
rect 646 288 650 292
rect 638 278 642 282
rect 710 318 714 322
rect 918 758 922 762
rect 910 748 914 752
rect 986 903 990 907
rect 993 903 997 907
rect 982 878 986 882
rect 998 878 1002 882
rect 1038 1108 1042 1112
rect 1054 1118 1058 1122
rect 1046 1078 1050 1082
rect 1070 1068 1074 1072
rect 1046 1048 1050 1052
rect 1038 1018 1042 1022
rect 1046 998 1050 1002
rect 1062 988 1066 992
rect 1038 958 1042 962
rect 1054 958 1058 962
rect 1022 948 1026 952
rect 1054 948 1058 952
rect 1046 848 1050 852
rect 982 828 986 832
rect 1014 828 1018 832
rect 950 788 954 792
rect 1046 818 1050 822
rect 1030 798 1034 802
rect 1022 788 1026 792
rect 998 768 1002 772
rect 958 758 962 762
rect 1014 748 1018 752
rect 958 738 962 742
rect 1030 738 1034 742
rect 966 728 970 732
rect 910 718 914 722
rect 894 698 898 702
rect 902 688 906 692
rect 886 668 890 672
rect 814 658 818 662
rect 854 658 858 662
rect 862 658 866 662
rect 870 658 874 662
rect 798 648 802 652
rect 918 678 922 682
rect 926 678 930 682
rect 966 708 970 712
rect 950 698 954 702
rect 986 703 990 707
rect 993 703 997 707
rect 1102 1108 1106 1112
rect 1086 1088 1090 1092
rect 1086 1078 1090 1082
rect 1158 1168 1162 1172
rect 1142 1088 1146 1092
rect 1190 1248 1194 1252
rect 1230 1268 1234 1272
rect 1246 1258 1250 1262
rect 1246 1238 1250 1242
rect 1278 1238 1282 1242
rect 1326 1288 1330 1292
rect 1318 1278 1322 1282
rect 1318 1268 1322 1272
rect 1318 1248 1322 1252
rect 1254 1228 1258 1232
rect 1286 1228 1290 1232
rect 1206 1158 1210 1162
rect 1182 1128 1186 1132
rect 1198 1118 1202 1122
rect 1174 1108 1178 1112
rect 1190 1078 1194 1082
rect 1222 1098 1226 1102
rect 1222 1078 1226 1082
rect 1118 1068 1122 1072
rect 1174 1068 1178 1072
rect 1102 1058 1106 1062
rect 1198 1058 1202 1062
rect 1070 978 1074 982
rect 1070 868 1074 872
rect 1070 848 1074 852
rect 1110 1038 1114 1042
rect 1150 1038 1154 1042
rect 1094 998 1098 1002
rect 1142 998 1146 1002
rect 1134 948 1138 952
rect 1094 918 1098 922
rect 1102 918 1106 922
rect 1102 878 1106 882
rect 1110 868 1114 872
rect 1070 838 1074 842
rect 1054 808 1058 812
rect 1102 858 1106 862
rect 1134 908 1138 912
rect 1238 1188 1242 1192
rect 1254 1168 1258 1172
rect 1254 1158 1258 1162
rect 1246 1078 1250 1082
rect 1286 1178 1290 1182
rect 1302 1178 1306 1182
rect 1278 1158 1282 1162
rect 1342 1268 1346 1272
rect 1342 1238 1346 1242
rect 1318 1228 1322 1232
rect 1326 1168 1330 1172
rect 1294 1158 1298 1162
rect 1334 1158 1338 1162
rect 1286 1138 1290 1142
rect 1310 1138 1314 1142
rect 1374 1358 1378 1362
rect 1398 1358 1402 1362
rect 1430 1358 1434 1362
rect 1382 1348 1386 1352
rect 1430 1338 1434 1342
rect 1390 1318 1394 1322
rect 1454 1318 1458 1322
rect 1374 1278 1378 1282
rect 1438 1288 1442 1292
rect 1430 1278 1434 1282
rect 1390 1268 1394 1272
rect 1414 1268 1418 1272
rect 1374 1238 1378 1242
rect 1422 1258 1426 1262
rect 1422 1248 1426 1252
rect 1382 1228 1386 1232
rect 1414 1228 1418 1232
rect 1406 1218 1410 1222
rect 1358 1198 1362 1202
rect 1358 1168 1362 1172
rect 1270 1068 1274 1072
rect 1302 1068 1306 1072
rect 1270 1058 1274 1062
rect 1294 1058 1298 1062
rect 1262 1048 1266 1052
rect 1326 1088 1330 1092
rect 1342 1108 1346 1112
rect 1358 1138 1362 1142
rect 1446 1218 1450 1222
rect 1438 1168 1442 1172
rect 1382 1158 1386 1162
rect 1398 1158 1402 1162
rect 1398 1148 1402 1152
rect 1390 1138 1394 1142
rect 1406 1138 1410 1142
rect 1366 1128 1370 1132
rect 1350 1078 1354 1082
rect 1374 1078 1378 1082
rect 1382 1078 1386 1082
rect 1398 1078 1402 1082
rect 1342 1068 1346 1072
rect 1366 1068 1370 1072
rect 1334 1058 1338 1062
rect 1318 1048 1322 1052
rect 1278 1038 1282 1042
rect 1222 1018 1226 1022
rect 1206 1008 1210 1012
rect 1150 968 1154 972
rect 1174 968 1178 972
rect 1182 968 1186 972
rect 1254 1008 1258 1012
rect 1246 958 1250 962
rect 1206 948 1210 952
rect 1238 948 1242 952
rect 1262 948 1266 952
rect 1222 938 1226 942
rect 1174 928 1178 932
rect 1214 928 1218 932
rect 1286 928 1290 932
rect 1302 968 1306 972
rect 1206 908 1210 912
rect 1142 898 1146 902
rect 1254 918 1258 922
rect 1238 898 1242 902
rect 1270 898 1274 902
rect 1238 888 1242 892
rect 1254 888 1258 892
rect 1294 878 1298 882
rect 1326 968 1330 972
rect 1398 1068 1402 1072
rect 1350 1048 1354 1052
rect 1358 1018 1362 1022
rect 1438 1138 1442 1142
rect 1446 1138 1450 1142
rect 1462 1138 1466 1142
rect 1470 1138 1474 1142
rect 1446 1128 1450 1132
rect 1470 1088 1474 1092
rect 1414 1058 1418 1062
rect 1438 1058 1442 1062
rect 1422 1048 1426 1052
rect 1446 1048 1450 1052
rect 1398 1028 1402 1032
rect 1342 988 1346 992
rect 1374 988 1378 992
rect 1406 988 1410 992
rect 1366 968 1370 972
rect 1326 958 1330 962
rect 1374 958 1378 962
rect 1318 928 1322 932
rect 1318 908 1322 912
rect 1182 868 1186 872
rect 1190 868 1194 872
rect 1214 868 1218 872
rect 1294 868 1298 872
rect 1302 868 1306 872
rect 1310 868 1314 872
rect 1166 858 1170 862
rect 1142 848 1146 852
rect 1174 838 1178 842
rect 1118 828 1122 832
rect 1342 948 1346 952
rect 1358 948 1362 952
rect 1398 938 1402 942
rect 1358 928 1362 932
rect 1390 928 1394 932
rect 1350 858 1354 862
rect 1326 848 1330 852
rect 1334 848 1338 852
rect 1406 918 1410 922
rect 1366 908 1370 912
rect 1398 878 1402 882
rect 1374 848 1378 852
rect 1390 848 1394 852
rect 1214 838 1218 842
rect 1286 838 1290 842
rect 1294 838 1298 842
rect 1310 838 1314 842
rect 1326 838 1330 842
rect 1342 838 1346 842
rect 1198 808 1202 812
rect 1270 798 1274 802
rect 1310 798 1314 802
rect 1326 798 1330 802
rect 1158 788 1162 792
rect 1294 788 1298 792
rect 1094 768 1098 772
rect 1158 768 1162 772
rect 1254 768 1258 772
rect 1294 768 1298 772
rect 1086 758 1090 762
rect 1118 758 1122 762
rect 1214 758 1218 762
rect 1318 788 1322 792
rect 1438 1038 1442 1042
rect 1454 1038 1458 1042
rect 1430 1018 1434 1022
rect 1470 998 1474 1002
rect 1430 968 1434 972
rect 1478 968 1482 972
rect 1438 958 1442 962
rect 1446 938 1450 942
rect 1454 938 1458 942
rect 1478 928 1482 932
rect 1422 878 1426 882
rect 1406 848 1410 852
rect 1318 768 1322 772
rect 1358 768 1362 772
rect 1334 758 1338 762
rect 1038 688 1042 692
rect 1310 738 1314 742
rect 1358 738 1362 742
rect 1182 718 1186 722
rect 1206 708 1210 712
rect 1230 698 1234 702
rect 1054 678 1058 682
rect 1118 678 1122 682
rect 894 638 898 642
rect 1118 668 1122 672
rect 1254 668 1258 672
rect 1254 658 1258 662
rect 1270 658 1274 662
rect 1022 648 1026 652
rect 1302 688 1306 692
rect 1294 678 1298 682
rect 1318 678 1322 682
rect 1294 668 1298 672
rect 1286 658 1290 662
rect 1278 648 1282 652
rect 1094 638 1098 642
rect 1214 638 1218 642
rect 870 628 874 632
rect 990 628 994 632
rect 846 618 850 622
rect 838 558 842 562
rect 790 548 794 552
rect 1014 608 1018 612
rect 934 568 938 572
rect 918 558 922 562
rect 942 558 946 562
rect 998 558 1002 562
rect 1310 648 1314 652
rect 1102 568 1106 572
rect 1110 568 1114 572
rect 1150 568 1154 572
rect 1214 568 1218 572
rect 1222 568 1226 572
rect 1238 568 1242 572
rect 1254 568 1258 572
rect 1118 558 1122 562
rect 1166 558 1170 562
rect 1262 558 1266 562
rect 1070 548 1074 552
rect 1150 548 1154 552
rect 798 538 802 542
rect 918 538 922 542
rect 950 538 954 542
rect 958 538 962 542
rect 998 538 1002 542
rect 1022 538 1026 542
rect 1046 538 1050 542
rect 774 498 778 502
rect 758 478 762 482
rect 942 518 946 522
rect 806 508 810 512
rect 830 508 834 512
rect 806 498 810 502
rect 790 468 794 472
rect 822 468 826 472
rect 846 468 850 472
rect 870 458 874 462
rect 886 458 890 462
rect 790 448 794 452
rect 758 438 762 442
rect 806 438 810 442
rect 750 308 754 312
rect 790 408 794 412
rect 814 408 818 412
rect 790 358 794 362
rect 806 358 810 362
rect 838 428 842 432
rect 838 398 842 402
rect 838 358 842 362
rect 774 348 778 352
rect 790 348 794 352
rect 806 348 810 352
rect 766 328 770 332
rect 654 268 658 272
rect 686 268 690 272
rect 630 258 634 262
rect 646 248 650 252
rect 702 248 706 252
rect 662 228 666 232
rect 694 228 698 232
rect 702 228 706 232
rect 622 218 626 222
rect 686 188 690 192
rect 702 188 706 192
rect 662 178 666 182
rect 630 158 634 162
rect 414 148 418 152
rect 486 148 490 152
rect 518 148 522 152
rect 446 138 450 142
rect 462 128 466 132
rect 422 118 426 122
rect 558 138 562 142
rect 534 128 538 132
rect 518 98 522 102
rect 462 78 466 82
rect 526 88 530 92
rect 598 118 602 122
rect 574 108 578 112
rect 550 98 554 102
rect 438 68 442 72
rect 462 68 466 72
rect 542 68 546 72
rect 574 88 578 92
rect 558 78 562 82
rect 574 78 578 82
rect 398 58 402 62
rect 422 48 426 52
rect 342 38 346 42
rect 334 18 338 22
rect 510 48 514 52
rect 494 28 498 32
rect 550 28 554 32
rect 438 8 442 12
rect 454 8 458 12
rect 474 3 478 7
rect 481 3 485 7
rect 622 148 626 152
rect 622 108 626 112
rect 622 78 626 82
rect 566 48 570 52
rect 598 48 602 52
rect 622 38 626 42
rect 742 258 746 262
rect 734 248 738 252
rect 726 198 730 202
rect 718 178 722 182
rect 822 338 826 342
rect 774 278 778 282
rect 766 268 770 272
rect 710 158 714 162
rect 710 138 714 142
rect 646 128 650 132
rect 646 118 650 122
rect 710 128 714 132
rect 686 108 690 112
rect 670 88 674 92
rect 662 78 666 82
rect 694 78 698 82
rect 662 48 666 52
rect 710 48 714 52
rect 718 38 722 42
rect 734 128 738 132
rect 758 138 762 142
rect 798 248 802 252
rect 782 228 786 232
rect 790 228 794 232
rect 806 228 810 232
rect 814 208 818 212
rect 862 438 866 442
rect 974 528 978 532
rect 1046 528 1050 532
rect 1070 528 1074 532
rect 942 478 946 482
rect 926 468 930 472
rect 878 438 882 442
rect 894 438 898 442
rect 918 438 922 442
rect 878 408 882 412
rect 870 358 874 362
rect 862 338 866 342
rect 986 503 990 507
rect 993 503 997 507
rect 990 488 994 492
rect 1022 468 1026 472
rect 1038 468 1042 472
rect 1102 518 1106 522
rect 1142 528 1146 532
rect 1078 488 1082 492
rect 1110 488 1114 492
rect 1118 488 1122 492
rect 1086 478 1090 482
rect 1110 478 1114 482
rect 1134 478 1138 482
rect 1158 478 1162 482
rect 1118 468 1122 472
rect 1134 468 1138 472
rect 982 458 986 462
rect 1030 458 1034 462
rect 1046 458 1050 462
rect 1070 458 1074 462
rect 966 448 970 452
rect 1038 448 1042 452
rect 966 428 970 432
rect 950 408 954 412
rect 974 408 978 412
rect 918 398 922 402
rect 886 378 890 382
rect 910 368 914 372
rect 1022 418 1026 422
rect 1062 448 1066 452
rect 1078 448 1082 452
rect 1046 408 1050 412
rect 1038 368 1042 372
rect 1078 368 1082 372
rect 926 358 930 362
rect 950 358 954 362
rect 1022 358 1026 362
rect 1046 358 1050 362
rect 918 348 922 352
rect 902 338 906 342
rect 838 308 842 312
rect 846 308 850 312
rect 870 308 874 312
rect 926 288 930 292
rect 902 268 906 272
rect 910 268 914 272
rect 822 198 826 202
rect 862 248 866 252
rect 838 228 842 232
rect 846 198 850 202
rect 838 188 842 192
rect 774 178 778 182
rect 814 178 818 182
rect 830 178 834 182
rect 774 148 778 152
rect 790 138 794 142
rect 774 128 778 132
rect 782 88 786 92
rect 742 78 746 82
rect 758 78 762 82
rect 734 48 738 52
rect 766 28 770 32
rect 726 8 730 12
rect 750 8 754 12
rect 806 128 810 132
rect 806 108 810 112
rect 798 58 802 62
rect 790 38 794 42
rect 878 248 882 252
rect 862 228 866 232
rect 870 228 874 232
rect 950 338 954 342
rect 990 328 994 332
rect 942 308 946 312
rect 986 303 990 307
rect 993 303 997 307
rect 942 268 946 272
rect 966 268 970 272
rect 990 268 994 272
rect 934 248 938 252
rect 950 248 954 252
rect 974 248 978 252
rect 982 248 986 252
rect 902 228 906 232
rect 886 208 890 212
rect 894 208 898 212
rect 878 198 882 202
rect 838 158 842 162
rect 830 138 834 142
rect 846 138 850 142
rect 830 128 834 132
rect 822 108 826 112
rect 958 238 962 242
rect 894 188 898 192
rect 910 188 914 192
rect 934 188 938 192
rect 902 168 906 172
rect 974 228 978 232
rect 1030 348 1034 352
rect 1014 308 1018 312
rect 1070 298 1074 302
rect 1102 458 1106 462
rect 1142 458 1146 462
rect 1174 468 1178 472
rect 1166 448 1170 452
rect 1190 538 1194 542
rect 1238 518 1242 522
rect 1214 488 1218 492
rect 1214 468 1218 472
rect 1238 468 1242 472
rect 1286 568 1290 572
rect 1350 648 1354 652
rect 1318 638 1322 642
rect 1350 638 1354 642
rect 1318 618 1322 622
rect 1270 548 1274 552
rect 1278 468 1282 472
rect 1190 458 1194 462
rect 1230 458 1234 462
rect 1246 458 1250 462
rect 1254 448 1258 452
rect 1190 438 1194 442
rect 1198 438 1202 442
rect 1262 438 1266 442
rect 1222 428 1226 432
rect 1142 418 1146 422
rect 1182 418 1186 422
rect 1150 408 1154 412
rect 1110 388 1114 392
rect 1214 388 1218 392
rect 1158 378 1162 382
rect 1126 348 1130 352
rect 1214 368 1218 372
rect 1182 358 1186 362
rect 1134 338 1138 342
rect 1086 328 1090 332
rect 1182 328 1186 332
rect 1118 308 1122 312
rect 1126 308 1130 312
rect 1086 288 1090 292
rect 1110 288 1114 292
rect 1198 278 1202 282
rect 1038 268 1042 272
rect 1062 268 1066 272
rect 1078 268 1082 272
rect 1046 258 1050 262
rect 1094 248 1098 252
rect 1038 238 1042 242
rect 1006 208 1010 212
rect 958 178 962 182
rect 918 168 922 172
rect 886 158 890 162
rect 862 138 866 142
rect 854 128 858 132
rect 918 138 922 142
rect 1022 158 1026 162
rect 966 148 970 152
rect 1030 148 1034 152
rect 942 128 946 132
rect 958 98 962 102
rect 830 88 834 92
rect 910 88 914 92
rect 926 88 930 92
rect 822 78 826 82
rect 870 68 874 72
rect 862 48 866 52
rect 966 88 970 92
rect 910 68 914 72
rect 926 68 930 72
rect 958 68 962 72
rect 966 58 970 62
rect 1006 128 1010 132
rect 986 103 990 107
rect 993 103 997 107
rect 1006 98 1010 102
rect 1046 158 1050 162
rect 1070 138 1074 142
rect 1062 128 1066 132
rect 1054 88 1058 92
rect 1094 118 1098 122
rect 1134 268 1138 272
rect 1150 268 1154 272
rect 1110 248 1114 252
rect 1118 238 1122 242
rect 1110 168 1114 172
rect 1118 138 1122 142
rect 1102 98 1106 102
rect 1094 88 1098 92
rect 1006 78 1010 82
rect 1014 78 1018 82
rect 1078 78 1082 82
rect 982 58 986 62
rect 902 48 906 52
rect 990 48 994 52
rect 886 28 890 32
rect 894 28 898 32
rect 886 18 890 22
rect 918 18 922 22
rect 934 8 938 12
rect 958 8 962 12
rect 1022 58 1026 62
rect 1182 258 1186 262
rect 1174 248 1178 252
rect 1238 418 1242 422
rect 1318 558 1322 562
rect 1294 548 1298 552
rect 1302 538 1306 542
rect 1294 498 1298 502
rect 1342 548 1346 552
rect 1310 498 1314 502
rect 1302 468 1306 472
rect 1326 458 1330 462
rect 1278 418 1282 422
rect 1286 418 1290 422
rect 1254 408 1258 412
rect 1246 398 1250 402
rect 1262 398 1266 402
rect 1286 378 1290 382
rect 1254 368 1258 372
rect 1302 438 1306 442
rect 1478 848 1482 852
rect 1478 818 1482 822
rect 1438 788 1442 792
rect 1462 758 1466 762
rect 1446 748 1450 752
rect 1446 728 1450 732
rect 1438 648 1442 652
rect 1406 558 1410 562
rect 1358 538 1362 542
rect 1358 458 1362 462
rect 1374 448 1378 452
rect 1470 428 1474 432
rect 1414 418 1418 422
rect 1342 408 1346 412
rect 1342 388 1346 392
rect 1302 378 1306 382
rect 1326 378 1330 382
rect 1358 378 1362 382
rect 1238 358 1242 362
rect 1270 358 1274 362
rect 1294 358 1298 362
rect 1230 308 1234 312
rect 1214 268 1218 272
rect 1222 268 1226 272
rect 1238 268 1242 272
rect 1142 238 1146 242
rect 1150 238 1154 242
rect 1166 238 1170 242
rect 1190 238 1194 242
rect 1222 258 1226 262
rect 1214 248 1218 252
rect 1230 248 1234 252
rect 1198 198 1202 202
rect 1222 198 1226 202
rect 1214 188 1218 192
rect 1230 188 1234 192
rect 1150 168 1154 172
rect 1166 168 1170 172
rect 1142 158 1146 162
rect 1166 158 1170 162
rect 1294 348 1298 352
rect 1246 248 1250 252
rect 1254 238 1258 242
rect 1246 208 1250 212
rect 1278 268 1282 272
rect 1286 258 1290 262
rect 1334 358 1338 362
rect 1318 338 1322 342
rect 1302 248 1306 252
rect 1270 238 1274 242
rect 1302 228 1306 232
rect 1310 218 1314 222
rect 1262 178 1266 182
rect 1294 178 1298 182
rect 1238 168 1242 172
rect 1270 168 1274 172
rect 1294 168 1298 172
rect 1158 148 1162 152
rect 1182 148 1186 152
rect 1198 148 1202 152
rect 1222 148 1226 152
rect 1206 138 1210 142
rect 1222 138 1226 142
rect 1214 128 1218 132
rect 1142 88 1146 92
rect 1182 88 1186 92
rect 1102 78 1106 82
rect 1110 78 1114 82
rect 1158 78 1162 82
rect 1078 68 1082 72
rect 1270 148 1274 152
rect 1254 128 1258 132
rect 1422 388 1426 392
rect 1374 368 1378 372
rect 1390 368 1394 372
rect 1414 368 1418 372
rect 1382 358 1386 362
rect 1398 358 1402 362
rect 1358 348 1362 352
rect 1342 278 1346 282
rect 1358 258 1362 262
rect 1350 238 1354 242
rect 1374 238 1378 242
rect 1358 228 1362 232
rect 1350 208 1354 212
rect 1334 188 1338 192
rect 1318 178 1322 182
rect 1278 78 1282 82
rect 1302 78 1306 82
rect 1374 228 1378 232
rect 1366 218 1370 222
rect 1366 198 1370 202
rect 1326 158 1330 162
rect 1350 158 1354 162
rect 1334 148 1338 152
rect 1326 138 1330 142
rect 1342 128 1346 132
rect 1326 108 1330 112
rect 1118 68 1122 72
rect 1198 68 1202 72
rect 1230 68 1234 72
rect 1302 68 1306 72
rect 1102 58 1106 62
rect 1126 58 1130 62
rect 1142 58 1146 62
rect 1158 58 1162 62
rect 1254 58 1258 62
rect 1062 28 1066 32
rect 1078 18 1082 22
rect 1070 8 1074 12
rect 1166 48 1170 52
rect 1198 48 1202 52
rect 1238 48 1242 52
rect 1262 48 1266 52
rect 1286 48 1290 52
rect 1278 38 1282 42
rect 1238 28 1242 32
rect 1166 18 1170 22
rect 1382 208 1386 212
rect 1382 198 1386 202
rect 1406 328 1410 332
rect 1406 318 1410 322
rect 1414 278 1418 282
rect 1422 248 1426 252
rect 1414 238 1418 242
rect 1390 158 1394 162
rect 1406 148 1410 152
rect 1366 138 1370 142
rect 1382 128 1386 132
rect 1390 118 1394 122
rect 1382 98 1386 102
rect 1374 78 1378 82
rect 1454 378 1458 382
rect 1478 338 1482 342
rect 1454 298 1458 302
rect 1446 248 1450 252
rect 1446 238 1450 242
rect 1406 88 1410 92
rect 1430 78 1434 82
rect 1470 288 1474 292
rect 1478 278 1482 282
rect 1478 168 1482 172
rect 1478 108 1482 112
rect 1422 68 1426 72
rect 1358 48 1362 52
rect 1334 38 1338 42
<< metal3 >>
rect 346 1408 350 1411
rect 618 1408 654 1411
rect 722 1408 726 1411
rect 882 1408 886 1411
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 486 1403 488 1407
rect 530 1398 726 1401
rect 730 1398 758 1401
rect 762 1398 1334 1401
rect 426 1388 998 1391
rect 1002 1388 1062 1391
rect 346 1378 377 1381
rect 514 1378 718 1381
rect 722 1378 742 1381
rect 746 1378 774 1381
rect 778 1378 1358 1381
rect 282 1368 366 1371
rect 374 1371 377 1378
rect 374 1368 694 1371
rect 698 1368 798 1371
rect 802 1368 1177 1371
rect 1266 1368 1294 1371
rect 58 1358 94 1361
rect 114 1358 118 1361
rect 138 1358 142 1361
rect 218 1358 262 1361
rect 270 1361 273 1368
rect 1174 1362 1177 1368
rect 270 1358 438 1361
rect 458 1358 478 1361
rect 554 1358 654 1361
rect 770 1358 814 1361
rect 922 1358 1046 1361
rect 1050 1358 1118 1361
rect 1158 1358 1166 1361
rect 1194 1358 1214 1361
rect 1234 1358 1310 1361
rect 1378 1358 1398 1361
rect 1418 1358 1430 1361
rect 202 1348 222 1351
rect 226 1348 238 1351
rect 250 1348 286 1351
rect 290 1348 326 1351
rect 330 1348 350 1351
rect 354 1348 398 1351
rect 402 1348 454 1351
rect 602 1348 622 1351
rect 634 1348 638 1351
rect 762 1348 790 1351
rect 794 1348 814 1351
rect 818 1348 878 1351
rect 882 1348 902 1351
rect 906 1348 950 1351
rect 954 1348 1014 1351
rect 1074 1348 1110 1351
rect 1130 1348 1262 1351
rect 1362 1348 1382 1351
rect 34 1338 62 1341
rect 66 1338 102 1341
rect 106 1338 150 1341
rect 154 1338 185 1341
rect 226 1338 257 1341
rect 282 1338 334 1341
rect 362 1338 382 1341
rect 482 1338 510 1341
rect 646 1341 649 1348
rect 646 1338 678 1341
rect 682 1338 694 1341
rect 842 1338 889 1341
rect 914 1338 974 1341
rect 1034 1338 1190 1341
rect 1298 1338 1318 1341
rect 1322 1338 1350 1341
rect 1354 1338 1430 1341
rect 182 1332 185 1338
rect 254 1332 257 1338
rect 614 1332 617 1338
rect 886 1332 889 1338
rect -26 1331 -22 1332
rect -26 1328 6 1331
rect 82 1328 86 1331
rect 394 1328 398 1331
rect 730 1328 774 1331
rect 906 1328 942 1331
rect 946 1328 1046 1331
rect 1054 1328 1086 1331
rect 1146 1328 1166 1331
rect 1054 1322 1057 1328
rect 10 1318 230 1321
rect 266 1318 270 1321
rect 314 1318 718 1321
rect 722 1318 726 1321
rect 730 1318 782 1321
rect 786 1318 1022 1321
rect 1066 1318 1094 1321
rect 1098 1318 1134 1321
rect 1138 1318 1158 1321
rect 1178 1318 1206 1321
rect 1210 1318 1262 1321
rect 1266 1318 1390 1321
rect 1394 1318 1454 1321
rect 1454 1312 1457 1318
rect -26 1311 -22 1312
rect -26 1308 6 1311
rect 10 1308 62 1311
rect 66 1308 118 1311
rect 122 1308 222 1311
rect 258 1308 350 1311
rect 354 1308 846 1311
rect 850 1308 854 1311
rect 858 1308 894 1311
rect 970 1308 974 1311
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 146 1298 222 1301
rect 234 1298 558 1301
rect 562 1298 638 1301
rect 810 1298 822 1301
rect 834 1298 862 1301
rect 178 1288 678 1291
rect 682 1288 766 1291
rect 770 1288 1230 1291
rect 1330 1288 1438 1291
rect 226 1278 230 1281
rect 234 1278 310 1281
rect 314 1278 334 1281
rect 386 1278 414 1281
rect 418 1278 446 1281
rect 450 1278 526 1281
rect 530 1278 534 1281
rect 538 1278 574 1281
rect 618 1278 630 1281
rect 642 1278 950 1281
rect 954 1278 958 1281
rect 1018 1278 1038 1281
rect 1226 1278 1318 1281
rect 1378 1278 1430 1281
rect 126 1272 129 1278
rect -26 1271 -22 1272
rect -26 1268 38 1271
rect 106 1268 110 1271
rect 226 1268 590 1271
rect 606 1268 614 1271
rect 618 1268 622 1271
rect 818 1268 1102 1271
rect 1202 1268 1230 1271
rect 1394 1268 1414 1271
rect 118 1261 121 1268
rect 54 1258 81 1261
rect 118 1258 126 1261
rect 190 1261 193 1268
rect 186 1258 193 1261
rect 226 1258 238 1261
rect 282 1258 318 1261
rect 354 1258 526 1261
rect 530 1258 662 1261
rect 706 1258 742 1261
rect 806 1258 830 1261
rect 842 1258 1070 1261
rect 1118 1261 1121 1268
rect 1118 1258 1182 1261
rect 1202 1258 1246 1261
rect 1318 1261 1321 1268
rect 1342 1261 1345 1268
rect 1318 1258 1345 1261
rect 1402 1258 1422 1261
rect 54 1252 57 1258
rect 78 1252 81 1258
rect 806 1252 809 1258
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 34 1248 46 1251
rect 90 1248 118 1251
rect 122 1248 174 1251
rect 178 1248 254 1251
rect 282 1248 302 1251
rect 394 1248 462 1251
rect 482 1248 502 1251
rect 522 1248 534 1251
rect 538 1248 582 1251
rect 586 1248 622 1251
rect 626 1248 702 1251
rect 854 1248 878 1251
rect 898 1248 902 1251
rect 914 1248 918 1251
rect 1086 1251 1089 1258
rect 1086 1248 1142 1251
rect 1162 1248 1190 1251
rect 1194 1248 1254 1251
rect 1258 1248 1318 1251
rect 1322 1248 1422 1251
rect 1502 1248 1506 1252
rect 854 1242 857 1248
rect 202 1238 214 1241
rect 226 1238 446 1241
rect 450 1238 838 1241
rect 906 1238 1038 1241
rect 1058 1238 1126 1241
rect 1250 1238 1278 1241
rect 1282 1238 1342 1241
rect 1346 1238 1374 1241
rect 1502 1241 1505 1248
rect 1378 1238 1505 1241
rect 298 1228 422 1231
rect 610 1228 654 1231
rect 890 1228 918 1231
rect 1146 1228 1254 1231
rect 1290 1228 1318 1231
rect 1386 1228 1409 1231
rect 1418 1228 1449 1231
rect 1406 1222 1409 1228
rect 1446 1222 1449 1228
rect 594 1218 814 1221
rect 834 1218 910 1221
rect 914 1218 974 1221
rect 930 1208 950 1211
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 486 1203 488 1207
rect 74 1198 86 1201
rect 98 1198 158 1201
rect 266 1198 382 1201
rect 1146 1198 1358 1201
rect 42 1188 486 1191
rect 626 1188 630 1191
rect 926 1191 929 1198
rect 874 1188 929 1191
rect 18 1178 38 1181
rect 138 1178 142 1181
rect 410 1178 654 1181
rect 658 1178 1142 1181
rect 1238 1181 1241 1188
rect 1238 1178 1286 1181
rect 126 1172 129 1178
rect 1302 1172 1305 1178
rect -26 1171 -22 1172
rect -26 1168 49 1171
rect 626 1168 710 1171
rect 882 1168 886 1171
rect 906 1168 910 1171
rect 946 1168 985 1171
rect 1122 1168 1158 1171
rect 1258 1168 1281 1171
rect 1330 1168 1358 1171
rect 1434 1168 1438 1171
rect 46 1162 49 1168
rect 270 1162 273 1168
rect 50 1158 134 1161
rect 138 1158 198 1161
rect 202 1158 246 1161
rect 298 1158 350 1161
rect 418 1158 510 1161
rect 746 1158 750 1161
rect 830 1161 833 1168
rect 982 1162 985 1168
rect 1278 1162 1281 1168
rect 810 1158 833 1161
rect 882 1158 894 1161
rect 1002 1158 1022 1161
rect 1106 1158 1134 1161
rect 1210 1158 1254 1161
rect 1298 1158 1334 1161
rect 1370 1158 1382 1161
rect 1502 1161 1506 1162
rect 1402 1158 1506 1161
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 50 1148 54 1151
rect 82 1148 94 1151
rect 138 1148 142 1151
rect 286 1151 289 1158
rect 158 1148 289 1151
rect 306 1148 457 1151
rect 642 1148 662 1151
rect 710 1151 713 1158
rect 682 1148 713 1151
rect 722 1148 1134 1151
rect 1138 1148 1398 1151
rect 158 1142 161 1148
rect 454 1142 457 1148
rect 66 1138 150 1141
rect 230 1138 238 1141
rect 242 1138 326 1141
rect 330 1138 414 1141
rect 458 1138 462 1141
rect 474 1138 534 1141
rect 538 1138 614 1141
rect 618 1138 686 1141
rect 690 1138 718 1141
rect 722 1138 750 1141
rect 802 1138 822 1141
rect 858 1138 910 1141
rect 930 1138 1094 1141
rect 1290 1138 1310 1141
rect 1362 1138 1390 1141
rect 1410 1138 1430 1141
rect 1434 1138 1438 1141
rect 1442 1138 1446 1141
rect 1450 1138 1462 1141
rect 1474 1138 1478 1141
rect 1502 1141 1506 1142
rect 1482 1138 1506 1141
rect 194 1128 302 1131
rect 306 1128 358 1131
rect 434 1128 478 1131
rect 498 1128 502 1131
rect 522 1128 550 1131
rect 554 1128 638 1131
rect 1010 1128 1014 1131
rect 1026 1128 1182 1131
rect 1186 1128 1326 1131
rect 1370 1128 1446 1131
rect 114 1118 238 1121
rect 426 1118 462 1121
rect 518 1121 521 1128
rect 590 1122 593 1128
rect 466 1118 521 1121
rect 578 1118 582 1121
rect 706 1118 766 1121
rect 810 1118 862 1121
rect 874 1118 1054 1121
rect 1058 1118 1198 1121
rect 346 1108 350 1111
rect 354 1108 630 1111
rect 1042 1108 1102 1111
rect 1178 1108 1342 1111
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 154 1098 286 1101
rect 386 1098 430 1101
rect 618 1098 646 1101
rect 650 1098 670 1101
rect 1010 1098 1222 1101
rect 202 1088 393 1091
rect 594 1088 606 1091
rect 634 1088 849 1091
rect 978 1088 1086 1091
rect 1090 1088 1142 1091
rect 1502 1091 1506 1092
rect 1474 1088 1506 1091
rect 390 1082 393 1088
rect 846 1082 849 1088
rect 246 1078 334 1081
rect 394 1078 398 1081
rect 506 1078 558 1081
rect 746 1078 750 1081
rect 850 1078 854 1081
rect 942 1078 966 1081
rect 1050 1078 1086 1081
rect 1106 1078 1190 1081
rect 1226 1078 1246 1081
rect 1326 1081 1329 1088
rect 1250 1078 1329 1081
rect 1354 1078 1374 1081
rect 1402 1078 1406 1081
rect 246 1072 249 1078
rect 382 1072 385 1078
rect 194 1068 198 1071
rect 490 1068 494 1071
rect 610 1068 694 1071
rect 918 1071 921 1078
rect 906 1068 921 1071
rect 942 1072 945 1078
rect 1014 1071 1017 1078
rect 1014 1068 1070 1071
rect 1178 1068 1182 1071
rect 1274 1068 1286 1071
rect 1306 1068 1310 1071
rect 1382 1071 1385 1078
rect 1370 1068 1385 1071
rect 1502 1071 1506 1072
rect 1402 1068 1506 1071
rect 106 1058 110 1061
rect 170 1058 182 1061
rect 258 1058 270 1061
rect 318 1061 321 1068
rect 306 1058 321 1061
rect 502 1061 505 1068
rect 502 1058 518 1061
rect 538 1058 550 1061
rect 570 1058 598 1061
rect 830 1061 833 1068
rect 794 1058 833 1061
rect 842 1058 886 1061
rect 890 1058 1014 1061
rect 1118 1061 1121 1068
rect 1106 1058 1121 1061
rect 1202 1058 1270 1061
rect 1286 1058 1294 1061
rect 1298 1058 1334 1061
rect 1342 1061 1345 1068
rect 1342 1058 1374 1061
rect 1378 1058 1414 1061
rect 1442 1058 1449 1061
rect 1422 1052 1425 1058
rect 1446 1052 1449 1058
rect -26 1051 -22 1052
rect -26 1048 62 1051
rect 154 1048 206 1051
rect 242 1048 246 1051
rect 266 1048 273 1051
rect 306 1048 326 1051
rect 538 1048 542 1051
rect 578 1048 606 1051
rect 610 1048 646 1051
rect 650 1048 654 1051
rect 858 1048 870 1051
rect 882 1048 894 1051
rect 922 1048 1046 1051
rect 1266 1048 1318 1051
rect 1502 1051 1506 1052
rect 1482 1048 1506 1051
rect 50 1038 102 1041
rect 146 1038 262 1041
rect 270 1041 273 1048
rect 270 1038 305 1041
rect 438 1041 441 1048
rect 426 1038 441 1041
rect 626 1038 734 1041
rect 870 1038 878 1041
rect 882 1038 886 1041
rect 1114 1038 1150 1041
rect 1350 1041 1353 1048
rect 1282 1038 1353 1041
rect 1442 1038 1454 1041
rect 138 1028 166 1031
rect 274 1028 294 1031
rect 302 1031 305 1038
rect 302 1028 518 1031
rect 642 1028 646 1031
rect 810 1028 926 1031
rect 938 1028 1398 1031
rect 74 1018 150 1021
rect 338 1018 681 1021
rect 830 1018 838 1021
rect 842 1018 854 1021
rect 1042 1018 1049 1021
rect 1214 1018 1222 1021
rect 1226 1018 1358 1021
rect 1366 1018 1430 1021
rect 678 1012 681 1018
rect 1046 1012 1049 1018
rect 290 1008 334 1011
rect 530 1008 582 1011
rect 682 1008 934 1011
rect 1210 1008 1254 1011
rect 1258 1008 1262 1011
rect 1366 1011 1369 1018
rect 1338 1008 1369 1011
rect 1502 1011 1506 1012
rect 1394 1008 1506 1011
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 486 1003 488 1007
rect 290 998 406 1001
rect 450 998 462 1001
rect 562 998 654 1001
rect 850 998 862 1001
rect 1050 998 1094 1001
rect 1146 998 1470 1001
rect 226 988 270 991
rect 274 988 281 991
rect 314 988 446 991
rect 578 988 598 991
rect 866 988 966 991
rect 970 988 1062 991
rect 1346 988 1374 991
rect 1502 991 1506 992
rect 1410 988 1506 991
rect 202 978 246 981
rect 258 978 270 981
rect 274 978 302 981
rect 354 978 494 981
rect 498 978 574 981
rect 630 981 633 988
rect 594 978 633 981
rect 714 978 726 981
rect 854 981 857 988
rect 854 978 910 981
rect 930 978 1070 981
rect 1150 978 1390 981
rect 1150 972 1153 978
rect 130 968 206 971
rect 258 968 262 971
rect 330 968 342 971
rect 466 968 614 971
rect 626 968 630 971
rect 642 968 806 971
rect 810 968 830 971
rect 834 968 1150 971
rect 1178 968 1182 971
rect 1306 968 1326 971
rect 1370 968 1430 971
rect 1502 971 1506 972
rect 1482 968 1506 971
rect 118 961 121 968
rect 118 958 126 961
rect 166 958 174 961
rect 178 958 238 961
rect 338 958 390 961
rect 434 958 502 961
rect 634 958 654 961
rect 666 958 710 961
rect 746 958 774 961
rect 838 958 854 961
rect 954 958 982 961
rect 1042 958 1054 961
rect 1250 958 1254 961
rect 1330 958 1334 961
rect 1442 958 1446 961
rect -26 951 -22 952
rect -26 948 6 951
rect 94 951 97 958
rect 94 948 174 951
rect 258 948 318 951
rect 342 948 369 951
rect 450 948 462 951
rect 542 951 545 958
rect 530 948 545 951
rect 586 948 606 951
rect 654 951 657 958
rect 654 948 734 951
rect 798 951 801 958
rect 786 948 801 951
rect 838 952 841 958
rect 902 951 905 958
rect 890 948 905 951
rect 934 951 937 958
rect 930 948 937 951
rect 1026 948 1054 951
rect 1058 948 1134 951
rect 1210 948 1238 951
rect 1266 948 1318 951
rect 1322 948 1342 951
rect 1374 951 1377 958
rect 1502 951 1506 952
rect 1362 948 1377 951
rect 1390 948 1506 951
rect 342 942 345 948
rect 366 942 369 948
rect 410 938 446 941
rect 458 938 510 941
rect 562 938 566 941
rect 602 938 654 941
rect 674 938 822 941
rect 826 938 958 941
rect 962 938 1222 941
rect 1390 941 1393 948
rect 1226 938 1393 941
rect 1402 938 1406 941
rect 1410 938 1446 941
rect 1450 938 1454 941
rect 134 932 137 938
rect 154 928 166 931
rect 538 928 590 931
rect 730 928 798 931
rect 802 928 814 931
rect 818 928 838 931
rect 850 928 1097 931
rect 1178 928 1214 931
rect 1290 928 1294 931
rect 1322 928 1358 931
rect 1386 928 1390 931
rect 1394 928 1478 931
rect 1502 928 1506 932
rect 1094 922 1097 928
rect 362 918 390 921
rect 538 918 1086 921
rect 1106 918 1254 921
rect 1362 918 1406 921
rect 1502 921 1505 928
rect 1442 918 1505 921
rect 130 908 142 911
rect 162 908 174 911
rect 354 908 390 911
rect 538 908 566 911
rect 634 908 846 911
rect 874 908 950 911
rect 1138 908 1206 911
rect 1322 908 1366 911
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 506 898 534 901
rect 794 898 822 901
rect 1090 898 1142 901
rect 1242 898 1270 901
rect 1274 898 1438 901
rect -26 891 -22 892
rect -26 888 166 891
rect 378 888 702 891
rect 706 888 1238 891
rect 1502 891 1506 892
rect 1258 888 1506 891
rect 282 878 430 881
rect 530 878 622 881
rect 714 878 734 881
rect 842 878 926 881
rect 986 878 998 881
rect 1002 878 1102 881
rect 1298 878 1398 881
rect -26 871 -22 872
rect 6 871 9 878
rect -26 868 9 871
rect 322 868 326 871
rect 338 868 358 871
rect 362 868 374 871
rect 378 868 398 871
rect 426 868 438 871
rect 522 868 550 871
rect 554 868 598 871
rect 690 868 718 871
rect 794 868 798 871
rect 866 868 878 871
rect 1074 868 1110 871
rect 1194 868 1198 871
rect 1218 868 1294 871
rect 1298 868 1302 871
rect 1422 871 1425 878
rect 1314 868 1425 871
rect 142 862 145 868
rect 310 861 313 868
rect 298 858 313 861
rect 558 858 577 861
rect 586 858 598 861
rect 618 858 646 861
rect 698 858 742 861
rect 758 861 761 868
rect 774 861 777 868
rect 758 858 777 861
rect 850 858 870 861
rect 1182 861 1185 868
rect 1170 858 1185 861
rect -26 848 -22 852
rect 98 848 142 851
rect 354 848 358 851
rect 430 851 433 858
rect 410 848 433 851
rect 558 852 561 858
rect 574 852 577 858
rect 582 848 718 851
rect 878 851 881 858
rect 1046 852 1049 858
rect 722 848 881 851
rect 898 848 942 851
rect 1102 851 1105 858
rect 1074 848 1142 851
rect 1322 848 1326 851
rect 1350 851 1353 858
rect 1406 852 1409 858
rect 1338 848 1353 851
rect 1370 848 1374 851
rect 1502 851 1506 852
rect 1482 848 1506 851
rect -26 841 -23 848
rect -26 838 278 841
rect 306 838 350 841
rect 394 838 526 841
rect 582 841 585 848
rect 570 838 585 841
rect 642 838 646 841
rect 666 838 686 841
rect 754 838 838 841
rect 858 838 862 841
rect 874 838 1070 841
rect 1178 838 1214 841
rect 1290 838 1294 841
rect 1314 838 1326 841
rect 1390 841 1393 848
rect 1346 838 1393 841
rect -26 831 -22 832
rect -26 828 6 831
rect 250 828 430 831
rect 442 828 982 831
rect 1018 828 1118 831
rect 466 818 926 821
rect 930 818 1046 821
rect 1050 818 1478 821
rect -26 811 -22 812
rect -26 808 30 811
rect 498 808 790 811
rect 802 808 886 811
rect 946 808 1054 811
rect 1202 808 1366 811
rect 472 803 474 807
rect 478 803 481 807
rect 486 803 488 807
rect 594 798 614 801
rect 626 798 630 801
rect 642 798 646 801
rect 658 798 670 801
rect 698 798 814 801
rect 818 798 854 801
rect 858 798 870 801
rect 874 798 1030 801
rect 1274 798 1302 801
rect 1314 798 1326 801
rect 1502 801 1506 802
rect 1482 798 1506 801
rect -26 791 -22 792
rect -26 788 78 791
rect 458 788 462 791
rect 530 788 934 791
rect 954 788 1022 791
rect 1034 788 1158 791
rect 1298 788 1318 791
rect 50 778 174 781
rect 442 778 726 781
rect 738 778 798 781
rect 842 778 870 781
rect 878 778 902 781
rect 938 778 1390 781
rect 1438 781 1441 788
rect 1502 781 1506 782
rect 1438 778 1506 781
rect -26 771 -22 772
rect -26 768 62 771
rect 178 768 222 771
rect 402 768 494 771
rect 626 768 710 771
rect 722 768 742 771
rect 782 768 790 771
rect 810 768 814 771
rect 878 771 881 778
rect 826 768 881 771
rect 890 768 998 771
rect 1002 768 1094 771
rect 1162 768 1254 771
rect 1290 768 1294 771
rect 1322 768 1358 771
rect 138 758 262 761
rect 266 758 382 761
rect 386 758 798 761
rect 874 758 878 761
rect 962 758 1030 761
rect 1122 758 1214 761
rect 1218 758 1334 761
rect 1378 758 1462 761
rect 1502 761 1506 762
rect 1466 758 1506 761
rect -26 751 -22 752
rect -26 748 14 751
rect 54 751 57 758
rect 34 748 57 751
rect 66 748 230 751
rect 246 748 342 751
rect 366 748 422 751
rect 434 748 550 751
rect 554 748 870 751
rect 918 751 921 758
rect 1086 752 1089 758
rect 914 748 921 751
rect 1018 748 1033 751
rect 246 742 249 748
rect 366 742 369 748
rect 1030 742 1033 748
rect 122 738 161 741
rect 158 732 161 738
rect 538 738 574 741
rect 586 738 606 741
rect 634 738 670 741
rect 690 738 694 741
rect 706 738 758 741
rect 770 738 774 741
rect 810 738 830 741
rect 866 738 958 741
rect 1314 738 1358 741
rect 1446 741 1449 748
rect 1386 738 1449 741
rect 166 732 169 738
rect -26 728 -22 732
rect 322 728 406 731
rect 514 728 558 731
rect 618 728 646 731
rect 682 728 718 731
rect 730 728 734 731
rect 810 728 961 731
rect 970 728 1358 731
rect 1502 731 1506 732
rect 1450 728 1506 731
rect -26 721 -23 728
rect -26 718 222 721
rect 226 718 462 721
rect 466 718 910 721
rect 958 721 961 728
rect 958 718 1182 721
rect -26 711 -22 712
rect -26 708 142 711
rect 146 708 550 711
rect 554 708 750 711
rect 754 708 830 711
rect 886 708 966 711
rect 1502 711 1506 712
rect 1210 708 1506 711
rect 338 698 446 701
rect 450 698 622 701
rect 626 698 686 701
rect 690 698 702 701
rect 886 701 889 708
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 730 698 889 701
rect 898 698 950 701
rect 1234 698 1505 701
rect 1502 692 1505 698
rect -26 688 -22 692
rect 10 688 334 691
rect 346 688 758 691
rect 906 688 1038 691
rect 1306 688 1318 691
rect 1502 688 1506 692
rect -26 681 -23 688
rect -26 678 17 681
rect 50 678 102 681
rect 106 678 190 681
rect 618 678 654 681
rect 682 678 758 681
rect 770 678 782 681
rect 922 678 926 681
rect 1058 678 1118 681
rect 1298 678 1318 681
rect -26 671 -22 672
rect -26 668 6 671
rect 14 671 17 678
rect 14 668 54 671
rect 70 668 94 671
rect 130 668 166 671
rect 234 668 246 671
rect 250 668 342 671
rect 442 668 462 671
rect 534 671 537 678
rect 522 668 537 671
rect 562 668 566 671
rect 602 668 686 671
rect 722 668 734 671
rect 754 668 766 671
rect 810 668 814 671
rect 850 668 854 671
rect 890 668 1118 671
rect 1262 671 1265 678
rect 1258 668 1265 671
rect 1298 668 1302 671
rect 1502 671 1506 672
rect 1482 668 1506 671
rect 70 662 73 668
rect 702 662 705 668
rect 1270 662 1273 668
rect 82 658 118 661
rect 122 658 550 661
rect 654 658 670 661
rect 762 658 814 661
rect 858 658 862 661
rect 874 658 1025 661
rect 1250 658 1254 661
rect 1290 658 1353 661
rect -26 648 -22 652
rect 42 648 86 651
rect 114 648 166 651
rect 170 648 214 651
rect 266 648 286 651
rect 362 648 366 651
rect 402 648 462 651
rect 466 648 598 651
rect 630 651 633 658
rect 602 648 633 651
rect 638 652 641 658
rect 654 652 657 658
rect 686 652 689 658
rect 1022 652 1025 658
rect 1350 652 1353 658
rect 698 648 798 651
rect 1282 648 1310 651
rect 1502 651 1506 652
rect 1442 648 1506 651
rect -26 641 -23 648
rect -26 638 302 641
rect 306 638 366 641
rect 370 638 462 641
rect 466 638 590 641
rect 658 638 662 641
rect 682 638 894 641
rect 1098 638 1214 641
rect 1322 638 1350 641
rect 670 632 673 638
rect 18 628 230 631
rect 278 628 318 631
rect 342 628 350 631
rect 354 628 382 631
rect 394 628 422 631
rect 474 628 494 631
rect 522 628 550 631
rect 562 628 606 631
rect 802 628 870 631
rect 874 628 990 631
rect 278 622 281 628
rect 298 618 318 621
rect 330 618 390 621
rect 394 618 401 621
rect 418 618 526 621
rect 586 618 630 621
rect 850 618 1318 621
rect 58 608 366 611
rect 554 608 1014 611
rect 472 603 474 607
rect 478 603 481 607
rect 486 603 488 607
rect 274 598 294 601
rect 346 598 414 601
rect 530 598 606 601
rect 610 598 622 601
rect 458 588 534 591
rect -26 578 -22 582
rect 78 581 81 588
rect 78 578 150 581
rect 162 578 166 581
rect 346 578 494 581
rect 498 578 550 581
rect 554 578 654 581
rect -26 571 -23 578
rect -26 568 110 571
rect 134 568 142 571
rect 146 568 158 571
rect 274 568 318 571
rect 410 568 502 571
rect 514 568 518 571
rect 682 568 718 571
rect 938 568 1102 571
rect 1114 568 1150 571
rect 1218 568 1222 571
rect 1242 568 1254 571
rect 1282 568 1286 571
rect 110 562 113 568
rect 126 562 129 568
rect 174 562 177 568
rect -26 561 -22 562
rect -26 558 54 561
rect 82 558 86 561
rect 138 558 174 561
rect 242 558 334 561
rect 394 558 502 561
rect 922 558 942 561
rect 1002 558 1118 561
rect 1170 558 1262 561
rect 34 548 38 551
rect 70 551 73 558
rect 70 548 86 551
rect 106 548 126 551
rect 130 548 206 551
rect 210 548 222 551
rect 350 551 353 558
rect 346 548 353 551
rect 386 548 702 551
rect 706 548 774 551
rect 838 551 841 558
rect 1318 552 1321 558
rect 794 548 841 551
rect 1062 548 1070 551
rect 1074 548 1150 551
rect 1274 548 1294 551
rect 1406 551 1409 558
rect 1346 548 1409 551
rect -26 541 -22 542
rect -26 538 6 541
rect 58 538 62 541
rect 90 538 126 541
rect 154 538 158 541
rect 170 538 174 541
rect 186 538 206 541
rect 274 538 294 541
rect 406 538 422 541
rect 458 538 462 541
rect 634 538 646 541
rect 770 538 798 541
rect 802 538 918 541
rect 922 538 950 541
rect 954 538 958 541
rect 962 538 998 541
rect 1026 538 1046 541
rect 1058 538 1190 541
rect 1274 538 1302 541
rect 1346 538 1358 541
rect 366 532 369 538
rect 406 532 409 538
rect 566 532 569 538
rect 138 528 150 531
rect 234 528 238 531
rect 282 528 286 531
rect 758 531 761 538
rect 666 528 974 531
rect 1050 528 1070 531
rect 1074 528 1142 531
rect 46 522 49 528
rect 66 518 750 521
rect 754 518 942 521
rect 946 518 1054 521
rect 1094 518 1102 521
rect 1106 518 1238 521
rect 314 508 502 511
rect 578 508 630 511
rect 642 508 702 511
rect 810 508 830 511
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 170 498 198 501
rect 290 498 382 501
rect 386 498 430 501
rect 778 498 806 501
rect 1298 498 1310 501
rect -26 491 -22 492
rect -26 488 6 491
rect 10 488 278 491
rect 298 488 334 491
rect 338 488 366 491
rect 466 488 494 491
rect 562 488 614 491
rect 626 488 678 491
rect 682 488 990 491
rect 998 488 1078 491
rect 1114 488 1118 491
rect 1122 488 1214 491
rect 1218 488 1246 491
rect 98 478 126 481
rect 378 478 398 481
rect 458 478 462 481
rect 506 478 510 481
rect 614 481 617 488
rect 614 478 662 481
rect 666 478 694 481
rect 698 478 710 481
rect 778 478 942 481
rect 998 481 1001 488
rect 946 478 1001 481
rect 1090 478 1110 481
rect 1138 478 1158 481
rect 342 472 345 478
rect -26 471 -22 472
rect -26 468 6 471
rect 34 468 54 471
rect 362 468 382 471
rect 398 471 401 478
rect 398 468 414 471
rect 442 468 470 471
rect 554 468 582 471
rect 742 468 745 478
rect 758 472 761 478
rect 786 468 790 471
rect 826 468 846 471
rect 1026 468 1038 471
rect 42 458 78 461
rect 118 461 121 468
rect 166 461 169 468
rect 118 458 169 461
rect 218 458 230 461
rect 262 461 265 468
rect 662 462 665 468
rect 250 458 265 461
rect 378 458 457 461
rect 538 458 566 461
rect 570 458 622 461
rect 738 458 790 461
rect 794 458 870 461
rect 926 461 929 468
rect 1102 462 1105 471
rect 1114 468 1118 471
rect 1178 468 1214 471
rect 1234 468 1238 471
rect 1282 468 1302 471
rect 890 458 929 461
rect 986 458 1030 461
rect 1050 458 1070 461
rect 1134 461 1137 468
rect 1134 458 1142 461
rect 1194 458 1230 461
rect 1234 458 1246 461
rect 1250 458 1326 461
rect 1362 458 1377 461
rect -26 451 -22 452
rect -26 448 70 451
rect 122 448 214 451
rect 362 448 366 451
rect 454 451 457 458
rect 426 448 449 451
rect 454 448 598 451
rect 650 448 654 451
rect 726 451 729 458
rect 1374 452 1377 458
rect 726 448 790 451
rect 794 448 966 451
rect 1042 448 1062 451
rect 1082 448 1166 451
rect 446 442 449 448
rect 146 438 150 441
rect 210 438 238 441
rect 258 438 294 441
rect 522 438 542 441
rect 762 438 806 441
rect 866 438 878 441
rect 898 438 918 441
rect 1194 438 1198 441
rect 1254 441 1257 448
rect 1254 438 1262 441
rect 1298 438 1302 441
rect 574 432 577 438
rect 10 428 182 431
rect 186 428 374 431
rect 514 428 518 431
rect 842 428 966 431
rect 1226 428 1470 431
rect 74 418 318 421
rect 322 418 726 421
rect 730 418 1022 421
rect 1146 418 1182 421
rect 1186 418 1201 421
rect 1242 418 1278 421
rect 1290 418 1414 421
rect 70 408 190 411
rect 194 408 278 411
rect 282 408 294 411
rect 506 408 558 411
rect 562 408 702 411
rect 794 408 814 411
rect 882 408 950 411
rect 954 408 974 411
rect 1050 408 1150 411
rect 1198 411 1201 418
rect 1198 408 1254 411
rect 1258 408 1342 411
rect 46 402 49 408
rect 70 402 73 408
rect 472 403 474 407
rect 478 403 481 407
rect 486 403 488 407
rect 58 398 70 401
rect 498 398 550 401
rect 770 398 838 401
rect 922 398 934 401
rect 1250 398 1262 401
rect 122 388 134 391
rect 138 388 166 391
rect 210 388 246 391
rect 514 388 1110 391
rect 1218 388 1318 391
rect 1346 388 1422 391
rect -26 381 -22 382
rect -26 378 118 381
rect 414 381 417 388
rect 394 378 417 381
rect 426 378 590 381
rect 602 378 886 381
rect 890 378 1158 381
rect 1306 378 1326 381
rect 1330 378 1358 381
rect 130 368 134 371
rect 194 368 222 371
rect 258 368 318 371
rect 338 368 374 371
rect 402 368 454 371
rect 490 368 550 371
rect 658 368 910 371
rect 1042 368 1078 371
rect 1286 371 1289 378
rect 1286 368 1374 371
rect 1382 368 1390 371
rect 1454 371 1457 378
rect 1418 368 1457 371
rect 98 358 102 361
rect 150 361 153 368
rect 138 358 190 361
rect 310 358 350 361
rect 378 358 438 361
rect 514 358 518 361
rect 586 358 606 361
rect 674 358 774 361
rect 794 358 806 361
rect 874 358 926 361
rect 954 358 1022 361
rect 1214 361 1217 368
rect 1254 362 1257 368
rect 1382 362 1385 368
rect 1214 358 1238 361
rect 1274 358 1278 361
rect 1298 358 1334 361
rect 1402 358 1454 361
rect 1502 361 1506 362
rect 1482 358 1506 361
rect -26 348 -22 352
rect 6 348 14 351
rect 18 348 22 351
rect 26 348 46 351
rect 74 348 94 351
rect 262 351 265 358
rect 250 348 265 351
rect 310 352 313 358
rect 614 351 617 358
rect 838 352 841 358
rect 578 348 617 351
rect 698 348 774 351
rect 810 348 814 351
rect 902 348 918 351
rect 1046 351 1049 358
rect 1034 348 1049 351
rect 1130 348 1166 351
rect 1182 351 1185 358
rect 1334 352 1337 358
rect 1182 348 1238 351
rect 1250 348 1294 351
rect 1354 348 1358 351
rect -26 341 -23 348
rect 454 342 457 348
rect 790 342 793 348
rect 902 342 905 348
rect -26 338 78 341
rect 114 338 158 341
rect 218 338 246 341
rect 282 338 286 341
rect 714 338 726 341
rect 826 338 862 341
rect 914 338 950 341
rect 1138 338 1198 341
rect 1202 338 1318 341
rect 1502 341 1506 342
rect 1482 338 1506 341
rect 566 332 569 338
rect 26 328 278 331
rect 282 328 318 331
rect 378 328 430 331
rect 434 328 462 331
rect 474 328 510 331
rect 546 328 550 331
rect 602 328 654 331
rect 690 328 742 331
rect 770 328 990 331
rect 1074 328 1086 331
rect 1186 328 1246 331
rect 1410 328 1478 331
rect 82 318 494 321
rect 498 318 574 321
rect 578 318 662 321
rect 682 318 710 321
rect 714 318 1406 321
rect 354 308 678 311
rect 754 308 838 311
rect 850 308 870 311
rect 874 308 942 311
rect 1018 308 1118 311
rect 1130 308 1230 311
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 58 298 446 301
rect 514 298 929 301
rect 1010 298 1070 301
rect 1074 298 1454 301
rect 926 292 929 298
rect -26 291 -22 292
rect -26 288 6 291
rect 10 288 510 291
rect 530 288 582 291
rect 650 288 654 291
rect 930 288 1086 291
rect 1114 288 1470 291
rect 26 278 38 281
rect 162 278 270 281
rect 322 278 342 281
rect 370 278 374 281
rect 378 278 390 281
rect 450 278 454 281
rect 466 278 518 281
rect 522 278 534 281
rect 538 278 622 281
rect 626 278 638 281
rect 770 278 774 281
rect 1018 278 1198 281
rect 1346 278 1414 281
rect 1502 281 1506 282
rect 1482 278 1506 281
rect -26 271 -22 272
rect -26 268 54 271
rect 106 268 230 271
rect 234 268 262 271
rect 274 268 326 271
rect 362 268 366 271
rect 402 268 406 271
rect 410 268 470 271
rect 474 268 494 271
rect 570 268 590 271
rect 618 268 654 271
rect 658 268 686 271
rect 758 268 766 271
rect 770 268 902 271
rect 914 268 942 271
rect 970 268 990 271
rect 994 268 1038 271
rect 1042 268 1062 271
rect 1074 268 1078 271
rect 1138 268 1150 271
rect 1226 268 1238 271
rect 70 258 86 261
rect 210 258 238 261
rect 426 258 438 261
rect 450 258 630 261
rect 634 258 742 261
rect 746 258 1014 261
rect 1034 258 1046 261
rect 1170 258 1177 261
rect 70 252 73 258
rect 206 252 209 258
rect 294 251 297 258
rect 218 248 297 251
rect 438 252 441 258
rect 1174 252 1177 258
rect 1214 261 1217 268
rect 1214 258 1222 261
rect 1278 261 1281 268
rect 1278 258 1286 261
rect 1354 258 1358 261
rect 1182 252 1185 258
rect 506 248 574 251
rect 650 248 702 251
rect 726 248 734 251
rect 738 248 782 251
rect 802 248 862 251
rect 882 248 910 251
rect 938 248 950 251
rect 970 248 974 251
rect 1098 248 1110 251
rect 1210 248 1214 251
rect 1226 248 1230 251
rect 1234 248 1246 251
rect 1306 248 1310 251
rect 1426 248 1446 251
rect 42 238 78 241
rect 98 238 126 241
rect 138 238 142 241
rect 202 238 230 241
rect 290 238 302 241
rect 314 238 550 241
rect 554 238 958 241
rect 982 241 985 248
rect 982 238 1038 241
rect 1110 238 1118 241
rect 1122 238 1142 241
rect 1170 238 1190 241
rect 1194 238 1254 241
rect 1258 238 1270 241
rect 1274 238 1350 241
rect 1354 238 1374 241
rect 1378 238 1414 241
rect 1418 238 1446 241
rect 42 228 502 231
rect 654 228 662 231
rect 666 228 694 231
rect 706 228 782 231
rect 794 228 806 231
rect 842 228 862 231
rect 874 228 902 231
rect 914 228 974 231
rect 1150 231 1153 238
rect 1150 228 1302 231
rect 1354 228 1358 231
rect 1378 228 1438 231
rect 82 218 118 221
rect 146 218 166 221
rect 258 218 318 221
rect 626 218 662 221
rect 666 218 1310 221
rect 1362 218 1366 221
rect 66 208 150 211
rect 170 208 182 211
rect 818 208 886 211
rect 898 208 1006 211
rect 1250 208 1302 211
rect 1354 208 1382 211
rect 472 203 474 207
rect 478 203 481 207
rect 486 203 488 207
rect 730 198 822 201
rect 826 198 846 201
rect 850 198 878 201
rect 890 198 1198 201
rect 1226 198 1286 201
rect 1330 198 1366 201
rect 1386 198 1446 201
rect 90 188 118 191
rect 122 188 206 191
rect 234 188 337 191
rect 678 188 686 191
rect 690 188 702 191
rect 842 188 894 191
rect 914 188 934 191
rect 1218 188 1230 191
rect 1294 188 1334 191
rect 334 182 337 188
rect 1294 182 1297 188
rect -26 178 38 181
rect 410 178 422 181
rect 466 178 662 181
rect 666 178 718 181
rect 770 178 774 181
rect 818 178 830 181
rect 962 178 1262 181
rect 1322 178 1422 181
rect -26 172 -23 178
rect -26 168 -22 172
rect 26 168 73 171
rect 238 171 241 178
rect 138 168 241 171
rect 702 168 886 171
rect 906 168 918 171
rect 1114 168 1150 171
rect 1170 168 1230 171
rect 1242 168 1270 171
rect 1298 168 1358 171
rect 1502 171 1506 172
rect 1482 168 1506 171
rect 70 162 73 168
rect 186 158 262 161
rect 362 158 630 161
rect 702 161 705 168
rect 634 158 705 161
rect 714 158 838 161
rect 890 158 1022 161
rect 1170 158 1222 161
rect 1226 158 1326 161
rect 1354 158 1390 161
rect -26 151 -22 152
rect 6 151 9 158
rect -26 148 14 151
rect 18 148 86 151
rect 270 151 273 158
rect 266 148 273 151
rect 330 148 414 151
rect 490 148 518 151
rect 626 148 758 151
rect 778 148 966 151
rect 1046 151 1049 158
rect 1034 148 1049 151
rect 1142 151 1145 158
rect 1142 148 1158 151
rect 1178 148 1182 151
rect 1202 148 1222 151
rect 1234 148 1270 151
rect 1326 148 1334 151
rect 1378 148 1406 151
rect 1502 148 1506 152
rect 198 142 201 148
rect 1326 142 1329 148
rect 54 138 78 141
rect 298 138 446 141
rect 450 138 454 141
rect 554 138 558 141
rect 646 138 710 141
rect 778 138 790 141
rect 806 138 830 141
rect 850 138 862 141
rect 922 138 945 141
rect 1074 138 1118 141
rect 1122 138 1129 141
rect 1210 138 1222 141
rect 1502 141 1505 148
rect 1370 138 1505 141
rect 54 132 57 138
rect 646 132 649 138
rect 162 128 230 131
rect 422 128 462 131
rect 538 128 614 131
rect 714 128 734 131
rect 758 131 761 138
rect 806 132 809 138
rect 942 132 945 138
rect 1342 132 1345 138
rect 758 128 774 131
rect 834 128 854 131
rect 1010 128 1062 131
rect 1218 128 1254 131
rect 1386 128 1390 131
rect 1502 131 1506 132
rect 1394 128 1506 131
rect 422 122 425 128
rect 90 118 206 121
rect 602 118 646 121
rect 650 118 1094 121
rect 1394 118 1406 121
rect 162 108 390 111
rect 394 108 574 111
rect 626 108 686 111
rect 810 108 822 111
rect 1330 108 1414 111
rect 1502 111 1506 112
rect 1482 108 1506 111
rect 114 98 166 101
rect 170 98 206 101
rect 210 98 262 101
rect 266 98 294 101
rect 298 98 318 101
rect 522 98 550 101
rect 622 101 625 108
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect 554 98 625 101
rect 658 98 958 101
rect 1010 98 1102 101
rect 1370 98 1382 101
rect 1386 98 1505 101
rect 1502 92 1505 98
rect -26 91 -22 92
rect -26 88 6 91
rect 10 88 38 91
rect 178 88 246 91
rect 346 88 526 91
rect 578 88 670 91
rect 786 88 830 91
rect 834 88 910 91
rect 930 88 966 91
rect 970 88 1017 91
rect 150 81 153 88
rect 1014 82 1017 88
rect 1098 88 1142 91
rect 1402 88 1406 91
rect 1502 88 1506 92
rect 98 78 153 81
rect 250 78 262 81
rect 338 78 358 81
rect 466 78 558 81
rect 562 78 574 81
rect 578 78 622 81
rect 698 78 742 81
rect 746 78 758 81
rect 958 78 1006 81
rect 1054 81 1057 88
rect 1034 78 1078 81
rect 1114 78 1158 81
rect 1182 81 1185 88
rect 1430 82 1433 88
rect 1162 78 1278 81
rect 1282 78 1302 81
rect 1378 78 1382 81
rect -26 71 -22 72
rect 46 71 49 78
rect -26 68 118 71
rect 282 68 318 71
rect 378 68 390 71
rect 394 68 438 71
rect 442 68 462 71
rect 466 68 542 71
rect 662 71 665 78
rect 662 68 814 71
rect 822 71 825 78
rect 958 72 961 78
rect 822 68 870 71
rect 874 68 910 71
rect 914 68 926 71
rect 1102 71 1105 78
rect 1082 68 1105 71
rect 1122 68 1190 71
rect 1234 68 1302 71
rect 1306 68 1310 71
rect 1426 68 1462 71
rect 1502 71 1506 72
rect 1466 68 1506 71
rect 1198 62 1201 68
rect 42 58 78 61
rect 202 58 398 61
rect 402 58 798 61
rect 802 58 966 61
rect 986 58 1022 61
rect 1106 58 1126 61
rect 1146 58 1158 61
rect 1162 58 1198 61
rect 1258 58 1265 61
rect 1262 52 1265 58
rect 82 48 102 51
rect 154 48 238 51
rect 258 48 278 51
rect 306 48 422 51
rect 426 48 486 51
rect 514 48 566 51
rect 602 48 662 51
rect 714 48 734 51
rect 866 48 902 51
rect 994 48 1166 51
rect 1194 48 1198 51
rect 1226 48 1238 51
rect 1290 48 1294 51
rect 1338 48 1358 51
rect 1502 51 1506 52
rect 1362 48 1506 51
rect 122 38 342 41
rect 346 38 622 41
rect 626 38 718 41
rect 794 38 1278 41
rect 1322 38 1334 41
rect 322 28 494 31
rect 542 28 550 31
rect 554 28 766 31
rect 890 28 894 31
rect 898 28 1062 31
rect 1166 28 1238 31
rect 1166 22 1169 28
rect 338 18 886 21
rect 906 18 918 21
rect 922 18 1078 21
rect 442 8 454 11
rect 730 8 750 11
rect 930 8 934 11
rect 962 8 966 11
rect 1074 8 1078 11
rect 472 3 474 7
rect 478 3 481 7
rect 486 3 488 7
<< m4contact >>
rect 350 1408 354 1412
rect 726 1408 730 1412
rect 886 1408 890 1412
rect 474 1403 478 1407
rect 482 1403 485 1407
rect 485 1403 486 1407
rect 278 1368 282 1372
rect 1262 1368 1266 1372
rect 110 1358 114 1362
rect 134 1358 138 1362
rect 918 1358 922 1362
rect 1166 1358 1170 1362
rect 1414 1358 1418 1362
rect 638 1348 642 1352
rect 78 1328 82 1332
rect 390 1328 394 1332
rect 614 1328 618 1332
rect 902 1328 906 1332
rect 1142 1328 1146 1332
rect 230 1318 234 1322
rect 270 1318 274 1322
rect 718 1318 722 1322
rect 974 1308 978 1312
rect 1454 1308 1458 1312
rect 986 1303 990 1307
rect 994 1303 997 1307
rect 997 1303 998 1307
rect 230 1298 234 1302
rect 638 1298 642 1302
rect 630 1278 634 1282
rect 638 1278 642 1282
rect 102 1268 106 1272
rect 126 1268 130 1272
rect 662 1258 666 1262
rect 1398 1258 1402 1262
rect 6 1248 10 1252
rect 534 1248 538 1252
rect 902 1248 906 1252
rect 910 1248 914 1252
rect 1254 1248 1258 1252
rect 1422 1248 1426 1252
rect 222 1238 226 1242
rect 474 1203 478 1207
rect 482 1203 485 1207
rect 485 1203 486 1207
rect 486 1188 490 1192
rect 622 1188 626 1192
rect 134 1178 138 1182
rect 126 1168 130 1172
rect 270 1168 274 1172
rect 878 1168 882 1172
rect 902 1168 906 1172
rect 1302 1168 1306 1172
rect 1430 1168 1434 1172
rect 294 1158 298 1162
rect 1366 1158 1370 1162
rect 46 1148 50 1152
rect 134 1148 138 1152
rect 718 1148 722 1152
rect 454 1138 458 1142
rect 614 1138 618 1142
rect 1430 1138 1434 1142
rect 1478 1138 1482 1142
rect 478 1128 482 1132
rect 502 1128 506 1132
rect 1006 1128 1010 1132
rect 1022 1128 1026 1132
rect 1326 1128 1330 1132
rect 574 1118 578 1122
rect 806 1118 810 1122
rect 870 1118 874 1122
rect 342 1108 346 1112
rect 986 1103 990 1107
rect 994 1103 997 1107
rect 997 1103 998 1107
rect 1006 1098 1010 1102
rect 382 1078 386 1082
rect 390 1078 394 1082
rect 750 1078 754 1082
rect 846 1078 850 1082
rect 1102 1078 1106 1082
rect 1406 1078 1410 1082
rect 486 1068 490 1072
rect 1182 1068 1186 1072
rect 1286 1068 1290 1072
rect 1310 1068 1314 1072
rect 254 1058 258 1062
rect 1374 1058 1378 1062
rect 1422 1058 1426 1062
rect 534 1048 538 1052
rect 878 1048 882 1052
rect 1478 1048 1482 1052
rect 646 1028 650 1032
rect 854 1018 858 1022
rect 582 1008 586 1012
rect 1046 1008 1050 1012
rect 1262 1008 1266 1012
rect 1334 1008 1338 1012
rect 1390 1008 1394 1012
rect 474 1003 478 1007
rect 482 1003 485 1007
rect 485 1003 486 1007
rect 462 998 466 1002
rect 654 998 658 1002
rect 1390 978 1394 982
rect 254 968 258 972
rect 462 968 466 972
rect 630 968 634 972
rect 1254 958 1258 962
rect 1334 958 1338 962
rect 1446 958 1450 962
rect 582 948 586 952
rect 1318 948 1322 952
rect 134 938 138 942
rect 558 938 562 942
rect 670 938 674 942
rect 1406 938 1410 942
rect 1294 928 1298 932
rect 1382 928 1386 932
rect 1086 918 1090 922
rect 1094 918 1098 922
rect 1358 918 1362 922
rect 1438 918 1442 922
rect 174 908 178 912
rect 534 908 538 912
rect 986 903 990 907
rect 994 903 997 907
rect 997 903 998 907
rect 1086 898 1090 902
rect 1438 898 1442 902
rect 326 868 330 872
rect 438 868 442 872
rect 598 868 602 872
rect 718 868 722 872
rect 790 868 794 872
rect 1198 868 1202 872
rect 142 858 146 862
rect 1046 858 1050 862
rect 1406 858 1410 862
rect 1318 848 1322 852
rect 1366 848 1370 852
rect 646 838 650 842
rect 750 838 754 842
rect 854 838 858 842
rect 870 838 874 842
rect 438 828 442 832
rect 494 808 498 812
rect 798 808 802 812
rect 1366 808 1370 812
rect 474 803 478 807
rect 482 803 485 807
rect 485 803 486 807
rect 622 798 626 802
rect 646 798 650 802
rect 654 798 658 802
rect 1302 798 1306 802
rect 1478 798 1482 802
rect 78 788 82 792
rect 462 788 466 792
rect 1030 788 1034 792
rect 726 778 730 782
rect 798 778 802 782
rect 870 778 874 782
rect 1390 778 1394 782
rect 494 768 498 772
rect 790 768 794 772
rect 814 768 818 772
rect 1286 768 1290 772
rect 798 758 802 762
rect 878 758 882 762
rect 1030 758 1034 762
rect 1374 758 1378 762
rect 342 748 346 752
rect 1086 748 1090 752
rect 166 738 170 742
rect 606 738 610 742
rect 670 738 674 742
rect 694 738 698 742
rect 702 738 706 742
rect 766 738 770 742
rect 1382 738 1386 742
rect 734 728 738 732
rect 1358 728 1362 732
rect 686 698 690 702
rect 986 703 990 707
rect 994 703 997 707
rect 997 703 998 707
rect 6 688 10 692
rect 342 688 346 692
rect 1318 688 1322 692
rect 654 678 658 682
rect 758 678 762 682
rect 1262 678 1266 682
rect 6 668 10 672
rect 342 668 346 672
rect 566 668 570 672
rect 598 668 602 672
rect 702 668 706 672
rect 718 668 722 672
rect 750 668 754 672
rect 814 668 818 672
rect 854 668 858 672
rect 1270 668 1274 672
rect 1302 668 1306 672
rect 1478 668 1482 672
rect 78 658 82 662
rect 638 658 642 662
rect 758 658 762 662
rect 1246 658 1250 662
rect 366 648 370 652
rect 686 648 690 652
rect 694 648 698 652
rect 670 638 674 642
rect 230 628 234 632
rect 382 628 386 632
rect 494 628 498 632
rect 550 628 554 632
rect 798 628 802 632
rect 366 608 370 612
rect 474 603 478 607
rect 482 603 485 607
rect 485 603 486 607
rect 158 578 162 582
rect 342 578 346 582
rect 126 568 130 572
rect 510 568 514 572
rect 1278 568 1282 572
rect 54 558 58 562
rect 78 558 82 562
rect 110 558 114 562
rect 174 558 178 562
rect 334 558 338 562
rect 38 548 42 552
rect 206 548 210 552
rect 382 548 386 552
rect 774 548 778 552
rect 1318 548 1322 552
rect 6 538 10 542
rect 54 538 58 542
rect 126 538 130 542
rect 150 538 154 542
rect 166 538 170 542
rect 366 538 370 542
rect 454 538 458 542
rect 1054 538 1058 542
rect 1270 538 1274 542
rect 1342 538 1346 542
rect 46 528 50 532
rect 134 528 138 532
rect 230 528 234 532
rect 286 528 290 532
rect 566 528 570 532
rect 662 528 666 532
rect 62 518 66 522
rect 1054 518 1058 522
rect 986 503 990 507
rect 994 503 997 507
rect 997 503 998 507
rect 430 498 434 502
rect 278 488 282 492
rect 558 488 562 492
rect 622 488 626 492
rect 1246 488 1250 492
rect 462 478 466 482
rect 742 478 746 482
rect 774 478 778 482
rect 342 468 346 472
rect 358 468 362 472
rect 662 468 666 472
rect 758 468 762 472
rect 782 468 786 472
rect 790 458 794 462
rect 1110 468 1114 472
rect 1230 468 1234 472
rect 1102 458 1106 462
rect 358 448 362 452
rect 422 448 426 452
rect 598 448 602 452
rect 150 438 154 442
rect 1294 438 1298 442
rect 510 428 514 432
rect 574 428 578 432
rect 46 408 50 412
rect 502 408 506 412
rect 702 408 706 412
rect 474 403 478 407
rect 482 403 485 407
rect 485 403 486 407
rect 494 398 498 402
rect 766 398 770 402
rect 934 398 938 402
rect 1318 388 1322 392
rect 598 378 602 382
rect 134 368 138 372
rect 334 368 338 372
rect 774 358 778 362
rect 1254 358 1258 362
rect 1278 358 1282 362
rect 1454 358 1458 362
rect 1478 358 1482 362
rect 454 348 458 352
rect 814 348 818 352
rect 838 348 842 352
rect 1166 348 1170 352
rect 1238 348 1242 352
rect 1246 348 1250 352
rect 1334 348 1338 352
rect 1350 348 1354 352
rect 110 338 114 342
rect 278 338 282 342
rect 566 338 570 342
rect 790 338 794 342
rect 910 338 914 342
rect 1198 338 1202 342
rect 462 328 466 332
rect 550 328 554 332
rect 1070 328 1074 332
rect 1246 328 1250 332
rect 1478 328 1482 332
rect 1014 308 1018 312
rect 986 303 990 307
rect 994 303 997 307
rect 997 303 998 307
rect 1006 298 1010 302
rect 654 288 658 292
rect 446 278 450 282
rect 766 278 770 282
rect 1014 278 1018 282
rect 358 268 362 272
rect 1070 268 1074 272
rect 438 258 442 262
rect 1014 258 1018 262
rect 1030 258 1034 262
rect 1166 258 1170 262
rect 206 248 210 252
rect 1350 258 1354 262
rect 574 248 578 252
rect 782 248 786 252
rect 910 248 914 252
rect 966 248 970 252
rect 1182 248 1186 252
rect 1206 248 1210 252
rect 1222 248 1226 252
rect 1310 248 1314 252
rect 134 238 138 242
rect 502 228 506 232
rect 910 228 914 232
rect 1350 228 1354 232
rect 1438 228 1442 232
rect 662 218 666 222
rect 1358 218 1362 222
rect 1302 208 1306 212
rect 474 203 478 207
rect 482 203 485 207
rect 485 203 486 207
rect 886 198 890 202
rect 1286 198 1290 202
rect 1326 198 1330 202
rect 1446 198 1450 202
rect 206 188 210 192
rect 422 178 426 182
rect 462 178 466 182
rect 766 178 770 182
rect 958 178 962 182
rect 1422 178 1426 182
rect 886 168 890 172
rect 1230 168 1234 172
rect 1358 168 1362 172
rect 1222 158 1226 162
rect 758 148 762 152
rect 1174 148 1178 152
rect 1230 148 1234 152
rect 1374 148 1378 152
rect 198 138 202 142
rect 454 138 458 142
rect 550 138 554 142
rect 774 138 778 142
rect 1070 138 1074 142
rect 1342 138 1346 142
rect 614 128 618 132
rect 1390 128 1394 132
rect 1406 118 1410 122
rect 1414 108 1418 112
rect 986 103 990 107
rect 994 103 997 107
rect 997 103 998 107
rect 654 98 658 102
rect 1366 98 1370 102
rect 38 88 42 92
rect 1398 88 1402 92
rect 1430 88 1434 92
rect 262 78 266 82
rect 1030 78 1034 82
rect 1382 78 1386 82
rect 814 68 818 72
rect 1190 68 1194 72
rect 1310 68 1314 72
rect 1462 68 1466 72
rect 1198 58 1202 62
rect 486 48 490 52
rect 1190 48 1194 52
rect 1222 48 1226 52
rect 1294 48 1298 52
rect 1334 48 1338 52
rect 1318 38 1322 42
rect 902 18 906 22
rect 438 8 442 12
rect 926 8 930 12
rect 966 8 970 12
rect 1078 8 1082 12
rect 474 3 478 7
rect 482 3 485 7
rect 485 3 486 7
<< metal4 >>
rect 342 1408 350 1411
rect 718 1408 726 1411
rect 878 1408 886 1411
rect 278 1362 281 1368
rect 138 1358 142 1361
rect 110 1352 113 1358
rect 6 1252 9 1268
rect 50 1148 54 1151
rect 78 1112 81 1328
rect 230 1302 233 1318
rect 106 1268 110 1271
rect 126 1172 129 1268
rect 222 1242 225 1268
rect 134 1152 137 1178
rect 270 1172 273 1318
rect 294 1152 297 1158
rect 342 1112 345 1408
rect 472 1403 474 1407
rect 478 1403 481 1407
rect 486 1403 488 1407
rect 634 1348 638 1351
rect 394 1328 398 1331
rect 472 1203 474 1207
rect 478 1203 481 1207
rect 486 1203 488 1207
rect 458 1138 462 1141
rect 478 1122 481 1128
rect 382 1082 385 1088
rect 390 1062 393 1078
rect 486 1072 489 1188
rect 494 1128 502 1131
rect 494 1112 497 1128
rect 490 1068 494 1071
rect 254 972 257 1058
rect 534 1052 537 1248
rect 614 1142 617 1328
rect 718 1322 721 1408
rect 638 1282 641 1298
rect 630 1191 633 1278
rect 662 1252 665 1258
rect 626 1188 633 1191
rect 878 1172 881 1408
rect 1258 1368 1262 1371
rect 1166 1362 1169 1368
rect 918 1352 921 1358
rect 898 1328 902 1331
rect 1138 1328 1142 1331
rect 974 1312 977 1328
rect 984 1303 986 1307
rect 990 1303 993 1307
rect 998 1303 1000 1307
rect 914 1248 918 1251
rect 902 1172 905 1248
rect 718 1142 721 1148
rect 1010 1128 1017 1131
rect 1014 1122 1017 1128
rect 578 1118 582 1121
rect 750 1082 753 1088
rect 472 1003 474 1007
rect 478 1003 481 1007
rect 486 1003 488 1007
rect 462 972 465 998
rect 6 672 9 688
rect 78 662 81 788
rect 82 558 86 561
rect 38 552 41 558
rect 54 552 57 558
rect 54 542 57 548
rect 10 538 14 541
rect 46 412 49 528
rect 62 522 65 538
rect 110 342 113 558
rect 126 542 129 568
rect 134 532 137 938
rect 534 912 537 1048
rect 582 952 585 1008
rect 562 938 566 941
rect 142 441 145 858
rect 158 541 161 578
rect 154 538 161 541
rect 166 542 169 738
rect 174 562 177 908
rect 330 868 334 871
rect 438 832 441 868
rect 472 803 474 807
rect 478 803 481 807
rect 486 803 488 807
rect 458 788 462 791
rect 494 772 497 808
rect 342 692 345 748
rect 598 672 601 868
rect 630 801 633 968
rect 646 842 649 1028
rect 654 802 657 998
rect 666 938 670 941
rect 794 868 798 871
rect 626 798 633 801
rect 606 682 609 738
rect 646 692 649 798
rect 674 738 678 741
rect 706 738 710 741
rect 654 672 657 678
rect 558 668 566 671
rect 142 438 150 441
rect 38 92 41 328
rect 134 242 137 368
rect 206 252 209 548
rect 230 532 233 628
rect 342 582 345 668
rect 358 648 366 651
rect 234 528 238 531
rect 278 528 286 531
rect 278 512 281 528
rect 278 492 281 508
rect 334 372 337 558
rect 342 472 345 578
rect 358 472 361 648
rect 382 632 385 638
rect 550 632 553 648
rect 366 542 369 608
rect 472 603 474 607
rect 478 603 481 607
rect 486 603 488 607
rect 378 548 382 551
rect 458 538 465 541
rect 366 482 369 538
rect 282 338 286 341
rect 358 272 361 448
rect 206 192 209 248
rect 422 182 425 448
rect 430 322 433 498
rect 462 482 465 538
rect 472 403 474 407
rect 478 403 481 407
rect 486 403 488 407
rect 494 402 497 628
rect 510 432 513 568
rect 558 492 561 668
rect 638 652 641 658
rect 686 652 689 698
rect 694 652 697 738
rect 702 672 705 678
rect 718 672 721 868
rect 750 792 753 838
rect 798 782 801 808
rect 726 731 729 778
rect 806 771 809 1118
rect 870 1112 873 1118
rect 984 1103 986 1107
rect 990 1103 993 1107
rect 998 1103 1000 1107
rect 850 1078 854 1081
rect 1006 1072 1009 1098
rect 1022 1092 1025 1128
rect 1098 1078 1102 1081
rect 1178 1068 1182 1071
rect 854 842 857 1018
rect 870 782 873 838
rect 806 768 814 771
rect 790 752 793 768
rect 878 762 881 1048
rect 1254 1011 1257 1248
rect 1302 1071 1305 1168
rect 1302 1068 1310 1071
rect 1254 1008 1262 1011
rect 984 903 986 907
rect 990 903 993 907
rect 998 903 1000 907
rect 1046 862 1049 1008
rect 1086 902 1089 918
rect 1030 762 1033 788
rect 726 728 734 731
rect 750 672 753 688
rect 758 662 761 678
rect 666 638 670 641
rect 658 528 662 531
rect 454 281 457 348
rect 450 278 457 281
rect 198 132 201 138
rect 262 82 265 88
rect 438 12 441 258
rect 462 182 465 328
rect 502 232 505 408
rect 566 342 569 528
rect 622 492 625 508
rect 742 472 745 478
rect 758 472 761 478
rect 546 328 550 331
rect 574 252 577 428
rect 598 382 601 448
rect 662 342 665 468
rect 702 342 705 408
rect 766 402 769 738
rect 798 632 801 758
rect 1082 748 1086 751
rect 984 703 986 707
rect 990 703 993 707
rect 998 703 1000 707
rect 850 668 854 671
rect 774 482 777 548
rect 778 468 782 471
rect 778 358 782 361
rect 790 342 793 458
rect 814 352 817 668
rect 1054 522 1057 538
rect 984 503 986 507
rect 990 503 993 507
rect 998 503 1000 507
rect 842 348 846 351
rect 910 342 913 348
rect 472 203 474 207
rect 478 203 481 207
rect 486 203 488 207
rect 450 138 454 141
rect 550 132 553 138
rect 614 82 617 128
rect 654 102 657 288
rect 662 222 665 338
rect 766 182 769 278
rect 786 248 790 251
rect 910 232 913 248
rect 886 172 889 198
rect 762 148 766 151
rect 770 138 774 141
rect 654 92 657 98
rect 814 52 817 68
rect 486 22 489 48
rect 898 18 902 21
rect 934 11 937 398
rect 1070 332 1073 338
rect 984 303 986 307
rect 990 303 993 307
rect 998 303 1000 307
rect 1006 302 1009 318
rect 1014 312 1017 328
rect 1014 262 1017 278
rect 1070 272 1073 328
rect 1026 258 1030 261
rect 974 251 977 258
rect 970 248 977 251
rect 930 8 937 11
rect 958 11 961 178
rect 1070 132 1073 138
rect 1094 132 1097 918
rect 1194 868 1198 871
rect 1254 661 1257 958
rect 1286 772 1289 1068
rect 1262 672 1265 678
rect 1294 671 1297 928
rect 1318 852 1321 948
rect 1302 792 1305 798
rect 1294 668 1302 671
rect 1250 658 1257 661
rect 1270 542 1273 668
rect 1282 568 1289 571
rect 1110 472 1113 478
rect 1234 468 1238 471
rect 1102 462 1105 468
rect 1246 352 1249 488
rect 1274 358 1278 361
rect 1254 352 1257 358
rect 1170 348 1174 351
rect 1238 342 1241 348
rect 1170 258 1174 261
rect 1178 248 1182 251
rect 1178 148 1182 151
rect 984 103 986 107
rect 990 103 993 107
rect 998 103 1000 107
rect 1026 78 1030 81
rect 958 8 966 11
rect 1070 11 1073 128
rect 1190 52 1193 68
rect 1198 62 1201 338
rect 1246 332 1249 348
rect 1214 251 1217 258
rect 1210 248 1217 251
rect 1222 162 1225 248
rect 1286 202 1289 568
rect 1318 552 1321 688
rect 1298 438 1305 441
rect 1302 212 1305 438
rect 1222 52 1225 158
rect 1230 152 1233 168
rect 1310 72 1313 248
rect 1290 48 1294 51
rect 1318 42 1321 388
rect 1326 202 1329 1128
rect 1334 962 1337 1008
rect 1358 732 1361 918
rect 1366 852 1369 1158
rect 1334 52 1337 348
rect 1342 142 1345 538
rect 1354 348 1361 351
rect 1358 342 1361 348
rect 1350 232 1353 258
rect 1358 172 1361 218
rect 1366 102 1369 808
rect 1374 762 1377 1058
rect 1390 982 1393 1008
rect 1386 928 1393 931
rect 1390 782 1393 928
rect 1374 152 1377 758
rect 1382 82 1385 738
rect 1390 132 1393 138
rect 1398 92 1401 1258
rect 1406 942 1409 1078
rect 1414 892 1417 1358
rect 1422 1062 1425 1248
rect 1434 1168 1441 1171
rect 1406 122 1409 858
rect 1414 112 1417 818
rect 1422 182 1425 1048
rect 1430 92 1433 1138
rect 1438 1052 1441 1168
rect 1438 902 1441 918
rect 1438 232 1441 888
rect 1446 202 1449 958
rect 1454 362 1457 1308
rect 1462 72 1465 1248
rect 1478 1122 1481 1138
rect 1478 1052 1481 1068
rect 1478 822 1481 1048
rect 1474 798 1478 801
rect 1474 668 1478 671
rect 1478 332 1481 358
rect 1070 8 1078 11
rect 472 3 474 7
rect 478 3 481 7
rect 486 3 488 7
<< m5contact >>
rect 142 1358 146 1362
rect 278 1358 282 1362
rect 110 1348 114 1352
rect 6 1268 10 1272
rect 54 1148 58 1152
rect 110 1268 114 1272
rect 222 1268 226 1272
rect 294 1148 298 1152
rect 474 1403 478 1407
rect 481 1403 482 1407
rect 482 1403 485 1407
rect 630 1348 634 1352
rect 398 1328 402 1332
rect 474 1203 478 1207
rect 481 1203 482 1207
rect 482 1203 485 1207
rect 462 1138 466 1142
rect 478 1118 482 1122
rect 78 1108 82 1112
rect 382 1088 386 1092
rect 494 1108 498 1112
rect 494 1068 498 1072
rect 390 1058 394 1062
rect 662 1248 666 1252
rect 1166 1368 1170 1372
rect 1254 1368 1258 1372
rect 918 1348 922 1352
rect 894 1328 898 1332
rect 974 1328 978 1332
rect 1134 1328 1138 1332
rect 986 1303 990 1307
rect 993 1303 994 1307
rect 994 1303 997 1307
rect 918 1248 922 1252
rect 718 1138 722 1142
rect 582 1118 586 1122
rect 1014 1118 1018 1122
rect 750 1088 754 1092
rect 474 1003 478 1007
rect 481 1003 482 1007
rect 482 1003 485 1007
rect 38 558 42 562
rect 86 558 90 562
rect 54 548 58 552
rect 14 538 18 542
rect 62 538 66 542
rect 566 938 570 942
rect 334 868 338 872
rect 474 803 478 807
rect 481 803 482 807
rect 482 803 485 807
rect 454 788 458 792
rect 662 938 666 942
rect 798 868 802 872
rect 678 738 682 742
rect 710 738 714 742
rect 646 688 650 692
rect 606 678 610 682
rect 654 668 658 672
rect 38 328 42 332
rect 550 648 554 652
rect 238 528 242 532
rect 278 508 282 512
rect 382 638 386 642
rect 474 603 478 607
rect 481 603 482 607
rect 482 603 485 607
rect 374 548 378 552
rect 366 478 370 482
rect 286 338 290 342
rect 474 403 478 407
rect 481 403 482 407
rect 482 403 485 407
rect 702 678 706 682
rect 750 788 754 792
rect 870 1108 874 1112
rect 986 1103 990 1107
rect 993 1103 994 1107
rect 994 1103 997 1107
rect 854 1078 858 1082
rect 1022 1088 1026 1092
rect 1094 1078 1098 1082
rect 1006 1068 1010 1072
rect 1174 1068 1178 1072
rect 986 903 990 907
rect 993 903 994 907
rect 994 903 997 907
rect 790 748 794 752
rect 750 688 754 692
rect 638 648 642 652
rect 662 638 666 642
rect 654 528 658 532
rect 430 318 434 322
rect 198 128 202 132
rect 262 88 266 92
rect 622 508 626 512
rect 758 478 762 482
rect 742 468 746 472
rect 542 328 546 332
rect 1078 748 1082 752
rect 986 703 990 707
rect 993 703 994 707
rect 994 703 997 707
rect 846 668 850 672
rect 774 468 778 472
rect 782 358 786 362
rect 986 503 990 507
rect 993 503 994 507
rect 994 503 997 507
rect 846 348 850 352
rect 910 348 914 352
rect 662 338 666 342
rect 702 338 706 342
rect 474 203 478 207
rect 481 203 482 207
rect 482 203 485 207
rect 446 138 450 142
rect 550 128 554 132
rect 790 248 794 252
rect 766 148 770 152
rect 766 138 770 142
rect 654 88 658 92
rect 614 78 618 82
rect 814 48 818 52
rect 486 18 490 22
rect 894 18 898 22
rect 1070 338 1074 342
rect 1014 328 1018 332
rect 1006 318 1010 322
rect 986 303 990 307
rect 993 303 994 307
rect 994 303 997 307
rect 974 258 978 262
rect 1022 258 1026 262
rect 1190 868 1194 872
rect 1262 668 1266 672
rect 1302 788 1306 792
rect 1110 478 1114 482
rect 1102 468 1106 472
rect 1238 468 1242 472
rect 1270 358 1274 362
rect 1174 348 1178 352
rect 1254 348 1258 352
rect 1238 338 1242 342
rect 1174 258 1178 262
rect 1174 248 1178 252
rect 1182 148 1186 152
rect 1070 128 1074 132
rect 1094 128 1098 132
rect 986 103 990 107
rect 993 103 994 107
rect 994 103 997 107
rect 1022 78 1026 82
rect 1214 258 1218 262
rect 1286 48 1290 52
rect 1358 338 1362 342
rect 1390 138 1394 142
rect 1422 1048 1426 1052
rect 1414 888 1418 892
rect 1414 818 1418 822
rect 1438 1048 1442 1052
rect 1438 888 1442 892
rect 1462 1248 1466 1252
rect 1478 1118 1482 1122
rect 1478 1068 1482 1072
rect 1478 818 1482 822
rect 1470 798 1474 802
rect 1470 668 1474 672
rect 474 3 478 7
rect 481 3 482 7
rect 482 3 485 7
<< metal5 >>
rect 478 1403 481 1407
rect 478 1402 482 1403
rect 1170 1368 1254 1371
rect 146 1358 278 1361
rect 114 1348 630 1351
rect 634 1348 918 1351
rect 402 1328 894 1331
rect 978 1328 1134 1331
rect 990 1303 993 1307
rect 990 1302 994 1303
rect 10 1268 110 1271
rect 114 1268 222 1271
rect 666 1248 918 1251
rect 922 1248 1462 1251
rect 478 1203 481 1207
rect 478 1202 482 1203
rect 58 1148 294 1151
rect 466 1138 718 1141
rect 482 1118 582 1121
rect 586 1118 1014 1121
rect 1018 1118 1478 1121
rect 82 1108 494 1111
rect 498 1108 870 1111
rect 990 1103 993 1107
rect 990 1102 994 1103
rect 386 1088 750 1091
rect 754 1088 1022 1091
rect 858 1078 1094 1081
rect 498 1068 1006 1071
rect 1178 1068 1478 1071
rect 1174 1061 1177 1068
rect 394 1058 1177 1061
rect 1426 1048 1438 1051
rect 478 1003 481 1007
rect 478 1002 482 1003
rect 570 938 662 941
rect 990 903 993 907
rect 990 902 994 903
rect 1418 888 1438 891
rect 338 868 798 871
rect 802 868 1190 871
rect 1418 818 1478 821
rect 478 803 481 807
rect 478 802 482 803
rect 1302 798 1470 801
rect 1302 792 1305 798
rect 458 788 750 791
rect 794 748 1078 751
rect 682 738 710 741
rect 990 703 993 707
rect 990 702 994 703
rect 650 688 750 691
rect 610 678 702 681
rect 658 668 846 671
rect 1266 668 1470 671
rect 554 648 638 651
rect 386 638 662 641
rect 478 603 481 607
rect 478 602 482 603
rect 42 558 86 561
rect 58 548 374 551
rect 18 538 62 541
rect 242 528 654 531
rect 282 508 622 511
rect 990 503 993 507
rect 990 502 994 503
rect 370 478 758 481
rect 762 478 1110 481
rect 746 468 774 471
rect 1106 468 1238 471
rect 478 403 481 407
rect 478 402 482 403
rect 786 358 1270 361
rect 850 348 910 351
rect 1178 348 1254 351
rect 290 338 662 341
rect 706 338 1070 341
rect 1242 338 1358 341
rect 42 328 542 331
rect 546 328 1014 331
rect 434 318 1006 321
rect 990 303 993 307
rect 990 302 994 303
rect 978 258 1022 261
rect 1178 258 1214 261
rect 794 248 1174 251
rect 478 203 481 207
rect 478 202 482 203
rect 770 148 1182 151
rect 450 138 766 141
rect 202 128 550 131
rect 554 128 1070 131
rect 1390 131 1393 138
rect 1098 128 1393 131
rect 990 103 993 107
rect 990 102 994 103
rect 266 88 654 91
rect 618 78 1022 81
rect 818 48 1286 51
rect 490 18 894 21
rect 478 3 481 7
rect 478 2 482 3
<< m6contact >>
rect 472 1407 478 1408
rect 482 1407 488 1408
rect 472 1403 474 1407
rect 474 1403 478 1407
rect 482 1403 485 1407
rect 485 1403 488 1407
rect 472 1402 478 1403
rect 482 1402 488 1403
rect 984 1307 990 1308
rect 994 1307 1000 1308
rect 984 1303 986 1307
rect 986 1303 990 1307
rect 994 1303 997 1307
rect 997 1303 1000 1307
rect 984 1302 990 1303
rect 994 1302 1000 1303
rect 472 1207 478 1208
rect 482 1207 488 1208
rect 472 1203 474 1207
rect 474 1203 478 1207
rect 482 1203 485 1207
rect 485 1203 488 1207
rect 472 1202 478 1203
rect 482 1202 488 1203
rect 984 1107 990 1108
rect 994 1107 1000 1108
rect 984 1103 986 1107
rect 986 1103 990 1107
rect 994 1103 997 1107
rect 997 1103 1000 1107
rect 984 1102 990 1103
rect 994 1102 1000 1103
rect 472 1007 478 1008
rect 482 1007 488 1008
rect 472 1003 474 1007
rect 474 1003 478 1007
rect 482 1003 485 1007
rect 485 1003 488 1007
rect 472 1002 478 1003
rect 482 1002 488 1003
rect 984 907 990 908
rect 994 907 1000 908
rect 984 903 986 907
rect 986 903 990 907
rect 994 903 997 907
rect 997 903 1000 907
rect 984 902 990 903
rect 994 902 1000 903
rect 472 807 478 808
rect 482 807 488 808
rect 472 803 474 807
rect 474 803 478 807
rect 482 803 485 807
rect 485 803 488 807
rect 472 802 478 803
rect 482 802 488 803
rect 984 707 990 708
rect 994 707 1000 708
rect 984 703 986 707
rect 986 703 990 707
rect 994 703 997 707
rect 997 703 1000 707
rect 984 702 990 703
rect 994 702 1000 703
rect 472 607 478 608
rect 482 607 488 608
rect 472 603 474 607
rect 474 603 478 607
rect 482 603 485 607
rect 485 603 488 607
rect 472 602 478 603
rect 482 602 488 603
rect 984 507 990 508
rect 994 507 1000 508
rect 984 503 986 507
rect 986 503 990 507
rect 994 503 997 507
rect 997 503 1000 507
rect 984 502 990 503
rect 994 502 1000 503
rect 472 407 478 408
rect 482 407 488 408
rect 472 403 474 407
rect 474 403 478 407
rect 482 403 485 407
rect 485 403 488 407
rect 472 402 478 403
rect 482 402 488 403
rect 984 307 990 308
rect 994 307 1000 308
rect 984 303 986 307
rect 986 303 990 307
rect 994 303 997 307
rect 997 303 1000 307
rect 984 302 990 303
rect 994 302 1000 303
rect 472 207 478 208
rect 482 207 488 208
rect 472 203 474 207
rect 474 203 478 207
rect 482 203 485 207
rect 485 203 488 207
rect 472 202 478 203
rect 482 202 488 203
rect 984 107 990 108
rect 994 107 1000 108
rect 984 103 986 107
rect 986 103 990 107
rect 994 103 997 107
rect 997 103 1000 107
rect 984 102 990 103
rect 994 102 1000 103
rect 472 7 478 8
rect 482 7 488 8
rect 472 3 474 7
rect 474 3 478 7
rect 482 3 485 7
rect 485 3 488 7
rect 472 2 478 3
rect 482 2 488 3
<< metal6 >>
rect 472 1408 488 1440
rect 478 1402 482 1408
rect 472 1208 488 1402
rect 478 1202 482 1208
rect 472 1008 488 1202
rect 478 1002 482 1008
rect 472 808 488 1002
rect 478 802 482 808
rect 472 608 488 802
rect 478 602 482 608
rect 472 408 488 602
rect 478 402 482 408
rect 472 208 488 402
rect 478 202 482 208
rect 472 8 488 202
rect 478 2 482 8
rect 472 -30 488 2
rect 984 1308 1000 1440
rect 990 1302 994 1308
rect 984 1108 1000 1302
rect 990 1102 994 1108
rect 984 908 1000 1102
rect 990 902 994 908
rect 984 708 1000 902
rect 990 702 994 708
rect 984 508 1000 702
rect 990 502 994 508
rect 984 308 1000 502
rect 990 302 994 308
rect 984 108 1000 302
rect 990 102 994 108
rect 984 -30 1000 102
use INVX1  _1287_
timestamp 1559787497
transform 1 0 4 0 1 1305
box -2 -3 18 103
use OAI21X1  _1289_
timestamp 1559787497
transform 1 0 20 0 1 1305
box -2 -3 34 103
use NAND2X1  _1276_
timestamp 1559787497
transform 1 0 52 0 1 1305
box -2 -3 26 103
use INVX1  _1275_
timestamp 1559787497
transform 1 0 76 0 1 1305
box -2 -3 18 103
use NAND2X1  _1288_
timestamp 1559787497
transform 1 0 92 0 1 1305
box -2 -3 26 103
use NAND2X1  _1251_
timestamp 1559787497
transform 1 0 116 0 1 1305
box -2 -3 26 103
use NAND2X1  _1207_
timestamp 1559787497
transform 1 0 140 0 1 1305
box -2 -3 26 103
use INVX1  _1206_
timestamp 1559787497
transform -1 0 180 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_insert38
timestamp 1559787497
transform -1 0 204 0 1 1305
box -2 -3 26 103
use NAND2X1  _1212_
timestamp 1559787497
transform -1 0 228 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert37
timestamp 1559787497
transform 1 0 228 0 1 1305
box -2 -3 26 103
use NAND2X1  _1171_
timestamp 1559787497
transform 1 0 252 0 1 1305
box -2 -3 26 103
use OAI21X1  _1211_
timestamp 1559787497
transform -1 0 308 0 1 1305
box -2 -3 34 103
use INVX1  _1209_
timestamp 1559787497
transform 1 0 308 0 1 1305
box -2 -3 18 103
use NAND2X1  _1210_
timestamp 1559787497
transform 1 0 324 0 1 1305
box -2 -3 26 103
use OAI21X1  _1250_
timestamp 1559787497
transform 1 0 348 0 1 1305
box -2 -3 34 103
use INVX1  _1248_
timestamp 1559787497
transform -1 0 396 0 1 1305
box -2 -3 18 103
use NAND2X1  _1249_
timestamp 1559787497
transform 1 0 396 0 1 1305
box -2 -3 26 103
use NAND2X1  _917_
timestamp 1559787497
transform -1 0 444 0 1 1305
box -2 -3 26 103
use OAI21X1  _1170_
timestamp 1559787497
transform -1 0 476 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1559787497
transform 1 0 476 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1559787497
transform 1 0 484 0 1 1305
box -2 -3 10 103
use NAND2X1  _1169_
timestamp 1559787497
transform 1 0 492 0 1 1305
box -2 -3 26 103
use INVX1  _1168_
timestamp 1559787497
transform -1 0 532 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_insert11
timestamp 1559787497
transform -1 0 556 0 1 1305
box -2 -3 26 103
use INVX1  _955_
timestamp 1559787497
transform 1 0 556 0 1 1305
box -2 -3 18 103
use OAI21X1  _957_
timestamp 1559787497
transform 1 0 572 0 1 1305
box -2 -3 34 103
use NAND2X1  _958_
timestamp 1559787497
transform -1 0 628 0 1 1305
box -2 -3 26 103
use NAND2X1  _956_
timestamp 1559787497
transform -1 0 652 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert12
timestamp 1559787497
transform 1 0 652 0 1 1305
box -2 -3 26 103
use NAND2X1  _878_
timestamp 1559787497
transform 1 0 676 0 1 1305
box -2 -3 26 103
use NAND2X1  _837_
timestamp 1559787497
transform 1 0 700 0 1 1305
box -2 -3 26 103
use INVX1  _670_
timestamp 1559787497
transform 1 0 724 0 1 1305
box -2 -3 18 103
use OAI21X1  _672_
timestamp 1559787497
transform 1 0 740 0 1 1305
box -2 -3 34 103
use NAND2X1  _671_
timestamp 1559787497
transform -1 0 796 0 1 1305
box -2 -3 26 103
use NAND2X1  _712_
timestamp 1559787497
transform -1 0 820 0 1 1305
box -2 -3 26 103
use NAND2X1  _673_
timestamp 1559787497
transform -1 0 844 0 1 1305
box -2 -3 26 103
use INVX1  _747_
timestamp 1559787497
transform 1 0 844 0 1 1305
box -2 -3 18 103
use NAND2X1  _748_
timestamp 1559787497
transform -1 0 884 0 1 1305
box -2 -3 26 103
use NAND2X1  _753_
timestamp 1559787497
transform 1 0 884 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert20
timestamp 1559787497
transform -1 0 932 0 1 1305
box -2 -3 26 103
use INVX1  _750_
timestamp 1559787497
transform 1 0 932 0 1 1305
box -2 -3 18 103
use OAI21X1  _752_
timestamp 1559787497
transform 1 0 948 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1559787497
transform -1 0 988 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1559787497
transform -1 0 996 0 1 1305
box -2 -3 10 103
use NAND2X1  _751_
timestamp 1559787497
transform -1 0 1020 0 1 1305
box -2 -3 26 103
use NAND2X1  _790_
timestamp 1559787497
transform 1 0 1020 0 1 1305
box -2 -3 26 103
use INVX1  _1082_
timestamp 1559787497
transform 1 0 1044 0 1 1305
box -2 -3 18 103
use NAND2X1  _1083_
timestamp 1559787497
transform -1 0 1084 0 1 1305
box -2 -3 26 103
use OAI21X1  _1084_
timestamp 1559787497
transform 1 0 1084 0 1 1305
box -2 -3 34 103
use NAND2X1  _1122_
timestamp 1559787497
transform -1 0 1140 0 1 1305
box -2 -3 26 103
use OAI21X1  _1123_
timestamp 1559787497
transform -1 0 1172 0 1 1305
box -2 -3 34 103
use NAND2X1  _1044_
timestamp 1559787497
transform -1 0 1196 0 1 1305
box -2 -3 26 103
use OAI21X1  _1045_
timestamp 1559787497
transform 1 0 1196 0 1 1305
box -2 -3 34 103
use INVX1  _1040_
timestamp 1559787497
transform 1 0 1228 0 1 1305
box -2 -3 18 103
use NAND2X1  _1041_
timestamp 1559787497
transform -1 0 1268 0 1 1305
box -2 -3 26 103
use NAND2X1  _1085_
timestamp 1559787497
transform -1 0 1292 0 1 1305
box -2 -3 26 103
use NAND2X1  _1124_
timestamp 1559787497
transform -1 0 1316 0 1 1305
box -2 -3 26 103
use NAND2X1  _1046_
timestamp 1559787497
transform -1 0 1340 0 1 1305
box -2 -3 26 103
use INVX1  _1002_
timestamp 1559787497
transform 1 0 1340 0 1 1305
box -2 -3 18 103
use NAND2X1  _1003_
timestamp 1559787497
transform -1 0 1380 0 1 1305
box -2 -3 26 103
use OAI21X1  _1004_
timestamp 1559787497
transform 1 0 1380 0 1 1305
box -2 -3 34 103
use NAND2X1  _1005_
timestamp 1559787497
transform -1 0 1436 0 1 1305
box -2 -3 26 103
use NAND2X1  _1119_
timestamp 1559787497
transform -1 0 1460 0 1 1305
box -2 -3 26 103
use FILL  FILL_14_1
timestamp 1559787497
transform 1 0 1460 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1559787497
transform 1 0 1468 0 1 1305
box -2 -3 10 103
use NAND2X1  _1290_
timestamp 1559787497
transform 1 0 4 0 -1 1305
box -2 -3 26 103
use OR2X2  _1274_
timestamp 1559787497
transform 1 0 28 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1277_
timestamp 1559787497
transform -1 0 92 0 -1 1305
box -2 -3 34 103
use OR2X2  _1244_
timestamp 1559787497
transform 1 0 92 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1247_
timestamp 1559787497
transform 1 0 124 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1208_
timestamp 1559787497
transform -1 0 188 0 -1 1305
box -2 -3 34 103
use OR2X2  _1205_
timestamp 1559787497
transform -1 0 220 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1246_
timestamp 1559787497
transform -1 0 244 0 -1 1305
box -2 -3 26 103
use INVX1  _1245_
timestamp 1559787497
transform -1 0 260 0 -1 1305
box -2 -3 18 103
use NAND3X1  _1167_
timestamp 1559787497
transform 1 0 260 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1166_
timestamp 1559787497
transform -1 0 316 0 -1 1305
box -2 -3 26 103
use OR2X2  _1164_
timestamp 1559787497
transform -1 0 348 0 -1 1305
box -2 -3 34 103
use INVX1  _913_
timestamp 1559787497
transform 1 0 348 0 -1 1305
box -2 -3 18 103
use NAND2X1  _914_
timestamp 1559787497
transform -1 0 388 0 -1 1305
box -2 -3 26 103
use INVX1  _916_
timestamp 1559787497
transform 1 0 388 0 -1 1305
box -2 -3 18 103
use OAI21X1  _918_
timestamp 1559787497
transform 1 0 404 0 -1 1305
box -2 -3 34 103
use OR2X2  _912_
timestamp 1559787497
transform 1 0 436 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1559787497
transform -1 0 476 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1559787497
transform -1 0 484 0 -1 1305
box -2 -3 10 103
use NAND3X1  _915_
timestamp 1559787497
transform -1 0 516 0 -1 1305
box -2 -3 34 103
use OR2X2  _832_
timestamp 1559787497
transform 1 0 516 0 -1 1305
box -2 -3 34 103
use NAND3X1  _835_
timestamp 1559787497
transform -1 0 580 0 -1 1305
box -2 -3 34 103
use OR2X2  _873_
timestamp 1559787497
transform 1 0 580 0 -1 1305
box -2 -3 34 103
use NAND3X1  _876_
timestamp 1559787497
transform 1 0 612 0 -1 1305
box -2 -3 34 103
use NAND2X1  _875_
timestamp 1559787497
transform 1 0 644 0 -1 1305
box -2 -3 26 103
use INVX1  _874_
timestamp 1559787497
transform -1 0 684 0 -1 1305
box -2 -3 18 103
use OAI21X1  _879_
timestamp 1559787497
transform -1 0 716 0 -1 1305
box -2 -3 34 103
use INVX1  _877_
timestamp 1559787497
transform -1 0 732 0 -1 1305
box -2 -3 18 103
use OAI21X1  _838_
timestamp 1559787497
transform -1 0 764 0 -1 1305
box -2 -3 34 103
use INVX1  _836_
timestamp 1559787497
transform -1 0 780 0 -1 1305
box -2 -3 18 103
use INVX1  _711_
timestamp 1559787497
transform 1 0 780 0 -1 1305
box -2 -3 18 103
use OAI21X1  _713_
timestamp 1559787497
transform 1 0 796 0 -1 1305
box -2 -3 34 103
use OR2X2  _746_
timestamp 1559787497
transform 1 0 828 0 -1 1305
box -2 -3 34 103
use NAND3X1  _749_
timestamp 1559787497
transform -1 0 892 0 -1 1305
box -2 -3 34 103
use INVX1  _1079_
timestamp 1559787497
transform 1 0 892 0 -1 1305
box -2 -3 18 103
use OR2X2  _666_
timestamp 1559787497
transform 1 0 908 0 -1 1305
box -2 -3 34 103
use INVX1  _789_
timestamp 1559787497
transform 1 0 940 0 -1 1305
box -2 -3 18 103
use INVX1  _1121_
timestamp 1559787497
transform 1 0 956 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_1_0
timestamp 1559787497
transform 1 0 972 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1559787497
transform 1 0 980 0 -1 1305
box -2 -3 10 103
use OAI21X1  _791_
timestamp 1559787497
transform 1 0 988 0 -1 1305
box -2 -3 34 103
use INVX1  _1043_
timestamp 1559787497
transform 1 0 1020 0 -1 1305
box -2 -3 18 103
use NAND2X1  _1080_
timestamp 1559787497
transform -1 0 1060 0 -1 1305
box -2 -3 26 103
use OR2X2  _1078_
timestamp 1559787497
transform 1 0 1060 0 -1 1305
box -2 -3 34 103
use OR2X2  _1039_
timestamp 1559787497
transform 1 0 1092 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1081_
timestamp 1559787497
transform -1 0 1156 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_insert7
timestamp 1559787497
transform -1 0 1180 0 -1 1305
box -2 -3 26 103
use NAND3X1  _1042_
timestamp 1559787497
transform 1 0 1180 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1047_
timestamp 1559787497
transform -1 0 1244 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1086_
timestamp 1559787497
transform 1 0 1244 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1125_
timestamp 1559787497
transform 1 0 1276 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1120_
timestamp 1559787497
transform 1 0 1308 0 -1 1305
box -2 -3 34 103
use OR2X2  _1117_
timestamp 1559787497
transform -1 0 1372 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1006_
timestamp 1559787497
transform 1 0 1372 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1001_
timestamp 1559787497
transform -1 0 1436 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1000_
timestamp 1559787497
transform 1 0 1436 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1559787497
transform -1 0 1468 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1559787497
transform -1 0 1476 0 -1 1305
box -2 -3 10 103
use BUFX2  _652_
timestamp 1559787497
transform -1 0 28 0 1 1105
box -2 -3 26 103
use NAND3X1  _1291_
timestamp 1559787497
transform -1 0 60 0 1 1105
box -2 -3 34 103
use INVX4  _1154_
timestamp 1559787497
transform 1 0 60 0 1 1105
box -2 -3 26 103
use NAND3X1  _1282_
timestamp 1559787497
transform -1 0 116 0 1 1105
box -2 -3 34 103
use NAND3X1  _1252_
timestamp 1559787497
transform -1 0 148 0 1 1105
box -2 -3 34 103
use NAND3X1  _1281_
timestamp 1559787497
transform 1 0 148 0 1 1105
box -2 -3 34 103
use NAND3X1  _1213_
timestamp 1559787497
transform 1 0 180 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert39
timestamp 1559787497
transform 1 0 212 0 1 1105
box -2 -3 26 103
use INVX2  _1153_
timestamp 1559787497
transform -1 0 252 0 1 1105
box -2 -3 18 103
use NAND3X1  _1172_
timestamp 1559787497
transform 1 0 252 0 1 1105
box -2 -3 34 103
use OR2X2  _1280_
timestamp 1559787497
transform -1 0 316 0 1 1105
box -2 -3 34 103
use NAND2X1  _1201_
timestamp 1559787497
transform 1 0 316 0 1 1105
box -2 -3 26 103
use INVX1  _1200_
timestamp 1559787497
transform -1 0 356 0 1 1105
box -2 -3 18 103
use NAND3X1  _1286_
timestamp 1559787497
transform -1 0 388 0 1 1105
box -2 -3 34 103
use OR2X2  _1283_
timestamp 1559787497
transform -1 0 420 0 1 1105
box -2 -3 34 103
use INVX1  _1165_
timestamp 1559787497
transform -1 0 436 0 1 1105
box -2 -3 18 103
use OR2X2  _948_
timestamp 1559787497
transform -1 0 468 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1559787497
transform 1 0 468 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1559787497
transform 1 0 476 0 1 1105
box -2 -3 10 103
use INVX1  _943_
timestamp 1559787497
transform 1 0 484 0 1 1105
box -2 -3 18 103
use NAND2X1  _944_
timestamp 1559787497
transform -1 0 524 0 1 1105
box -2 -3 26 103
use NAND2X1  _919_
timestamp 1559787497
transform -1 0 548 0 1 1105
box -2 -3 26 103
use NAND2X1  _834_
timestamp 1559787497
transform 1 0 548 0 1 1105
box -2 -3 26 103
use INVX1  _833_
timestamp 1559787497
transform -1 0 588 0 1 1105
box -2 -3 18 103
use BUFX2  BUFX2_insert13
timestamp 1559787497
transform -1 0 612 0 1 1105
box -2 -3 26 103
use NAND3X1  _959_
timestamp 1559787497
transform 1 0 612 0 1 1105
box -2 -3 34 103
use OR2X2  _951_
timestamp 1559787497
transform 1 0 644 0 1 1105
box -2 -3 34 103
use NAND2X1  _880_
timestamp 1559787497
transform 1 0 676 0 1 1105
box -2 -3 26 103
use NAND3X1  _954_
timestamp 1559787497
transform 1 0 700 0 1 1105
box -2 -3 34 103
use NAND2X1  _839_
timestamp 1559787497
transform -1 0 756 0 1 1105
box -2 -3 26 103
use INVX1  _708_
timestamp 1559787497
transform -1 0 772 0 1 1105
box -2 -3 18 103
use NAND2X1  _709_
timestamp 1559787497
transform -1 0 796 0 1 1105
box -2 -3 26 103
use OR2X2  _707_
timestamp 1559787497
transform -1 0 828 0 1 1105
box -2 -3 34 103
use NAND2X1  _714_
timestamp 1559787497
transform -1 0 852 0 1 1105
box -2 -3 26 103
use NAND3X1  _674_
timestamp 1559787497
transform -1 0 884 0 1 1105
box -2 -3 34 103
use NAND3X1  _754_
timestamp 1559787497
transform 1 0 884 0 1 1105
box -2 -3 34 103
use NAND3X1  _669_
timestamp 1559787497
transform 1 0 916 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert22
timestamp 1559787497
transform 1 0 948 0 1 1105
box -2 -3 26 103
use NAND2X1  _668_
timestamp 1559787497
transform 1 0 972 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1559787497
transform -1 0 1004 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1559787497
transform -1 0 1012 0 1 1105
box -2 -3 10 103
use INVX1  _667_
timestamp 1559787497
transform -1 0 1028 0 1 1105
box -2 -3 18 103
use NAND2X1  _792_
timestamp 1559787497
transform -1 0 1052 0 1 1105
box -2 -3 26 103
use INVX1  _777_
timestamp 1559787497
transform 1 0 1052 0 1 1105
box -2 -3 18 103
use NAND2X1  _778_
timestamp 1559787497
transform -1 0 1092 0 1 1105
box -2 -3 26 103
use NAND3X1  _788_
timestamp 1559787497
transform 1 0 1092 0 1 1105
box -2 -3 34 103
use OR2X2  _785_
timestamp 1559787497
transform -1 0 1156 0 1 1105
box -2 -3 34 103
use NAND2X1  _787_
timestamp 1559787497
transform 1 0 1156 0 1 1105
box -2 -3 26 103
use INVX1  _786_
timestamp 1559787497
transform -1 0 1196 0 1 1105
box -2 -3 18 103
use INVX1  _1109_
timestamp 1559787497
transform 1 0 1196 0 1 1105
box -2 -3 18 103
use OR2X2  _1108_
timestamp 1559787497
transform 1 0 1212 0 1 1105
box -2 -3 34 103
use NAND2X1  _1110_
timestamp 1559787497
transform 1 0 1244 0 1 1105
box -2 -3 26 103
use NAND3X1  _1111_
timestamp 1559787497
transform -1 0 1300 0 1 1105
box -2 -3 34 103
use NAND3X1  _1116_
timestamp 1559787497
transform 1 0 1300 0 1 1105
box -2 -3 34 103
use INVX2  _987_
timestamp 1559787497
transform -1 0 1348 0 1 1105
box -2 -3 18 103
use NAND3X1  _1115_
timestamp 1559787497
transform 1 0 1348 0 1 1105
box -2 -3 34 103
use OR2X2  _1114_
timestamp 1559787497
transform -1 0 1412 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert9
timestamp 1559787497
transform 1 0 1412 0 1 1105
box -2 -3 26 103
use NAND2X1  _1113_
timestamp 1559787497
transform -1 0 1460 0 1 1105
box -2 -3 26 103
use INVX1  _999_
timestamp 1559787497
transform -1 0 1476 0 1 1105
box -2 -3 18 103
use DFFPOSX1  _1316_
timestamp 1559787497
transform -1 0 100 0 -1 1105
box -2 -3 98 103
use NAND3X1  _1292_
timestamp 1559787497
transform -1 0 132 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1214_
timestamp 1559787497
transform 1 0 132 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1279_
timestamp 1559787497
transform -1 0 188 0 -1 1105
box -2 -3 26 103
use INVX1  _1278_
timestamp 1559787497
transform -1 0 204 0 -1 1105
box -2 -3 18 103
use BUFX2  BUFX2_insert36
timestamp 1559787497
transform -1 0 228 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert35
timestamp 1559787497
transform 1 0 228 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1204_
timestamp 1559787497
transform 1 0 252 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1203_
timestamp 1559787497
transform 1 0 284 0 -1 1105
box -2 -3 34 103
use OR2X2  _1202_
timestamp 1559787497
transform -1 0 348 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1285_
timestamp 1559787497
transform 1 0 348 0 -1 1105
box -2 -3 26 103
use INVX1  _1284_
timestamp 1559787497
transform -1 0 388 0 -1 1105
box -2 -3 18 103
use INVX1  _946_
timestamp 1559787497
transform 1 0 388 0 -1 1105
box -2 -3 18 103
use NAND2X1  _947_
timestamp 1559787497
transform -1 0 428 0 -1 1105
box -2 -3 26 103
use NAND3X1  _949_
timestamp 1559787497
transform -1 0 460 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1559787497
transform 1 0 460 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1559787497
transform 1 0 468 0 -1 1105
box -2 -3 10 103
use OR2X2  _942_
timestamp 1559787497
transform 1 0 476 0 -1 1105
box -2 -3 34 103
use NAND3X1  _945_
timestamp 1559787497
transform -1 0 540 0 -1 1105
box -2 -3 34 103
use NAND3X1  _920_
timestamp 1559787497
transform -1 0 572 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert14
timestamp 1559787497
transform -1 0 596 0 -1 1105
box -2 -3 26 103
use NAND3X1  _840_
timestamp 1559787497
transform 1 0 596 0 -1 1105
box -2 -3 34 103
use INVX1  _868_
timestamp 1559787497
transform 1 0 628 0 -1 1105
box -2 -3 18 103
use INVX2  _821_
timestamp 1559787497
transform 1 0 644 0 -1 1105
box -2 -3 18 103
use NAND3X1  _881_
timestamp 1559787497
transform 1 0 660 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert10
timestamp 1559787497
transform 1 0 692 0 -1 1105
box -2 -3 26 103
use NAND2X1  _953_
timestamp 1559787497
transform 1 0 716 0 -1 1105
box -2 -3 26 103
use INVX1  _952_
timestamp 1559787497
transform -1 0 756 0 -1 1105
box -2 -3 18 103
use INVX4  _822_
timestamp 1559787497
transform 1 0 756 0 -1 1105
box -2 -3 26 103
use NAND3X1  _710_
timestamp 1559787497
transform -1 0 812 0 -1 1105
box -2 -3 34 103
use NAND3X1  _715_
timestamp 1559787497
transform -1 0 844 0 -1 1105
box -2 -3 34 103
use INVX1  _702_
timestamp 1559787497
transform 1 0 844 0 -1 1105
box -2 -3 18 103
use NAND2X1  _703_
timestamp 1559787497
transform 1 0 860 0 -1 1105
box -2 -3 26 103
use NAND3X1  _705_
timestamp 1559787497
transform -1 0 916 0 -1 1105
box -2 -3 34 103
use OR2X2  _704_
timestamp 1559787497
transform -1 0 948 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert23
timestamp 1559787497
transform 1 0 948 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1559787497
transform 1 0 972 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1559787497
transform 1 0 980 0 -1 1105
box -2 -3 10 103
use OR2X2  _776_
timestamp 1559787497
transform 1 0 988 0 -1 1105
box -2 -3 34 103
use NAND3X1  _793_
timestamp 1559787497
transform 1 0 1020 0 -1 1105
box -2 -3 34 103
use NAND3X1  _779_
timestamp 1559787497
transform -1 0 1084 0 -1 1105
box -2 -3 34 103
use NAND3X1  _783_
timestamp 1559787497
transform 1 0 1084 0 -1 1105
box -2 -3 34 103
use OR2X2  _782_
timestamp 1559787497
transform -1 0 1148 0 -1 1105
box -2 -3 34 103
use NAND2X1  _781_
timestamp 1559787497
transform 1 0 1148 0 -1 1105
box -2 -3 26 103
use INVX1  _780_
timestamp 1559787497
transform 1 0 1172 0 -1 1105
box -2 -3 18 103
use INVX1  _1034_
timestamp 1559787497
transform 1 0 1188 0 -1 1105
box -2 -3 18 103
use NAND2X1  _1035_
timestamp 1559787497
transform -1 0 1228 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1048_
timestamp 1559787497
transform -1 0 1260 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1038_
timestamp 1559787497
transform -1 0 1292 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1126_
timestamp 1559787497
transform -1 0 1324 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert5
timestamp 1559787497
transform -1 0 1348 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1037_
timestamp 1559787497
transform -1 0 1380 0 -1 1105
box -2 -3 34 103
use OR2X2  _1036_
timestamp 1559787497
transform -1 0 1412 0 -1 1105
box -2 -3 34 103
use NAND3X1  _992_
timestamp 1559787497
transform 1 0 1412 0 -1 1105
box -2 -3 34 103
use OR2X2  _989_
timestamp 1559787497
transform -1 0 1476 0 -1 1105
box -2 -3 34 103
use BUFX2  _649_
timestamp 1559787497
transform -1 0 28 0 1 905
box -2 -3 26 103
use DFFPOSX1  _1313_
timestamp 1559787497
transform -1 0 124 0 1 905
box -2 -3 98 103
use AOI21X1  _1312_
timestamp 1559787497
transform 1 0 124 0 1 905
box -2 -3 34 103
use INVX2  _1152_
timestamp 1559787497
transform 1 0 156 0 1 905
box -2 -3 18 103
use AOI21X1  _1195_
timestamp 1559787497
transform -1 0 204 0 1 905
box -2 -3 34 103
use NAND3X1  _1253_
timestamp 1559787497
transform -1 0 236 0 1 905
box -2 -3 34 103
use NAND3X1  _1173_
timestamp 1559787497
transform 1 0 236 0 1 905
box -2 -3 34 103
use NAND3X1  _1243_
timestamp 1559787497
transform 1 0 268 0 1 905
box -2 -3 34 103
use NAND3X1  _1163_
timestamp 1559787497
transform 1 0 300 0 1 905
box -2 -3 34 103
use NAND3X1  _1162_
timestamp 1559787497
transform 1 0 332 0 1 905
box -2 -3 34 103
use OR2X2  _1161_
timestamp 1559787497
transform -1 0 396 0 1 905
box -2 -3 34 103
use NAND3X1  _1242_
timestamp 1559787497
transform 1 0 396 0 1 905
box -2 -3 34 103
use NAND3X1  _1158_
timestamp 1559787497
transform 1 0 428 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1559787497
transform -1 0 468 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1559787497
transform -1 0 476 0 1 905
box -2 -3 10 103
use OR2X2  _1155_
timestamp 1559787497
transform -1 0 508 0 1 905
box -2 -3 34 103
use NAND3X1  _1199_
timestamp 1559787497
transform 1 0 508 0 1 905
box -2 -3 34 103
use OR2X2  _1196_
timestamp 1559787497
transform -1 0 572 0 1 905
box -2 -3 34 103
use NAND2X1  _1198_
timestamp 1559787497
transform 1 0 572 0 1 905
box -2 -3 26 103
use NAND3X1  _950_
timestamp 1559787497
transform -1 0 628 0 1 905
box -2 -3 34 103
use INVX1  _1197_
timestamp 1559787497
transform -1 0 644 0 1 905
box -2 -3 18 103
use NAND2X1  _869_
timestamp 1559787497
transform -1 0 668 0 1 905
box -2 -3 26 103
use OR2X2  _870_
timestamp 1559787497
transform 1 0 668 0 1 905
box -2 -3 34 103
use NAND3X1  _871_
timestamp 1559787497
transform -1 0 732 0 1 905
box -2 -3 34 103
use NAND3X1  _872_
timestamp 1559787497
transform 1 0 732 0 1 905
box -2 -3 34 103
use NAND3X1  _867_
timestamp 1559787497
transform 1 0 764 0 1 905
box -2 -3 34 103
use OR2X2  _864_
timestamp 1559787497
transform -1 0 828 0 1 905
box -2 -3 34 103
use INVX1  _699_
timestamp 1559787497
transform 1 0 828 0 1 905
box -2 -3 18 103
use NAND2X1  _700_
timestamp 1559787497
transform 1 0 844 0 1 905
box -2 -3 26 103
use NAND3X1  _706_
timestamp 1559787497
transform 1 0 868 0 1 905
box -2 -3 34 103
use NAND3X1  _701_
timestamp 1559787497
transform -1 0 932 0 1 905
box -2 -3 34 103
use OR2X2  _698_
timestamp 1559787497
transform -1 0 964 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_insert24
timestamp 1559787497
transform -1 0 988 0 1 905
box -2 -3 26 103
use FILL  FILL_9_1_0
timestamp 1559787497
transform 1 0 988 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1559787497
transform 1 0 996 0 1 905
box -2 -3 10 103
use BUFX2  BUFX2_insert21
timestamp 1559787497
transform 1 0 1004 0 1 905
box -2 -3 26 103
use NAND3X1  _784_
timestamp 1559787497
transform 1 0 1028 0 1 905
box -2 -3 34 103
use NAND2X1  _659_
timestamp 1559787497
transform 1 0 1060 0 1 905
box -2 -3 26 103
use INVX1  _658_
timestamp 1559787497
transform -1 0 1100 0 1 905
box -2 -3 18 103
use INVX1  _741_
timestamp 1559787497
transform 1 0 1100 0 1 905
box -2 -3 18 103
use NAND2X1  _742_
timestamp 1559787497
transform -1 0 1140 0 1 905
box -2 -3 26 103
use INVX1  _1031_
timestamp 1559787497
transform -1 0 1156 0 1 905
box -2 -3 18 103
use NAND2X1  _1032_
timestamp 1559787497
transform -1 0 1180 0 1 905
box -2 -3 26 103
use NAND3X1  _1033_
timestamp 1559787497
transform -1 0 1212 0 1 905
box -2 -3 34 103
use OR2X2  _1030_
timestamp 1559787497
transform 1 0 1212 0 1 905
box -2 -3 34 103
use INVX4  _988_
timestamp 1559787497
transform -1 0 1268 0 1 905
box -2 -3 26 103
use INVX1  _1070_
timestamp 1559787497
transform 1 0 1268 0 1 905
box -2 -3 18 103
use NAND2X1  _1071_
timestamp 1559787497
transform -1 0 1308 0 1 905
box -2 -3 26 103
use NAND3X1  _997_
timestamp 1559787497
transform -1 0 1340 0 1 905
box -2 -3 34 103
use NAND3X1  _996_
timestamp 1559787497
transform 1 0 1340 0 1 905
box -2 -3 34 103
use OR2X2  _995_
timestamp 1559787497
transform -1 0 1404 0 1 905
box -2 -3 34 103
use INVX1  _993_
timestamp 1559787497
transform 1 0 1404 0 1 905
box -2 -3 18 103
use NAND2X1  _994_
timestamp 1559787497
transform -1 0 1444 0 1 905
box -2 -3 26 103
use NAND2X1  _991_
timestamp 1559787497
transform -1 0 1468 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1559787497
transform 1 0 1468 0 1 905
box -2 -3 10 103
use BUFX2  _650_
timestamp 1559787497
transform -1 0 28 0 -1 905
box -2 -3 26 103
use DFFPOSX1  _1314_
timestamp 1559787497
transform -1 0 124 0 -1 905
box -2 -3 98 103
use AOI21X1  _1234_
timestamp 1559787497
transform 1 0 124 0 -1 905
box -2 -3 34 103
use BUFX2  _638_
timestamp 1559787497
transform -1 0 180 0 -1 905
box -2 -3 26 103
use DFFPOSX1  _816_
timestamp 1559787497
transform -1 0 276 0 -1 905
box -2 -3 98 103
use NAND3X1  _1238_
timestamp 1559787497
transform 1 0 276 0 -1 905
box -2 -3 34 103
use OR2X2  _1235_
timestamp 1559787497
transform -1 0 340 0 -1 905
box -2 -3 34 103
use NAND2X1  _1237_
timestamp 1559787497
transform -1 0 364 0 -1 905
box -2 -3 26 103
use INVX1  _1236_
timestamp 1559787497
transform -1 0 380 0 -1 905
box -2 -3 18 103
use NAND2X1  _1160_
timestamp 1559787497
transform 1 0 380 0 -1 905
box -2 -3 26 103
use NAND2X1  _1240_
timestamp 1559787497
transform 1 0 404 0 -1 905
box -2 -3 26 103
use INVX1  _1159_
timestamp 1559787497
transform -1 0 444 0 -1 905
box -2 -3 18 103
use OR2X2  _1241_
timestamp 1559787497
transform -1 0 476 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1559787497
transform 1 0 476 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1559787497
transform 1 0 484 0 -1 905
box -2 -3 10 103
use NAND2X1  _1157_
timestamp 1559787497
transform 1 0 492 0 -1 905
box -2 -3 26 103
use INVX1  _1156_
timestamp 1559787497
transform -1 0 532 0 -1 905
box -2 -3 18 103
use OR2X2  _823_
timestamp 1559787497
transform 1 0 532 0 -1 905
box -2 -3 34 103
use NAND3X1  _826_
timestamp 1559787497
transform 1 0 564 0 -1 905
box -2 -3 34 103
use NAND2X1  _825_
timestamp 1559787497
transform 1 0 596 0 -1 905
box -2 -3 26 103
use INVX1  _824_
timestamp 1559787497
transform -1 0 636 0 -1 905
box -2 -3 18 103
use NAND3X1  _960_
timestamp 1559787497
transform -1 0 668 0 -1 905
box -2 -3 34 103
use NAND3X1  _882_
timestamp 1559787497
transform -1 0 700 0 -1 905
box -2 -3 34 103
use INVX1  _904_
timestamp 1559787497
transform 1 0 700 0 -1 905
box -2 -3 18 103
use NAND2X1  _905_
timestamp 1559787497
transform -1 0 740 0 -1 905
box -2 -3 26 103
use NAND3X1  _906_
timestamp 1559787497
transform -1 0 772 0 -1 905
box -2 -3 34 103
use OR2X2  _903_
timestamp 1559787497
transform -1 0 804 0 -1 905
box -2 -3 34 103
use INVX1  _865_
timestamp 1559787497
transform 1 0 804 0 -1 905
box -2 -3 18 103
use NAND2X1  _866_
timestamp 1559787497
transform -1 0 844 0 -1 905
box -2 -3 26 103
use NAND3X1  _716_
timestamp 1559787497
transform -1 0 876 0 -1 905
box -2 -3 34 103
use NAND3X1  _910_
timestamp 1559787497
transform 1 0 876 0 -1 905
box -2 -3 34 103
use OR2X2  _909_
timestamp 1559787497
transform -1 0 940 0 -1 905
box -2 -3 34 103
use NAND2X1  _908_
timestamp 1559787497
transform 1 0 940 0 -1 905
box -2 -3 26 103
use INVX1  _907_
timestamp 1559787497
transform -1 0 980 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_1_0
timestamp 1559787497
transform -1 0 988 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1559787497
transform -1 0 996 0 -1 905
box -2 -3 10 103
use INVX1  _1239_
timestamp 1559787497
transform -1 0 1012 0 -1 905
box -2 -3 18 103
use INVX2  _655_
timestamp 1559787497
transform 1 0 1012 0 -1 905
box -2 -3 18 103
use NAND3X1  _794_
timestamp 1559787497
transform 1 0 1028 0 -1 905
box -2 -3 34 103
use NAND3X1  _660_
timestamp 1559787497
transform 1 0 1060 0 -1 905
box -2 -3 34 103
use INVX4  _656_
timestamp 1559787497
transform 1 0 1092 0 -1 905
box -2 -3 26 103
use OR2X2  _657_
timestamp 1559787497
transform -1 0 1148 0 -1 905
box -2 -3 34 103
use NAND3X1  _740_
timestamp 1559787497
transform 1 0 1148 0 -1 905
box -2 -3 34 103
use OR2X2  _737_
timestamp 1559787497
transform -1 0 1212 0 -1 905
box -2 -3 34 103
use NAND2X1  _739_
timestamp 1559787497
transform 1 0 1212 0 -1 905
box -2 -3 26 103
use INVX1  _738_
timestamp 1559787497
transform 1 0 1236 0 -1 905
box -2 -3 18 103
use INVX1  _1073_
timestamp 1559787497
transform 1 0 1252 0 -1 905
box -2 -3 18 103
use NAND2X1  _1074_
timestamp 1559787497
transform -1 0 1292 0 -1 905
box -2 -3 26 103
use NAND3X1  _1076_
timestamp 1559787497
transform -1 0 1324 0 -1 905
box -2 -3 34 103
use NAND3X1  _1077_
timestamp 1559787497
transform -1 0 1356 0 -1 905
box -2 -3 34 103
use NAND3X1  _1007_
timestamp 1559787497
transform 1 0 1356 0 -1 905
box -2 -3 34 103
use NAND3X1  _1072_
timestamp 1559787497
transform -1 0 1420 0 -1 905
box -2 -3 34 103
use OR2X2  _1075_
timestamp 1559787497
transform -1 0 1452 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1559787497
transform -1 0 1460 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1559787497
transform -1 0 1468 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_3
timestamp 1559787497
transform -1 0 1476 0 -1 905
box -2 -3 10 103
use BUFX2  _651_
timestamp 1559787497
transform -1 0 28 0 1 705
box -2 -3 26 103
use BUFX2  _642_
timestamp 1559787497
transform -1 0 52 0 1 705
box -2 -3 26 103
use DFFPOSX1  _1315_
timestamp 1559787497
transform -1 0 148 0 1 705
box -2 -3 98 103
use AOI21X1  _1273_
timestamp 1559787497
transform -1 0 180 0 1 705
box -2 -3 34 103
use DFFPOSX1  _982_
timestamp 1559787497
transform -1 0 276 0 1 705
box -2 -3 98 103
use BUFX2  _637_
timestamp 1559787497
transform -1 0 300 0 1 705
box -2 -3 26 103
use DFFPOSX1  _815_
timestamp 1559787497
transform -1 0 396 0 1 705
box -2 -3 98 103
use AOI21X1  _697_
timestamp 1559787497
transform 1 0 396 0 1 705
box -2 -3 34 103
use AOI21X1  _736_
timestamp 1559787497
transform -1 0 460 0 1 705
box -2 -3 34 103
use INVX1  _796_
timestamp 1559787497
transform 1 0 460 0 1 705
box -2 -3 18 103
use FILL  FILL_7_0_0
timestamp 1559787497
transform -1 0 484 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1559787497
transform -1 0 492 0 1 705
box -2 -3 10 103
use NAND2X1  _797_
timestamp 1559787497
transform -1 0 516 0 1 705
box -2 -3 26 103
use OR2X2  _829_
timestamp 1559787497
transform 1 0 516 0 1 705
box -2 -3 34 103
use INVX2  _653_
timestamp 1559787497
transform -1 0 564 0 1 705
box -2 -3 18 103
use NAND3X1  _830_
timestamp 1559787497
transform 1 0 564 0 1 705
box -2 -3 34 103
use NAND3X1  _831_
timestamp 1559787497
transform -1 0 628 0 1 705
box -2 -3 34 103
use NAND3X1  _841_
timestamp 1559787497
transform -1 0 660 0 1 705
box -2 -3 34 103
use NAND3X1  _921_
timestamp 1559787497
transform -1 0 692 0 1 705
box -2 -3 34 103
use INVX2  _654_
timestamp 1559787497
transform -1 0 708 0 1 705
box -2 -3 18 103
use NAND3X1  _911_
timestamp 1559787497
transform 1 0 708 0 1 705
box -2 -3 34 103
use INVX2  _819_
timestamp 1559787497
transform -1 0 756 0 1 705
box -2 -3 18 103
use AOI21X1  _863_
timestamp 1559787497
transform 1 0 756 0 1 705
box -2 -3 34 103
use NAND3X1  _675_
timestamp 1559787497
transform -1 0 820 0 1 705
box -2 -3 34 103
use NAND3X1  _665_
timestamp 1559787497
transform -1 0 852 0 1 705
box -2 -3 34 103
use NAND3X1  _755_
timestamp 1559787497
transform 1 0 852 0 1 705
box -2 -3 34 103
use NAND3X1  _664_
timestamp 1559787497
transform 1 0 884 0 1 705
box -2 -3 34 103
use OR2X2  _663_
timestamp 1559787497
transform -1 0 948 0 1 705
box -2 -3 34 103
use NAND3X1  _745_
timestamp 1559787497
transform 1 0 948 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1559787497
transform 1 0 980 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1559787497
transform 1 0 988 0 1 705
box -2 -3 10 103
use NAND3X1  _744_
timestamp 1559787497
transform 1 0 996 0 1 705
box -2 -3 34 103
use OR2X2  _743_
timestamp 1559787497
transform -1 0 1060 0 1 705
box -2 -3 34 103
use DFFPOSX1  _981_
timestamp 1559787497
transform 1 0 1060 0 1 705
box -2 -3 98 103
use DFFPOSX1  _983_
timestamp 1559787497
transform 1 0 1156 0 1 705
box -2 -3 98 103
use BUFX2  _641_
timestamp 1559787497
transform 1 0 1252 0 1 705
box -2 -3 26 103
use INVX2  _986_
timestamp 1559787497
transform 1 0 1276 0 1 705
box -2 -3 18 103
use NAND3X1  _1087_
timestamp 1559787497
transform -1 0 1324 0 1 705
box -2 -3 34 103
use DFFPOSX1  _1150_
timestamp 1559787497
transform 1 0 1324 0 1 705
box -2 -3 98 103
use BUFX2  _648_
timestamp 1559787497
transform 1 0 1420 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_insert8
timestamp 1559787497
transform -1 0 1468 0 1 705
box -2 -3 26 103
use FILL  FILL_8_1
timestamp 1559787497
transform 1 0 1468 0 1 705
box -2 -3 10 103
use INVX1  _1186_
timestamp 1559787497
transform -1 0 20 0 -1 705
box -2 -3 18 103
use NAND2X1  _1187_
timestamp 1559787497
transform -1 0 44 0 -1 705
box -2 -3 26 103
use OR2X2  _1185_
timestamp 1559787497
transform 1 0 44 0 -1 705
box -2 -3 34 103
use NAND3X1  _1188_
timestamp 1559787497
transform -1 0 108 0 -1 705
box -2 -3 34 103
use OR2X2  _1293_
timestamp 1559787497
transform 1 0 108 0 -1 705
box -2 -3 34 103
use INVX2  _1151_
timestamp 1559787497
transform 1 0 140 0 -1 705
box -2 -3 18 103
use NAND3X1  _1296_
timestamp 1559787497
transform 1 0 156 0 -1 705
box -2 -3 34 103
use NAND2X1  _1295_
timestamp 1559787497
transform 1 0 188 0 -1 705
box -2 -3 26 103
use INVX1  _1294_
timestamp 1559787497
transform -1 0 228 0 -1 705
box -2 -3 18 103
use INVX4  _677_
timestamp 1559787497
transform 1 0 228 0 -1 705
box -2 -3 26 103
use NAND2X1  _694_
timestamp 1559787497
transform 1 0 252 0 -1 705
box -2 -3 26 103
use NAND3X1  _695_
timestamp 1559787497
transform -1 0 308 0 -1 705
box -2 -3 34 103
use NAND3X1  _696_
timestamp 1559787497
transform -1 0 340 0 -1 705
box -2 -3 34 103
use NAND3X1  _812_
timestamp 1559787497
transform -1 0 372 0 -1 705
box -2 -3 34 103
use INVX2  _676_
timestamp 1559787497
transform 1 0 372 0 -1 705
box -2 -3 18 103
use NAND3X1  _686_
timestamp 1559787497
transform 1 0 388 0 -1 705
box -2 -3 34 103
use NAND3X1  _735_
timestamp 1559787497
transform -1 0 452 0 -1 705
box -2 -3 34 103
use NAND3X1  _725_
timestamp 1559787497
transform 1 0 452 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1559787497
transform -1 0 492 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1559787497
transform -1 0 500 0 -1 705
box -2 -3 10 103
use NAND3X1  _798_
timestamp 1559787497
transform -1 0 532 0 -1 705
box -2 -3 34 103
use OR2X2  _795_
timestamp 1559787497
transform -1 0 564 0 -1 705
box -2 -3 34 103
use NAND3X1  _773_
timestamp 1559787497
transform -1 0 596 0 -1 705
box -2 -3 34 103
use NAND3X1  _774_
timestamp 1559787497
transform -1 0 628 0 -1 705
box -2 -3 34 103
use NAND3X1  _803_
timestamp 1559787497
transform 1 0 628 0 -1 705
box -2 -3 34 103
use NAND3X1  _813_
timestamp 1559787497
transform -1 0 692 0 -1 705
box -2 -3 34 103
use NAND2X1  _828_
timestamp 1559787497
transform 1 0 692 0 -1 705
box -2 -3 26 103
use INVX1  _827_
timestamp 1559787497
transform -1 0 732 0 -1 705
box -2 -3 18 103
use AOI21X1  _902_
timestamp 1559787497
transform 1 0 732 0 -1 705
box -2 -3 34 103
use AOI21X1  _980_
timestamp 1559787497
transform 1 0 764 0 -1 705
box -2 -3 34 103
use AOI21X1  _941_
timestamp 1559787497
transform -1 0 828 0 -1 705
box -2 -3 34 103
use INVX2  _985_
timestamp 1559787497
transform 1 0 828 0 -1 705
box -2 -3 18 103
use AOI21X1  _775_
timestamp 1559787497
transform 1 0 844 0 -1 705
box -2 -3 34 103
use AOI21X1  _814_
timestamp 1559787497
transform -1 0 908 0 -1 705
box -2 -3 34 103
use INVX1  _962_
timestamp 1559787497
transform 1 0 908 0 -1 705
box -2 -3 18 103
use INVX1  _1128_
timestamp 1559787497
transform 1 0 924 0 -1 705
box -2 -3 18 103
use NAND2X1  _662_
timestamp 1559787497
transform 1 0 940 0 -1 705
box -2 -3 26 103
use INVX1  _661_
timestamp 1559787497
transform 1 0 964 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_1_0
timestamp 1559787497
transform 1 0 980 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1559787497
transform 1 0 988 0 -1 705
box -2 -3 10 103
use DFFPOSX1  _817_
timestamp 1559787497
transform 1 0 996 0 -1 705
box -2 -3 98 103
use DFFPOSX1  _818_
timestamp 1559787497
transform 1 0 1092 0 -1 705
box -2 -3 98 103
use BUFX2  _640_
timestamp 1559787497
transform 1 0 1188 0 -1 705
box -2 -3 26 103
use BUFX2  _639_
timestamp 1559787497
transform 1 0 1212 0 -1 705
box -2 -3 26 103
use BUFX2  _643_
timestamp 1559787497
transform 1 0 1236 0 -1 705
box -2 -3 26 103
use AOI21X1  _1068_
timestamp 1559787497
transform 1 0 1260 0 -1 705
box -2 -3 34 103
use AOI21X1  _1146_
timestamp 1559787497
transform 1 0 1292 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1148_
timestamp 1559787497
transform 1 0 1324 0 -1 705
box -2 -3 98 103
use BUFX2  _646_
timestamp 1559787497
transform 1 0 1420 0 -1 705
box -2 -3 26 103
use BUFX2  _647_
timestamp 1559787497
transform -1 0 1468 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1559787497
transform -1 0 1476 0 -1 705
box -2 -3 10 103
use INVX1  _1297_
timestamp 1559787497
transform 1 0 4 0 1 505
box -2 -3 18 103
use NAND2X1  _1298_
timestamp 1559787497
transform -1 0 44 0 1 505
box -2 -3 26 103
use OR2X2  _1299_
timestamp 1559787497
transform 1 0 44 0 1 505
box -2 -3 34 103
use NAND3X1  _1300_
timestamp 1559787497
transform -1 0 108 0 1 505
box -2 -3 34 103
use NAND3X1  _1193_
timestamp 1559787497
transform 1 0 108 0 1 505
box -2 -3 34 103
use NAND3X1  _1301_
timestamp 1559787497
transform -1 0 172 0 1 505
box -2 -3 34 103
use NAND3X1  _1194_
timestamp 1559787497
transform 1 0 172 0 1 505
box -2 -3 34 103
use INVX4  _1175_
timestamp 1559787497
transform -1 0 228 0 1 505
box -2 -3 26 103
use INVX1  _688_
timestamp 1559787497
transform 1 0 228 0 1 505
box -2 -3 18 103
use NAND2X1  _689_
timestamp 1559787497
transform -1 0 268 0 1 505
box -2 -3 26 103
use INVX1  _691_
timestamp 1559787497
transform 1 0 268 0 1 505
box -2 -3 18 103
use OAI21X1  _693_
timestamp 1559787497
transform 1 0 284 0 1 505
box -2 -3 34 103
use NAND3X1  _690_
timestamp 1559787497
transform -1 0 348 0 1 505
box -2 -3 34 103
use OR2X2  _687_
timestamp 1559787497
transform -1 0 380 0 1 505
box -2 -3 34 103
use OR2X2  _678_
timestamp 1559787497
transform 1 0 380 0 1 505
box -2 -3 34 103
use NAND3X1  _681_
timestamp 1559787497
transform 1 0 412 0 1 505
box -2 -3 34 103
use NAND3X1  _734_
timestamp 1559787497
transform -1 0 476 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1559787497
transform 1 0 476 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1559787497
transform 1 0 484 0 1 505
box -2 -3 10 103
use NAND3X1  _685_
timestamp 1559787497
transform 1 0 492 0 1 505
box -2 -3 34 103
use NAND3X1  _724_
timestamp 1559787497
transform -1 0 556 0 1 505
box -2 -3 34 103
use NAND3X1  _763_
timestamp 1559787497
transform 1 0 556 0 1 505
box -2 -3 34 103
use NAND3X1  _764_
timestamp 1559787497
transform 1 0 588 0 1 505
box -2 -3 34 103
use NAND3X1  _768_
timestamp 1559787497
transform 1 0 620 0 1 505
box -2 -3 34 103
use NAND3X1  _802_
timestamp 1559787497
transform 1 0 652 0 1 505
box -2 -3 34 103
use OR2X2  _801_
timestamp 1559787497
transform -1 0 716 0 1 505
box -2 -3 34 103
use NAND2X1  _800_
timestamp 1559787497
transform 1 0 716 0 1 505
box -2 -3 26 103
use INVX1  _799_
timestamp 1559787497
transform -1 0 756 0 1 505
box -2 -3 18 103
use INVX1  _854_
timestamp 1559787497
transform 1 0 756 0 1 505
box -2 -3 18 103
use NAND2X1  _855_
timestamp 1559787497
transform -1 0 796 0 1 505
box -2 -3 26 103
use INVX2  _820_
timestamp 1559787497
transform -1 0 812 0 1 505
box -2 -3 18 103
use DFFPOSX1  _984_
timestamp 1559787497
transform 1 0 812 0 1 505
box -2 -3 98 103
use NAND2X1  _966_
timestamp 1559787497
transform 1 0 908 0 1 505
box -2 -3 26 103
use INVX1  _965_
timestamp 1559787497
transform -1 0 948 0 1 505
box -2 -3 18 103
use NAND2X1  _963_
timestamp 1559787497
transform -1 0 972 0 1 505
box -2 -3 26 103
use INVX1  _1020_
timestamp 1559787497
transform 1 0 972 0 1 505
box -2 -3 18 103
use FILL  FILL_5_1_0
timestamp 1559787497
transform 1 0 988 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1559787497
transform 1 0 996 0 1 505
box -2 -3 10 103
use OR2X2  _961_
timestamp 1559787497
transform 1 0 1004 0 1 505
box -2 -3 34 103
use OR2X2  _1127_
timestamp 1559787497
transform 1 0 1036 0 1 505
box -2 -3 34 103
use OR2X2  _1133_
timestamp 1559787497
transform 1 0 1068 0 1 505
box -2 -3 34 103
use NAND2X1  _1129_
timestamp 1559787497
transform -1 0 1124 0 1 505
box -2 -3 26 103
use NAND2X1  _1021_
timestamp 1559787497
transform -1 0 1148 0 1 505
box -2 -3 26 103
use NAND3X1  _1130_
timestamp 1559787497
transform -1 0 1180 0 1 505
box -2 -3 34 103
use INVX1  _1131_
timestamp 1559787497
transform -1 0 1196 0 1 505
box -2 -3 18 103
use NAND2X1  _1132_
timestamp 1559787497
transform -1 0 1220 0 1 505
box -2 -3 26 103
use NAND3X1  _1134_
timestamp 1559787497
transform -1 0 1252 0 1 505
box -2 -3 34 103
use NAND3X1  _1135_
timestamp 1559787497
transform -1 0 1284 0 1 505
box -2 -3 34 103
use NAND3X1  _1145_
timestamp 1559787497
transform -1 0 1316 0 1 505
box -2 -3 34 103
use AOI21X1  _1107_
timestamp 1559787497
transform 1 0 1316 0 1 505
box -2 -3 34 103
use AOI21X1  _1029_
timestamp 1559787497
transform -1 0 1380 0 1 505
box -2 -3 34 103
use DFFPOSX1  _1149_
timestamp 1559787497
transform 1 0 1380 0 1 505
box -2 -3 98 103
use INVX1  _1189_
timestamp 1559787497
transform 1 0 4 0 -1 505
box -2 -3 18 103
use OAI21X1  _1191_
timestamp 1559787497
transform 1 0 20 0 -1 505
box -2 -3 34 103
use NAND2X1  _1190_
timestamp 1559787497
transform 1 0 52 0 -1 505
box -2 -3 26 103
use NAND2X1  _1192_
timestamp 1559787497
transform -1 0 100 0 -1 505
box -2 -3 26 103
use NAND3X1  _1183_
timestamp 1559787497
transform -1 0 132 0 -1 505
box -2 -3 34 103
use NAND3X1  _1311_
timestamp 1559787497
transform 1 0 132 0 -1 505
box -2 -3 34 103
use OR2X2  _1182_
timestamp 1559787497
transform -1 0 196 0 -1 505
box -2 -3 34 103
use NAND3X1  _1184_
timestamp 1559787497
transform 1 0 196 0 -1 505
box -2 -3 34 103
use NAND3X1  _1179_
timestamp 1559787497
transform 1 0 228 0 -1 505
box -2 -3 34 103
use OR2X2  _1176_
timestamp 1559787497
transform -1 0 292 0 -1 505
box -2 -3 34 103
use NAND2X1  _1178_
timestamp 1559787497
transform 1 0 292 0 -1 505
box -2 -3 26 103
use NAND2X1  _692_
timestamp 1559787497
transform -1 0 340 0 -1 505
box -2 -3 26 103
use NAND2X1  _811_
timestamp 1559787497
transform 1 0 340 0 -1 505
box -2 -3 26 103
use OR2X2  _684_
timestamp 1559787497
transform 1 0 364 0 -1 505
box -2 -3 34 103
use BUFX2  BUFX2_insert30
timestamp 1559787497
transform -1 0 420 0 -1 505
box -2 -3 26 103
use NAND2X1  _680_
timestamp 1559787497
transform 1 0 420 0 -1 505
box -2 -3 26 103
use NAND2X1  _733_
timestamp 1559787497
transform -1 0 468 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1559787497
transform -1 0 476 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1559787497
transform -1 0 484 0 -1 505
box -2 -3 10 103
use INVX1  _679_
timestamp 1559787497
transform -1 0 500 0 -1 505
box -2 -3 18 103
use INVX1  _1177_
timestamp 1559787497
transform -1 0 516 0 -1 505
box -2 -3 18 103
use NAND2X1  _722_
timestamp 1559787497
transform -1 0 540 0 -1 505
box -2 -3 26 103
use OR2X2  _723_
timestamp 1559787497
transform -1 0 572 0 -1 505
box -2 -3 34 103
use NAND2X1  _772_
timestamp 1559787497
transform -1 0 596 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_insert32
timestamp 1559787497
transform 1 0 596 0 -1 505
box -2 -3 26 103
use NAND2X1  _761_
timestamp 1559787497
transform 1 0 620 0 -1 505
box -2 -3 26 103
use OR2X2  _765_
timestamp 1559787497
transform -1 0 676 0 -1 505
box -2 -3 34 103
use INVX1  _857_
timestamp 1559787497
transform 1 0 676 0 -1 505
box -2 -3 18 103
use NAND2X1  _767_
timestamp 1559787497
transform 1 0 692 0 -1 505
box -2 -3 26 103
use INVX4  _843_
timestamp 1559787497
transform -1 0 740 0 -1 505
box -2 -3 26 103
use OR2X2  _853_
timestamp 1559787497
transform -1 0 772 0 -1 505
box -2 -3 34 103
use NAND3X1  _856_
timestamp 1559787497
transform -1 0 804 0 -1 505
box -2 -3 34 103
use NAND3X1  _979_
timestamp 1559787497
transform -1 0 836 0 -1 505
box -2 -3 34 103
use NAND3X1  _969_
timestamp 1559787497
transform 1 0 836 0 -1 505
box -2 -3 34 103
use NAND3X1  _968_
timestamp 1559787497
transform 1 0 868 0 -1 505
box -2 -3 34 103
use BUFX2  _644_
timestamp 1559787497
transform 1 0 900 0 -1 505
box -2 -3 26 103
use OR2X2  _967_
timestamp 1559787497
transform -1 0 956 0 -1 505
box -2 -3 34 103
use NAND3X1  _964_
timestamp 1559787497
transform -1 0 988 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1559787497
transform 1 0 988 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1559787497
transform 1 0 996 0 -1 505
box -2 -3 10 103
use INVX1  _1023_
timestamp 1559787497
transform 1 0 1004 0 -1 505
box -2 -3 18 103
use NAND2X1  _1024_
timestamp 1559787497
transform -1 0 1044 0 -1 505
box -2 -3 26 103
use OAI21X1  _1025_
timestamp 1559787497
transform 1 0 1044 0 -1 505
box -2 -3 34 103
use OR2X2  _1055_
timestamp 1559787497
transform 1 0 1076 0 -1 505
box -2 -3 34 103
use OR2X2  _1019_
timestamp 1559787497
transform 1 0 1108 0 -1 505
box -2 -3 34 103
use NAND3X1  _1022_
timestamp 1559787497
transform 1 0 1140 0 -1 505
box -2 -3 34 103
use NAND2X1  _1026_
timestamp 1559787497
transform -1 0 1196 0 -1 505
box -2 -3 26 103
use NAND3X1  _1027_
timestamp 1559787497
transform -1 0 1228 0 -1 505
box -2 -3 34 103
use NAND3X1  _1056_
timestamp 1559787497
transform 1 0 1228 0 -1 505
box -2 -3 34 103
use NAND3X1  _1057_
timestamp 1559787497
transform -1 0 1292 0 -1 505
box -2 -3 34 103
use NAND3X1  _1067_
timestamp 1559787497
transform 1 0 1292 0 -1 505
box -2 -3 34 103
use INVX4  _1009_
timestamp 1559787497
transform 1 0 1324 0 -1 505
box -2 -3 26 103
use DFFPOSX1  _1147_
timestamp 1559787497
transform 1 0 1348 0 -1 505
box -2 -3 98 103
use FILL  FILL_5_1
timestamp 1559787497
transform -1 0 1452 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1559787497
transform -1 0 1460 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_3
timestamp 1559787497
transform -1 0 1468 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_4
timestamp 1559787497
transform -1 0 1476 0 -1 505
box -2 -3 10 103
use BUFX2  BUFX2_insert4
timestamp 1559787497
transform 1 0 4 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert2
timestamp 1559787497
transform 1 0 28 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert1
timestamp 1559787497
transform 1 0 52 0 1 305
box -2 -3 26 103
use INVX1  _1180_
timestamp 1559787497
transform 1 0 76 0 1 305
box -2 -3 18 103
use NAND2X1  _1181_
timestamp 1559787497
transform 1 0 92 0 1 305
box -2 -3 26 103
use NAND3X1  _1233_
timestamp 1559787497
transform 1 0 116 0 1 305
box -2 -3 34 103
use INVX2  _1174_
timestamp 1559787497
transform -1 0 164 0 1 305
box -2 -3 18 103
use NAND3X1  _1272_
timestamp 1559787497
transform 1 0 164 0 1 305
box -2 -3 34 103
use NAND3X1  _1271_
timestamp 1559787497
transform 1 0 196 0 1 305
box -2 -3 34 103
use NAND3X1  _1266_
timestamp 1559787497
transform 1 0 228 0 1 305
box -2 -3 34 103
use OR2X2  _1263_
timestamp 1559787497
transform -1 0 292 0 1 305
box -2 -3 34 103
use NAND2X1  _1304_
timestamp 1559787497
transform 1 0 292 0 1 305
box -2 -3 26 103
use NAND2X1  _1265_
timestamp 1559787497
transform 1 0 316 0 1 305
box -2 -3 26 103
use INVX1  _1264_
timestamp 1559787497
transform -1 0 356 0 1 305
box -2 -3 18 103
use INVX1  _1303_
timestamp 1559787497
transform -1 0 372 0 1 305
box -2 -3 18 103
use NAND3X1  _807_
timestamp 1559787497
transform 1 0 372 0 1 305
box -2 -3 34 103
use NAND2X1  _806_
timestamp 1559787497
transform 1 0 404 0 1 305
box -2 -3 26 103
use INVX1  _805_
timestamp 1559787497
transform -1 0 444 0 1 305
box -2 -3 18 103
use NAND3X1  _729_
timestamp 1559787497
transform 1 0 444 0 1 305
box -2 -3 34 103
use FILL  FILL_3_0_0
timestamp 1559787497
transform 1 0 476 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1559787497
transform 1 0 484 0 1 305
box -2 -3 10 103
use INVX1  _682_
timestamp 1559787497
transform 1 0 492 0 1 305
box -2 -3 18 103
use NAND2X1  _683_
timestamp 1559787497
transform 1 0 508 0 1 305
box -2 -3 26 103
use INVX1  _721_
timestamp 1559787497
transform 1 0 532 0 1 305
box -2 -3 18 103
use NAND3X1  _720_
timestamp 1559787497
transform -1 0 580 0 1 305
box -2 -3 34 103
use NAND3X1  _759_
timestamp 1559787497
transform -1 0 612 0 1 305
box -2 -3 34 103
use OR2X2  _717_
timestamp 1559787497
transform -1 0 644 0 1 305
box -2 -3 34 103
use INVX1  _760_
timestamp 1559787497
transform 1 0 644 0 1 305
box -2 -3 18 103
use INVX1  _1014_
timestamp 1559787497
transform 1 0 660 0 1 305
box -2 -3 18 103
use OAI21X1  _859_
timestamp 1559787497
transform 1 0 676 0 1 305
box -2 -3 34 103
use INVX1  _766_
timestamp 1559787497
transform 1 0 708 0 1 305
box -2 -3 18 103
use NAND2X1  _858_
timestamp 1559787497
transform -1 0 748 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert29
timestamp 1559787497
transform -1 0 772 0 1 305
box -2 -3 26 103
use NAND2X1  _860_
timestamp 1559787497
transform -1 0 796 0 1 305
box -2 -3 26 103
use NAND3X1  _861_
timestamp 1559787497
transform -1 0 828 0 1 305
box -2 -3 34 103
use NAND3X1  _862_
timestamp 1559787497
transform 1 0 828 0 1 305
box -2 -3 34 103
use INVX2  _842_
timestamp 1559787497
transform 1 0 860 0 1 305
box -2 -3 18 103
use OR2X2  _850_
timestamp 1559787497
transform 1 0 876 0 1 305
box -2 -3 34 103
use NAND3X1  _851_
timestamp 1559787497
transform -1 0 940 0 1 305
box -2 -3 34 103
use NAND3X1  _852_
timestamp 1559787497
transform 1 0 940 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert25
timestamp 1559787497
transform -1 0 996 0 1 305
box -2 -3 26 103
use FILL  FILL_3_1_0
timestamp 1559787497
transform 1 0 996 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1559787497
transform 1 0 1004 0 1 305
box -2 -3 10 103
use NAND3X1  _847_
timestamp 1559787497
transform 1 0 1012 0 1 305
box -2 -3 34 103
use OR2X2  _844_
timestamp 1559787497
transform -1 0 1076 0 1 305
box -2 -3 34 103
use NAND2X1  _846_
timestamp 1559787497
transform 1 0 1076 0 1 305
box -2 -3 26 103
use INVX1  _845_
timestamp 1559787497
transform -1 0 1116 0 1 305
box -2 -3 18 103
use INVX1  _1053_
timestamp 1559787497
transform 1 0 1116 0 1 305
box -2 -3 18 103
use BUFX2  BUFX2_insert17
timestamp 1559787497
transform 1 0 1132 0 1 305
box -2 -3 26 103
use OR2X2  _1016_
timestamp 1559787497
transform 1 0 1156 0 1 305
box -2 -3 34 103
use OR2X2  _1049_
timestamp 1559787497
transform 1 0 1188 0 1 305
box -2 -3 34 103
use NAND3X1  _1052_
timestamp 1559787497
transform -1 0 1252 0 1 305
box -2 -3 34 103
use NAND2X1  _1054_
timestamp 1559787497
transform -1 0 1276 0 1 305
box -2 -3 26 103
use NAND2X1  _1015_
timestamp 1559787497
transform -1 0 1300 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert19
timestamp 1559787497
transform -1 0 1324 0 1 305
box -2 -3 26 103
use NAND3X1  _1106_
timestamp 1559787497
transform 1 0 1324 0 1 305
box -2 -3 34 103
use NAND3X1  _1017_
timestamp 1559787497
transform 1 0 1356 0 1 305
box -2 -3 34 103
use NAND3X1  _1018_
timestamp 1559787497
transform -1 0 1420 0 1 305
box -2 -3 34 103
use NAND3X1  _1013_
timestamp 1559787497
transform 1 0 1420 0 1 305
box -2 -3 34 103
use INVX2  _1008_
timestamp 1559787497
transform -1 0 1468 0 1 305
box -2 -3 18 103
use FILL  FILL_4_1
timestamp 1559787497
transform 1 0 1468 0 1 305
box -2 -3 10 103
use INVX1  _1216_
timestamp 1559787497
transform 1 0 4 0 -1 305
box -2 -3 18 103
use NAND2X1  _1217_
timestamp 1559787497
transform -1 0 44 0 -1 305
box -2 -3 26 103
use OR2X2  _1215_
timestamp 1559787497
transform 1 0 44 0 -1 305
box -2 -3 34 103
use NAND3X1  _1218_
timestamp 1559787497
transform -1 0 108 0 -1 305
box -2 -3 34 103
use NAND3X1  _1223_
timestamp 1559787497
transform -1 0 140 0 -1 305
box -2 -3 34 103
use NAND3X1  _1310_
timestamp 1559787497
transform -1 0 172 0 -1 305
box -2 -3 34 103
use NAND3X1  _1262_
timestamp 1559787497
transform 1 0 172 0 -1 305
box -2 -3 34 103
use NAND3X1  _1261_
timestamp 1559787497
transform 1 0 204 0 -1 305
box -2 -3 34 103
use NAND2X1  _1270_
timestamp 1559787497
transform 1 0 236 0 -1 305
box -2 -3 26 103
use NAND3X1  _1305_
timestamp 1559787497
transform 1 0 260 0 -1 305
box -2 -3 34 103
use OR2X2  _1260_
timestamp 1559787497
transform -1 0 324 0 -1 305
box -2 -3 34 103
use OR2X2  _1302_
timestamp 1559787497
transform -1 0 356 0 -1 305
box -2 -3 34 103
use OR2X2  _804_
timestamp 1559787497
transform 1 0 356 0 -1 305
box -2 -3 34 103
use NAND2X1  _728_
timestamp 1559787497
transform 1 0 388 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert31
timestamp 1559787497
transform -1 0 436 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert33
timestamp 1559787497
transform 1 0 436 0 -1 305
box -2 -3 26 103
use NAND2X1  _719_
timestamp 1559787497
transform 1 0 460 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_0_0
timestamp 1559787497
transform -1 0 492 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1559787497
transform -1 0 500 0 -1 305
box -2 -3 10 103
use INVX1  _718_
timestamp 1559787497
transform -1 0 516 0 -1 305
box -2 -3 18 103
use NAND2X1  _758_
timestamp 1559787497
transform 1 0 516 0 -1 305
box -2 -3 26 103
use OR2X2  _762_
timestamp 1559787497
transform 1 0 540 0 -1 305
box -2 -3 34 103
use INVX1  _848_
timestamp 1559787497
transform 1 0 572 0 -1 305
box -2 -3 18 103
use NAND2X1  _849_
timestamp 1559787497
transform -1 0 612 0 -1 305
box -2 -3 26 103
use OR2X2  _931_
timestamp 1559787497
transform 1 0 612 0 -1 305
box -2 -3 34 103
use NAND2X1  _933_
timestamp 1559787497
transform 1 0 644 0 -1 305
box -2 -3 26 103
use INVX1  _932_
timestamp 1559787497
transform -1 0 684 0 -1 305
box -2 -3 18 103
use NAND3X1  _934_
timestamp 1559787497
transform -1 0 716 0 -1 305
box -2 -3 34 103
use INVX1  _1137_
timestamp 1559787497
transform 1 0 716 0 -1 305
box -2 -3 18 103
use OR2X2  _883_
timestamp 1559787497
transform 1 0 732 0 -1 305
box -2 -3 34 103
use NAND3X1  _939_
timestamp 1559787497
transform -1 0 796 0 -1 305
box -2 -3 34 103
use NAND3X1  _940_
timestamp 1559787497
transform -1 0 828 0 -1 305
box -2 -3 34 103
use NAND3X1  _901_
timestamp 1559787497
transform 1 0 828 0 -1 305
box -2 -3 34 103
use NAND3X1  _891_
timestamp 1559787497
transform 1 0 860 0 -1 305
box -2 -3 34 103
use NAND3X1  _886_
timestamp 1559787497
transform 1 0 892 0 -1 305
box -2 -3 34 103
use INVX1  _884_
timestamp 1559787497
transform 1 0 924 0 -1 305
box -2 -3 18 103
use NAND2X1  _885_
timestamp 1559787497
transform -1 0 964 0 -1 305
box -2 -3 26 103
use NAND3X1  _890_
timestamp 1559787497
transform 1 0 964 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1559787497
transform 1 0 996 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1559787497
transform 1 0 1004 0 -1 305
box -2 -3 10 103
use INVX1  _887_
timestamp 1559787497
transform 1 0 1012 0 -1 305
box -2 -3 18 103
use NAND2X1  _888_
timestamp 1559787497
transform -1 0 1052 0 -1 305
box -2 -3 26 103
use OR2X2  _889_
timestamp 1559787497
transform -1 0 1084 0 -1 305
box -2 -3 34 103
use INVX1  _1050_
timestamp 1559787497
transform 1 0 1084 0 -1 305
box -2 -3 18 103
use INVX1  _1092_
timestamp 1559787497
transform 1 0 1100 0 -1 305
box -2 -3 18 103
use NAND2X1  _1051_
timestamp 1559787497
transform -1 0 1140 0 -1 305
box -2 -3 26 103
use NAND2X1  _1093_
timestamp 1559787497
transform -1 0 1164 0 -1 305
box -2 -3 26 103
use NAND2X1  _1138_
timestamp 1559787497
transform 1 0 1164 0 -1 305
box -2 -3 26 103
use OR2X2  _1136_
timestamp 1559787497
transform 1 0 1188 0 -1 305
box -2 -3 34 103
use NAND3X1  _1139_
timestamp 1559787497
transform 1 0 1220 0 -1 305
box -2 -3 34 103
use OR2X2  _1094_
timestamp 1559787497
transform 1 0 1252 0 -1 305
box -2 -3 34 103
use NAND3X1  _1095_
timestamp 1559787497
transform 1 0 1284 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert16
timestamp 1559787497
transform 1 0 1316 0 -1 305
box -2 -3 26 103
use NAND3X1  _1105_
timestamp 1559787497
transform 1 0 1340 0 -1 305
box -2 -3 34 103
use NAND2X1  _1099_
timestamp 1559787497
transform 1 0 1372 0 -1 305
box -2 -3 26 103
use INVX1  _1098_
timestamp 1559787497
transform -1 0 1412 0 -1 305
box -2 -3 18 103
use NAND2X1  _1012_
timestamp 1559787497
transform 1 0 1412 0 -1 305
box -2 -3 26 103
use INVX1  _1011_
timestamp 1559787497
transform -1 0 1452 0 -1 305
box -2 -3 18 103
use FILL  FILL_3_1
timestamp 1559787497
transform -1 0 1460 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1559787497
transform -1 0 1468 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_3
timestamp 1559787497
transform -1 0 1476 0 -1 305
box -2 -3 10 103
use BUFX2  BUFX2_insert3
timestamp 1559787497
transform 1 0 4 0 1 105
box -2 -3 26 103
use OR2X2  _1221_
timestamp 1559787497
transform 1 0 28 0 1 105
box -2 -3 34 103
use NAND3X1  _1222_
timestamp 1559787497
transform -1 0 92 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert0
timestamp 1559787497
transform 1 0 92 0 1 105
box -2 -3 26 103
use NAND3X1  _1232_
timestamp 1559787497
transform -1 0 148 0 1 105
box -2 -3 34 103
use NAND3X1  _1257_
timestamp 1559787497
transform -1 0 180 0 1 105
box -2 -3 34 103
use OR2X2  _1254_
timestamp 1559787497
transform -1 0 212 0 1 105
box -2 -3 34 103
use NAND2X1  _1256_
timestamp 1559787497
transform 1 0 212 0 1 105
box -2 -3 26 103
use NAND3X1  _1227_
timestamp 1559787497
transform -1 0 268 0 1 105
box -2 -3 34 103
use OR2X2  _1224_
timestamp 1559787497
transform -1 0 300 0 1 105
box -2 -3 34 103
use OAI21X1  _1269_
timestamp 1559787497
transform -1 0 332 0 1 105
box -2 -3 34 103
use INVX1  _1255_
timestamp 1559787497
transform -1 0 348 0 1 105
box -2 -3 18 103
use OAI21X1  _810_
timestamp 1559787497
transform -1 0 380 0 1 105
box -2 -3 34 103
use INVX1  _808_
timestamp 1559787497
transform -1 0 396 0 1 105
box -2 -3 18 103
use INVX1  _727_
timestamp 1559787497
transform 1 0 396 0 1 105
box -2 -3 18 103
use INVX1  _1267_
timestamp 1559787497
transform -1 0 428 0 1 105
box -2 -3 18 103
use OR2X2  _726_
timestamp 1559787497
transform 1 0 428 0 1 105
box -2 -3 34 103
use INVX1  _769_
timestamp 1559787497
transform 1 0 460 0 1 105
box -2 -3 18 103
use FILL  FILL_1_0_0
timestamp 1559787497
transform 1 0 476 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1559787497
transform 1 0 484 0 1 105
box -2 -3 10 103
use OAI21X1  _771_
timestamp 1559787497
transform 1 0 492 0 1 105
box -2 -3 34 103
use INVX1  _757_
timestamp 1559787497
transform 1 0 524 0 1 105
box -2 -3 18 103
use OR2X2  _756_
timestamp 1559787497
transform 1 0 540 0 1 105
box -2 -3 34 103
use INVX1  _1140_
timestamp 1559787497
transform 1 0 572 0 1 105
box -2 -3 18 103
use OAI21X1  _1142_
timestamp 1559787497
transform 1 0 588 0 1 105
box -2 -3 34 103
use OR2X2  _970_
timestamp 1559787497
transform 1 0 620 0 1 105
box -2 -3 34 103
use INVX1  _971_
timestamp 1559787497
transform -1 0 668 0 1 105
box -2 -3 18 103
use NAND2X1  _972_
timestamp 1559787497
transform -1 0 692 0 1 105
box -2 -3 26 103
use NAND3X1  _973_
timestamp 1559787497
transform -1 0 724 0 1 105
box -2 -3 34 103
use NAND3X1  _978_
timestamp 1559787497
transform 1 0 724 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert26
timestamp 1559787497
transform -1 0 780 0 1 105
box -2 -3 26 103
use OR2X2  _892_
timestamp 1559787497
transform 1 0 780 0 1 105
box -2 -3 34 103
use NAND3X1  _895_
timestamp 1559787497
transform -1 0 844 0 1 105
box -2 -3 34 103
use NAND3X1  _900_
timestamp 1559787497
transform 1 0 844 0 1 105
box -2 -3 34 103
use NAND3X1  _930_
timestamp 1559787497
transform 1 0 876 0 1 105
box -2 -3 34 103
use NAND3X1  _929_
timestamp 1559787497
transform 1 0 908 0 1 105
box -2 -3 34 103
use OR2X2  _928_
timestamp 1559787497
transform -1 0 972 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert28
timestamp 1559787497
transform 1 0 972 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1559787497
transform 1 0 996 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1559787497
transform 1 0 1004 0 1 105
box -2 -3 10 103
use NAND3X1  _925_
timestamp 1559787497
transform 1 0 1012 0 1 105
box -2 -3 34 103
use OR2X2  _922_
timestamp 1559787497
transform -1 0 1076 0 1 105
box -2 -3 34 103
use INVX1  _1089_
timestamp 1559787497
transform 1 0 1076 0 1 105
box -2 -3 18 103
use NAND2X1  _1090_
timestamp 1559787497
transform -1 0 1116 0 1 105
box -2 -3 26 103
use OR2X2  _1088_
timestamp 1559787497
transform 1 0 1116 0 1 105
box -2 -3 34 103
use NAND3X1  _1091_
timestamp 1559787497
transform -1 0 1180 0 1 105
box -2 -3 34 103
use NAND2X1  _1143_
timestamp 1559787497
transform -1 0 1204 0 1 105
box -2 -3 26 103
use NAND3X1  _1144_
timestamp 1559787497
transform -1 0 1236 0 1 105
box -2 -3 34 103
use NAND3X1  _1066_
timestamp 1559787497
transform 1 0 1236 0 1 105
box -2 -3 34 103
use NAND3X1  _1096_
timestamp 1559787497
transform 1 0 1268 0 1 105
box -2 -3 34 103
use OR2X2  _1097_
timestamp 1559787497
transform 1 0 1300 0 1 105
box -2 -3 34 103
use NAND3X1  _1100_
timestamp 1559787497
transform 1 0 1332 0 1 105
box -2 -3 34 103
use INVX1  _1118_
timestamp 1559787497
transform 1 0 1364 0 1 105
box -2 -3 18 103
use INVX1  _990_
timestamp 1559787497
transform -1 0 1396 0 1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert6
timestamp 1559787497
transform -1 0 1420 0 1 105
box -2 -3 26 103
use BUFX2  _645_
timestamp 1559787497
transform 1 0 1420 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1559787497
transform 1 0 1444 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1559787497
transform 1 0 1452 0 1 105
box -2 -3 10 103
use FILL  FILL_2_3
timestamp 1559787497
transform 1 0 1460 0 1 105
box -2 -3 10 103
use FILL  FILL_2_4
timestamp 1559787497
transform 1 0 1468 0 1 105
box -2 -3 10 103
use INVX1  _1219_
timestamp 1559787497
transform 1 0 4 0 -1 105
box -2 -3 18 103
use NAND2X1  _1220_
timestamp 1559787497
transform -1 0 44 0 -1 105
box -2 -3 26 103
use NAND2X1  _1309_
timestamp 1559787497
transform 1 0 44 0 -1 105
box -2 -3 26 103
use OAI21X1  _1308_
timestamp 1559787497
transform -1 0 100 0 -1 105
box -2 -3 34 103
use NAND2X1  _1307_
timestamp 1559787497
transform 1 0 100 0 -1 105
box -2 -3 26 103
use NAND2X1  _1231_
timestamp 1559787497
transform 1 0 124 0 -1 105
box -2 -3 26 103
use INVX1  _1306_
timestamp 1559787497
transform -1 0 164 0 -1 105
box -2 -3 18 103
use NAND2X1  _1226_
timestamp 1559787497
transform 1 0 164 0 -1 105
box -2 -3 26 103
use INVX1  _1225_
timestamp 1559787497
transform -1 0 204 0 -1 105
box -2 -3 18 103
use NAND2X1  _1259_
timestamp 1559787497
transform 1 0 204 0 -1 105
box -2 -3 26 103
use INVX1  _1258_
timestamp 1559787497
transform -1 0 244 0 -1 105
box -2 -3 18 103
use OAI21X1  _1230_
timestamp 1559787497
transform -1 0 276 0 -1 105
box -2 -3 34 103
use NAND2X1  _1229_
timestamp 1559787497
transform 1 0 276 0 -1 105
box -2 -3 26 103
use NAND2X1  _1268_
timestamp 1559787497
transform 1 0 300 0 -1 105
box -2 -3 26 103
use INVX1  _1228_
timestamp 1559787497
transform -1 0 340 0 -1 105
box -2 -3 18 103
use NAND2X1  _809_
timestamp 1559787497
transform -1 0 364 0 -1 105
box -2 -3 26 103
use INVX1  _730_
timestamp 1559787497
transform 1 0 364 0 -1 105
box -2 -3 18 103
use OAI21X1  _732_
timestamp 1559787497
transform 1 0 380 0 -1 105
box -2 -3 34 103
use NAND2X1  _731_
timestamp 1559787497
transform -1 0 436 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert34
timestamp 1559787497
transform 1 0 436 0 -1 105
box -2 -3 26 103
use NAND2X1  _770_
timestamp 1559787497
transform 1 0 460 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1559787497
transform -1 0 492 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1559787497
transform -1 0 500 0 -1 105
box -2 -3 10 103
use NAND2X1  _936_
timestamp 1559787497
transform -1 0 524 0 -1 105
box -2 -3 26 103
use OAI21X1  _937_
timestamp 1559787497
transform -1 0 556 0 -1 105
box -2 -3 34 103
use INVX1  _935_
timestamp 1559787497
transform -1 0 572 0 -1 105
box -2 -3 18 103
use NAND2X1  _1102_
timestamp 1559787497
transform -1 0 596 0 -1 105
box -2 -3 26 103
use NAND2X1  _1141_
timestamp 1559787497
transform 1 0 596 0 -1 105
box -2 -3 26 103
use INVX1  _1101_
timestamp 1559787497
transform 1 0 620 0 -1 105
box -2 -3 18 103
use OAI21X1  _1103_
timestamp 1559787497
transform 1 0 636 0 -1 105
box -2 -3 34 103
use INVX1  _974_
timestamp 1559787497
transform 1 0 668 0 -1 105
box -2 -3 18 103
use OAI21X1  _976_
timestamp 1559787497
transform 1 0 684 0 -1 105
box -2 -3 34 103
use NAND2X1  _975_
timestamp 1559787497
transform -1 0 740 0 -1 105
box -2 -3 26 103
use NAND2X1  _977_
timestamp 1559787497
transform -1 0 764 0 -1 105
box -2 -3 26 103
use NAND2X1  _938_
timestamp 1559787497
transform -1 0 788 0 -1 105
box -2 -3 26 103
use INVX1  _893_
timestamp 1559787497
transform -1 0 804 0 -1 105
box -2 -3 18 103
use NAND2X1  _894_
timestamp 1559787497
transform -1 0 828 0 -1 105
box -2 -3 26 103
use NAND2X1  _899_
timestamp 1559787497
transform 1 0 828 0 -1 105
box -2 -3 26 103
use OAI21X1  _898_
timestamp 1559787497
transform -1 0 884 0 -1 105
box -2 -3 34 103
use INVX1  _896_
timestamp 1559787497
transform -1 0 900 0 -1 105
box -2 -3 18 103
use NAND2X1  _897_
timestamp 1559787497
transform 1 0 900 0 -1 105
box -2 -3 26 103
use NAND2X1  _927_
timestamp 1559787497
transform 1 0 924 0 -1 105
box -2 -3 26 103
use INVX1  _926_
timestamp 1559787497
transform -1 0 964 0 -1 105
box -2 -3 18 103
use INVX1  _1059_
timestamp 1559787497
transform 1 0 964 0 -1 105
box -2 -3 18 103
use FILL  FILL_0_1_0
timestamp 1559787497
transform 1 0 980 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1559787497
transform 1 0 988 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_insert27
timestamp 1559787497
transform 1 0 996 0 -1 105
box -2 -3 26 103
use NAND2X1  _924_
timestamp 1559787497
transform 1 0 1020 0 -1 105
box -2 -3 26 103
use INVX1  _923_
timestamp 1559787497
transform -1 0 1060 0 -1 105
box -2 -3 18 103
use INVX1  _1062_
timestamp 1559787497
transform 1 0 1060 0 -1 105
box -2 -3 18 103
use NAND2X1  _1063_
timestamp 1559787497
transform -1 0 1100 0 -1 105
box -2 -3 26 103
use OAI21X1  _1064_
timestamp 1559787497
transform 1 0 1100 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert15
timestamp 1559787497
transform -1 0 1156 0 -1 105
box -2 -3 26 103
use NAND2X1  _1060_
timestamp 1559787497
transform 1 0 1156 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert18
timestamp 1559787497
transform -1 0 1204 0 -1 105
box -2 -3 26 103
use NAND2X1  _1065_
timestamp 1559787497
transform -1 0 1228 0 -1 105
box -2 -3 26 103
use NAND3X1  _1061_
timestamp 1559787497
transform -1 0 1260 0 -1 105
box -2 -3 34 103
use OR2X2  _1058_
timestamp 1559787497
transform -1 0 1292 0 -1 105
box -2 -3 34 103
use NAND2X1  _1104_
timestamp 1559787497
transform -1 0 1316 0 -1 105
box -2 -3 26 103
use INVX1  _1112_
timestamp 1559787497
transform -1 0 1332 0 -1 105
box -2 -3 18 103
use NAND3X1  _1028_
timestamp 1559787497
transform -1 0 1364 0 -1 105
box -2 -3 34 103
use OR2X2  _1069_
timestamp 1559787497
transform 1 0 1364 0 -1 105
box -2 -3 34 103
use OR2X2  _998_
timestamp 1559787497
transform -1 0 1428 0 -1 105
box -2 -3 34 103
use OR2X2  _1010_
timestamp 1559787497
transform -1 0 1460 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1559787497
transform -1 0 1468 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1559787497
transform -1 0 1476 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 472 -30 488 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 984 -30 1000 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 CLK
port 2 nsew
flabel metal2 s 718 -22 722 -18 7 FreeSans 24 270 0 0 DATA_A[31]
port 3 nsew
flabel metal2 s 1006 -22 1010 -18 7 FreeSans 24 270 0 0 DATA_A[30]
port 4 nsew
flabel metal2 s 918 -22 922 -18 7 FreeSans 24 270 0 0 DATA_A[29]
port 5 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 DATA_A[28]
port 6 nsew
flabel metal3 s -26 538 -22 542 7 FreeSans 24 0 0 0 DATA_A[27]
port 7 nsew
flabel metal2 s 494 -22 498 -18 7 FreeSans 24 270 0 0 DATA_A[26]
port 8 nsew
flabel metal3 s -26 88 -22 92 7 FreeSans 24 0 0 0 DATA_A[25]
port 9 nsew
flabel metal3 s -26 348 -22 352 7 FreeSans 24 0 0 0 DATA_A[24]
port 10 nsew
flabel metal2 s 654 -22 658 -18 7 FreeSans 24 270 0 0 DATA_A[23]
port 11 nsew
flabel metal2 s 1046 -22 1050 -18 7 FreeSans 24 270 0 0 DATA_A[22]
port 12 nsew
flabel metal2 s 798 -22 802 -18 7 FreeSans 24 270 0 0 DATA_A[21]
port 13 nsew
flabel metal3 s -26 748 -22 752 7 FreeSans 24 0 0 0 DATA_A[20]
port 14 nsew
flabel metal3 s -26 728 -22 732 7 FreeSans 24 0 0 0 DATA_A[19]
port 15 nsew
flabel metal3 s 1502 358 1506 362 3 FreeSans 24 0 0 0 DATA_A[18]
port 16 nsew
flabel metal3 s -26 288 -22 292 7 FreeSans 24 0 0 0 DATA_A[17]
port 17 nsew
flabel metal3 s 1502 278 1506 282 3 FreeSans 24 0 0 0 DATA_A[16]
port 18 nsew
flabel metal2 s 670 -22 674 -18 7 FreeSans 24 270 0 0 DATA_A[15]
port 19 nsew
flabel metal2 s 958 -22 962 -18 7 FreeSans 24 270 0 0 DATA_A[14]
port 20 nsew
flabel metal2 s 886 -22 890 -18 7 FreeSans 24 270 0 0 DATA_A[13]
port 21 nsew
flabel metal3 s -26 488 -22 492 7 FreeSans 24 0 0 0 DATA_A[12]
port 22 nsew
flabel metal3 s -26 558 -22 562 7 FreeSans 24 0 0 0 DATA_A[11]
port 23 nsew
flabel metal2 s 558 -22 562 -18 7 FreeSans 24 270 0 0 DATA_A[10]
port 24 nsew
flabel metal3 s -26 168 -22 172 7 FreeSans 24 0 0 0 DATA_A[9]
port 25 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 DATA_A[8]
port 26 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 DATA_A[7]
port 27 nsew
flabel metal2 s 1070 -22 1074 -18 7 FreeSans 24 270 0 0 DATA_A[6]
port 28 nsew
flabel metal2 s 1270 -22 1274 -18 7 FreeSans 24 270 0 0 DATA_A[5]
port 29 nsew
flabel metal3 s -26 688 -22 692 7 FreeSans 24 0 0 0 DATA_A[4]
port 30 nsew
flabel metal3 s -26 788 -22 792 7 FreeSans 24 0 0 0 DATA_A[3]
port 31 nsew
flabel metal2 s 1318 -22 1322 -18 7 FreeSans 24 270 0 0 DATA_A[2]
port 32 nsew
flabel metal3 s -26 268 -22 272 7 FreeSans 24 0 0 0 DATA_A[1]
port 33 nsew
flabel metal3 s 1502 108 1506 112 3 FreeSans 24 0 0 0 DATA_A[0]
port 34 nsew
flabel metal2 s 630 1438 634 1442 3 FreeSans 24 90 0 0 DATA_B[31]
port 35 nsew
flabel metal2 s 422 1438 426 1442 3 FreeSans 24 90 0 0 DATA_B[30]
port 36 nsew
flabel metal2 s 694 1438 698 1442 3 FreeSans 24 90 0 0 DATA_B[29]
port 37 nsew
flabel metal2 s 742 1438 746 1442 3 FreeSans 24 90 0 0 DATA_B[28]
port 38 nsew
flabel metal3 s 1502 1048 1506 1052 3 FreeSans 24 0 0 0 DATA_B[27]
port 39 nsew
flabel metal3 s 1502 888 1506 892 3 FreeSans 24 0 0 0 DATA_B[26]
port 40 nsew
flabel metal2 s 342 1438 346 1442 3 FreeSans 24 90 0 0 DATA_B[25]
port 41 nsew
flabel metal3 s 1502 988 1506 992 3 FreeSans 24 0 0 0 DATA_B[24]
port 42 nsew
flabel metal3 s 1502 148 1506 152 3 FreeSans 24 0 0 0 DATA_B[23]
port 43 nsew
flabel metal2 s 854 1438 858 1442 3 FreeSans 24 90 0 0 DATA_B[22]
port 44 nsew
flabel metal2 s 166 1438 170 1442 3 FreeSans 24 90 0 0 DATA_B[21]
port 45 nsew
flabel metal3 s 1502 1138 1506 1142 3 FreeSans 24 0 0 0 DATA_B[20]
port 46 nsew
flabel metal2 s 86 1438 90 1442 3 FreeSans 24 90 0 0 DATA_B[19]
port 47 nsew
flabel metal3 s 1502 928 1506 932 3 FreeSans 24 0 0 0 DATA_B[18]
port 48 nsew
flabel metal3 s 1502 1008 1506 1012 3 FreeSans 24 0 0 0 DATA_B[17]
port 49 nsew
flabel metal3 s 1502 128 1506 132 3 FreeSans 24 0 0 0 DATA_B[16]
port 50 nsew
flabel metal3 s -26 1328 -22 1332 7 FreeSans 24 0 0 0 DATA_B[15]
port 51 nsew
flabel metal2 s 942 1438 946 1442 3 FreeSans 24 90 0 0 DATA_B[14]
port 52 nsew
flabel metal2 s 718 1438 722 1442 3 FreeSans 24 90 0 0 DATA_B[13]
port 53 nsew
flabel metal2 s 758 1438 762 1442 3 FreeSans 24 90 0 0 DATA_B[12]
port 54 nsew
flabel metal3 s 1502 1158 1506 1162 3 FreeSans 24 0 0 0 DATA_B[11]
port 55 nsew
flabel metal3 s 1502 848 1506 852 3 FreeSans 24 0 0 0 DATA_B[10]
port 56 nsew
flabel metal3 s 1502 1068 1506 1072 3 FreeSans 24 0 0 0 DATA_B[9]
port 57 nsew
flabel metal3 s 1502 968 1506 972 3 FreeSans 24 0 0 0 DATA_B[8]
port 58 nsew
flabel metal2 s 1366 1438 1370 1442 3 FreeSans 24 90 0 0 DATA_B[7]
port 59 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 DATA_B[6]
port 60 nsew
flabel metal2 s 590 1438 594 1442 3 FreeSans 24 90 0 0 DATA_B[5]
port 61 nsew
flabel metal3 s 1502 68 1506 72 3 FreeSans 24 0 0 0 DATA_B[4]
port 62 nsew
flabel metal3 s -26 1268 -22 1272 7 FreeSans 24 0 0 0 DATA_B[3]
port 63 nsew
flabel metal3 s 1502 88 1506 92 3 FreeSans 24 0 0 0 DATA_B[2]
port 64 nsew
flabel metal3 s 1502 948 1506 952 3 FreeSans 24 0 0 0 DATA_B[1]
port 65 nsew
flabel metal3 s 1502 1088 1506 1092 3 FreeSans 24 0 0 0 DATA_B[0]
port 66 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 NIBBLE_OUT[15]
port 67 nsew
flabel metal3 s -26 828 -22 832 7 FreeSans 24 0 0 0 NIBBLE_OUT[14]
port 68 nsew
flabel metal3 s -26 868 -22 872 7 FreeSans 24 0 0 0 NIBBLE_OUT[13]
port 69 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 NIBBLE_OUT[12]
port 70 nsew
flabel metal3 s 1502 778 1506 782 3 FreeSans 24 0 0 0 NIBBLE_OUT[11]
port 71 nsew
flabel metal3 s 1502 728 1506 732 3 FreeSans 24 0 0 0 NIBBLE_OUT[10]
port 72 nsew
flabel metal3 s 1502 648 1506 652 3 FreeSans 24 0 0 0 NIBBLE_OUT[9]
port 73 nsew
flabel metal3 s 1502 168 1506 172 3 FreeSans 24 0 0 0 NIBBLE_OUT[8]
port 74 nsew
flabel metal2 s 934 -22 938 -18 7 FreeSans 24 270 0 0 NIBBLE_OUT[7]
port 75 nsew
flabel metal3 s 1502 668 1506 672 3 FreeSans 24 0 0 0 NIBBLE_OUT[6]
port 76 nsew
flabel metal3 s -26 808 -22 812 7 FreeSans 24 0 0 0 NIBBLE_OUT[5]
port 77 nsew
flabel metal3 s 1502 798 1506 802 3 FreeSans 24 0 0 0 NIBBLE_OUT[4]
port 78 nsew
flabel metal3 s 1502 708 1506 712 3 FreeSans 24 0 0 0 NIBBLE_OUT[3]
port 79 nsew
flabel metal3 s 1502 688 1506 692 3 FreeSans 24 0 0 0 NIBBLE_OUT[2]
port 80 nsew
flabel metal3 s -26 888 -22 892 7 FreeSans 24 0 0 0 NIBBLE_OUT[1]
port 81 nsew
flabel metal3 s -26 848 -22 852 7 FreeSans 24 0 0 0 NIBBLE_OUT[0]
port 82 nsew
flabel metal3 s -26 708 -22 712 7 FreeSans 24 0 0 0 RESET_L
port 83 nsew
flabel metal3 s -26 378 -22 382 7 FreeSans 24 0 0 0 SEL[3]
port 84 nsew
flabel metal3 s 1502 48 1506 52 3 FreeSans 24 270 0 0 SEL[2]
port 85 nsew
flabel metal2 s 814 -22 818 -18 7 FreeSans 24 270 0 0 SEL[1]
port 86 nsew
flabel metal3 s -26 668 -22 672 7 FreeSans 24 0 0 0 SEL[0]
port 87 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 sel_A[11]
port 88 nsew
flabel metal3 s -26 68 -22 72 7 FreeSans 24 0 0 0 sel_A[10]
port 89 nsew
flabel metal3 s -26 578 -22 582 7 FreeSans 24 0 0 0 sel_A[9]
port 90 nsew
flabel metal2 s 1142 -22 1146 -18 7 FreeSans 24 270 0 0 sel_A[8]
port 91 nsew
flabel metal2 s 1302 -22 1306 -18 7 FreeSans 24 270 0 0 sel_A[7]
port 92 nsew
flabel metal3 s 1502 338 1506 342 3 FreeSans 24 0 0 0 sel_A[6]
port 93 nsew
flabel metal2 s 1022 -22 1026 -18 7 FreeSans 24 270 0 0 sel_A[5]
port 94 nsew
flabel metal2 s 774 -22 778 -18 7 FreeSans 24 270 0 0 sel_A[4]
port 95 nsew
flabel metal2 s 750 -22 754 -18 7 FreeSans 24 270 0 0 sel_A[3]
port 96 nsew
flabel metal2 s 454 -22 458 -18 7 FreeSans 24 270 0 0 sel_A[2]
port 97 nsew
flabel metal3 s -26 768 -22 772 7 FreeSans 24 0 0 0 sel_A[1]
port 98 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 sel_A[0]
port 99 nsew
flabel metal2 s 238 1438 242 1442 3 FreeSans 24 90 0 0 sel_B[11]
port 100 nsew
flabel metal3 s -26 1308 -22 1312 7 FreeSans 24 0 0 0 sel_B[10]
port 101 nsew
flabel metal3 s -26 1168 -22 1172 7 FreeSans 24 0 0 0 sel_B[9]
port 102 nsew
flabel metal3 s 1502 758 1506 762 3 FreeSans 24 0 0 0 sel_B[8]
port 103 nsew
flabel metal2 s 1350 1438 1354 1442 3 FreeSans 24 90 0 0 sel_B[7]
port 104 nsew
flabel metal3 s 1502 1248 1506 1252 3 FreeSans 24 0 0 0 sel_B[6]
port 105 nsew
flabel metal2 s 542 1438 546 1442 3 FreeSans 24 90 0 0 sel_B[5]
port 106 nsew
flabel metal2 s 654 1438 658 1442 3 FreeSans 24 90 0 0 sel_B[4]
port 107 nsew
flabel metal2 s 670 1438 674 1442 3 FreeSans 24 90 0 0 sel_B[3]
port 108 nsew
flabel metal2 s 918 1438 922 1442 3 FreeSans 24 90 0 0 sel_B[2]
port 109 nsew
flabel metal2 s 894 1438 898 1442 3 FreeSans 24 90 0 0 sel_B[1]
port 110 nsew
flabel metal2 s 878 1438 882 1442 3 FreeSans 24 90 0 0 sel_B[0]
port 111 nsew
<< end >>
