* NGSPICE file created from selector4.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

.subckt selector4 vdd gnd CLK DATA_A[31] DATA_A[30] DATA_A[29] DATA_A[28] DATA_A[27]
+ DATA_A[26] DATA_A[25] DATA_A[24] DATA_A[23] DATA_A[22] DATA_A[21] DATA_A[20] DATA_A[19]
+ DATA_A[18] DATA_A[17] DATA_A[16] DATA_A[15] DATA_A[14] DATA_A[13] DATA_A[12] DATA_A[11]
+ DATA_A[10] DATA_A[9] DATA_A[8] DATA_A[7] DATA_A[6] DATA_A[5] DATA_A[4] DATA_A[3]
+ DATA_A[2] DATA_A[1] DATA_A[0] DATA_B[31] DATA_B[30] DATA_B[29] DATA_B[28] DATA_B[27]
+ DATA_B[26] DATA_B[25] DATA_B[24] DATA_B[23] DATA_B[22] DATA_B[21] DATA_B[20] DATA_B[19]
+ DATA_B[18] DATA_B[17] DATA_B[16] DATA_B[15] DATA_B[14] DATA_B[13] DATA_B[12] DATA_B[11]
+ DATA_B[10] DATA_B[9] DATA_B[8] DATA_B[7] DATA_B[6] DATA_B[5] DATA_B[4] DATA_B[3]
+ DATA_B[2] DATA_B[1] DATA_B[0] NIBBLE_OUT[15] NIBBLE_OUT[14] NIBBLE_OUT[13] NIBBLE_OUT[12]
+ NIBBLE_OUT[11] NIBBLE_OUT[10] NIBBLE_OUT[9] NIBBLE_OUT[8] NIBBLE_OUT[7] NIBBLE_OUT[6]
+ NIBBLE_OUT[5] NIBBLE_OUT[4] NIBBLE_OUT[3] NIBBLE_OUT[2] NIBBLE_OUT[1] NIBBLE_OUT[0]
+ RESET_L SEL[3] SEL[2] SEL[1] SEL[0] sel_A[11] sel_A[10] sel_A[9] sel_A[8] sel_A[7]
+ sel_A[6] sel_A[5] sel_A[4] sel_A[3] sel_A[2] sel_A[1] sel_A[0] sel_B[11] sel_B[10]
+ sel_B[9] sel_B[8] sel_B[7] sel_B[6] sel_B[5] sel_B[4] sel_B[3] sel_B[2] sel_B[1]
+ sel_B[0]
X_668_ _662_/A _668_/B gnd _668_/Y vdd NAND2X1
X_1017_ sel_B[7] _1017_/B _1017_/C gnd _1017_/Y vdd NAND3X1
X_888_ _922_/A _887_/Y gnd _890_/C vdd NAND2X1
X_1237_ _1235_/A _1236_/Y gnd _1238_/C vdd NAND2X1
X_1118_ DATA_A[23] gnd _1118_/Y vdd INVX1
X_769_ DATA_B[10] gnd _771_/A vdd INVX1
X_989_ DATA_A[0] _991_/A gnd _992_/B vdd OR2X2
X_650_ _650_/A gnd NIBBLE_OUT[13] vdd BUFX2
XFILL_1_1_0 gnd vdd FILL
X_870_ _828_/A DATA_A[9] gnd _870_/Y vdd OR2X2
X_1219_ DATA_B[25] gnd _1219_/Y vdd INVX1
XFILL_9_1 gnd vdd FILL
X_751_ _751_/A DATA_A[30] gnd _752_/C vdd NAND2X1
X_1100_ _1091_/A _1097_/Y _1100_/C gnd _1100_/Y vdd NAND3X1
XFILL_8_1_0 gnd vdd FILL
X_971_ DATA_B[23] gnd _971_/Y vdd INVX1
X_852_ _939_/A _852_/B _851_/Y gnd _862_/B vdd NAND3X1
X_1201_ _1169_/A _1200_/Y gnd _1201_/Y vdd NAND2X1
X_1082_ DATA_A[14] gnd _1084_/A vdd INVX1
X_733_ sel_B[1] _733_/B gnd _734_/C vdd NAND2X1
X_953_ _957_/B _952_/Y gnd _953_/Y vdd NAND2X1
XBUFX2_insert9 sel_B[8] gnd _1058_/A vdd BUFX2
X_1302_ _1302_/A DATA_B[7] gnd _1302_/Y vdd OR2X2
X_834_ _828_/A _833_/Y gnd _834_/Y vdd NAND2X1
X_1183_ sel_B[10] _1182_/Y _1183_/C gnd _1184_/C vdd NAND3X1
X_715_ sel_A[0] _715_/B _715_/C gnd _716_/C vdd NAND3X1
X_1064_ _1064_/A _1133_/A _1064_/C gnd _1065_/B vdd OAI21X1
X_1284_ DATA_A[23] gnd _1284_/Y vdd INVX1
X_935_ DATA_B[10] gnd _935_/Y vdd INVX1
XFILL_1_1_1 gnd vdd FILL
X_816_ _638_/A CLK _816_/D gnd vdd DFFPOSX1
X_1165_ DATA_A[20] gnd _1165_/Y vdd INVX1
X_1046_ sel_A[7] _1046_/B gnd _1047_/C vdd NAND2X1
X_697_ _697_/A _697_/B _653_/Y gnd _815_/D vdd AOI21X1
X_917_ _823_/B DATA_A[30] gnd _918_/C vdd NAND2X1
XFILL_8_1_1 gnd vdd FILL
XBUFX2_insert10 sel_B[5] gnd _853_/A vdd BUFX2
X_1266_ _1188_/A _1266_/B _1266_/C gnd _1271_/B vdd NAND3X1
X_798_ _759_/A _795_/Y _798_/C gnd _803_/B vdd NAND3X1
X_1147_ _645_/A CLK _1147_/D gnd vdd DFFPOSX1
X_679_ DATA_B[16] gnd _679_/Y vdd INVX1
X_1028_ SEL[2] _1028_/B _1028_/C gnd _1029_/B vdd NAND3X1
X_899_ sel_B[4] _898_/Y gnd _900_/C vdd NAND2X1
X_1248_ DATA_A[14] gnd _1248_/Y vdd INVX1
X_780_ DATA_A[27] gnd _780_/Y vdd INVX1
X_1129_ _1133_/A _1128_/Y gnd _1130_/C vdd NAND2X1
X_661_ DATA_A[24] gnd _661_/Y vdd INVX1
X_1010_ DATA_B[0] _1019_/A gnd _1013_/B vdd OR2X2
X_881_ sel_A[3] _881_/B _881_/C gnd _882_/C vdd NAND3X1
X_1230_ _1230_/A _1304_/A _1230_/C gnd _1231_/B vdd OAI21X1
X_762_ _758_/A DATA_B[14] gnd _762_/Y vdd OR2X2
X_1111_ _992_/A _1111_/B _1111_/C gnd _1116_/B vdd NAND3X1
X_643_ _983_/Q gnd NIBBLE_OUT[6] vdd BUFX2
X_982_ _982_/Q CLK _982_/D gnd vdd DFFPOSX1
X_863_ _841_/Y _863_/B _980_/C gnd _863_/Y vdd AOI21X1
X_1212_ sel_A[10] _1212_/B gnd _1213_/C vdd NAND2X1
XBUFX2_insert11 sel_B[5] gnd _963_/A vdd BUFX2
X_744_ sel_A[1] _743_/Y _744_/C gnd _744_/Y vdd NAND3X1
XFILL_13_1 gnd vdd FILL
X_1093_ _1094_/A _1093_/B gnd _1095_/C vdd NAND2X1
X_964_ _856_/A _961_/Y _964_/C gnd _964_/Y vdd NAND3X1
X_1313_ _649_/A CLK _1195_/Y gnd vdd DFFPOSX1
X_845_ DATA_B[16] gnd _845_/Y vdd INVX1
X_1194_ SEL[3] _1194_/B _1194_/C gnd _1195_/B vdd NAND3X1
X_726_ _801_/A DATA_B[5] gnd _726_/Y vdd OR2X2
X_1075_ _1075_/A DATA_A[10] gnd _1076_/B vdd OR2X2
X_946_ DATA_A[27] gnd _946_/Y vdd INVX1
X_1295_ _1293_/A _1295_/B gnd _1296_/C vdd NAND2X1
X_827_ DATA_A[24] gnd _827_/Y vdd INVX1
X_1176_ DATA_B[0] _1187_/A gnd _1176_/Y vdd OR2X2
X_708_ DATA_A[21] gnd _708_/Y vdd INVX1
X_1057_ _1018_/A _1057_/B _1057_/C gnd _1067_/B vdd NAND3X1
X_928_ _853_/A DATA_B[14] gnd _928_/Y vdd OR2X2
X_1277_ _1158_/A _1277_/B _1276_/Y gnd _1277_/Y vdd NAND3X1
XFILL_4_0_0 gnd vdd FILL
X_1158_ _1158_/A _1158_/B _1157_/Y gnd _1163_/B vdd NAND3X1
X_809_ _795_/A DATA_B[31] gnd _810_/C vdd NAND2X1
X_690_ _759_/A _690_/B _690_/C gnd _695_/B vdd NAND3X1
X_1039_ _1030_/A DATA_A[5] gnd _1042_/B vdd OR2X2
XFILL_13_2 gnd vdd FILL
XBUFX2_insert12 sel_B[5] gnd _849_/A vdd BUFX2
X_910_ sel_A[4] _909_/Y _910_/C gnd _910_/Y vdd NAND3X1
X_1259_ _1191_/B _1259_/B gnd _1261_/C vdd NAND2X1
X_791_ _789_/Y _751_/A _791_/C gnd _791_/Y vdd OAI21X1
X_1140_ DATA_B[15] gnd _1142_/A vdd INVX1
X_672_ _670_/Y _662_/A _672_/C gnd _672_/Y vdd OAI21X1
X_1021_ _1019_/A _1021_/B gnd _1022_/C vdd NAND2X1
X_892_ _963_/A DATA_B[5] gnd _892_/Y vdd OR2X2
X_1241_ _1160_/A DATA_A[10] gnd _1242_/B vdd OR2X2
X_1122_ _1123_/B DATA_A[31] gnd _1123_/C vdd NAND2X1
X_773_ _773_/A _768_/Y _772_/Y gnd _774_/C vdd NAND3X1
X_993_ DATA_A[24] gnd _993_/Y vdd INVX1
X_654_ SEL[0] gnd _755_/A vdd INVX2
X_1003_ _1074_/A DATA_A[28] gnd _1004_/C vdd NAND2X1
X_874_ DATA_A[21] gnd _875_/B vdd INVX1
X_1223_ _1271_/A _1223_/B _1223_/C gnd _1233_/B vdd NAND3X1
XFILL_4_0_1 gnd vdd FILL
X_755_ _755_/A _745_/Y _755_/C gnd _775_/A vdd NAND3X1
X_1104_ sel_B[7] _1104_/B gnd _1105_/C vdd NAND2X1
X_975_ _963_/A DATA_B[31] gnd _975_/Y vdd NAND2X1
XFILL_13_3 gnd vdd FILL
XBUFX2_insert13 sel_B[5] gnd _922_/A vdd BUFX2
X_856_ _856_/A _853_/Y _855_/Y gnd _861_/B vdd NAND3X1
X_1205_ _1250_/B DATA_A[5] gnd _1205_/Y vdd OR2X2
X_1086_ sel_A[6] _1086_/B _1086_/C gnd _1087_/C vdd NAND3X1
X_737_ _737_/A DATA_A[2] gnd _737_/Y vdd OR2X2
X_957_ _955_/Y _957_/B _957_/C gnd _957_/Y vdd OAI21X1
X_1306_ DATA_B[15] gnd _1308_/A vdd INVX1
X_838_ _836_/Y _944_/A _838_/C gnd _838_/Y vdd OAI21X1
X_1187_ _1187_/A _1187_/B gnd _1187_/Y vdd NAND2X1
X_719_ _758_/A _718_/Y gnd _720_/C vdd NAND2X1
X_1068_ _1048_/Y _1068_/B _985_/Y gnd _1068_/Y vdd AOI21X1
XFILL_11_0_0 gnd vdd FILL
X_1288_ _1250_/B DATA_A[31] gnd _1289_/C vdd NAND2X1
X_939_ _939_/A _934_/Y _938_/Y gnd _940_/C vdd NAND3X1
X_820_ SEL[1] gnd _841_/A vdd INVX2
X_1169_ _1169_/A DATA_A[28] gnd _1169_/Y vdd NAND2X1
X_701_ _669_/A _698_/Y _701_/C gnd _706_/B vdd NAND3X1
X_1050_ DATA_B[17] gnd _1051_/B vdd INVX1
X_921_ _841_/A _911_/Y _920_/Y gnd _941_/A vdd NAND3X1
X_1270_ sel_B[10] _1270_/B gnd _1271_/C vdd NAND2X1
XFILL_5_1_0 gnd vdd FILL
XBUFX2_insert14 sel_B[5] gnd _972_/A vdd BUFX2
X_802_ sel_B[1] _801_/Y _800_/Y gnd _802_/Y vdd NAND3X1
X_1151_ RESET_L gnd _1195_/C vdd INVX2
X_683_ _801_/A _682_/Y gnd _683_/Y vdd NAND2X1
X_1032_ _1075_/A _1032_/B gnd _1033_/C vdd NAND2X1
X_903_ _823_/B DATA_A[2] gnd _903_/Y vdd OR2X2
X_1252_ sel_A[9] _1252_/B _1252_/C gnd _1253_/C vdd NAND3X1
X_784_ _665_/A _784_/B _783_/Y gnd _794_/B vdd NAND3X1
X_1133_ _1133_/A DATA_B[11] gnd _1134_/B vdd OR2X2
X_665_ _665_/A _660_/Y _664_/Y gnd _665_/Y vdd NAND3X1
X_1014_ DATA_B[24] gnd _1014_/Y vdd INVX1
XFILL_11_0_1 gnd vdd FILL
X_885_ _849_/A _884_/Y gnd _885_/Y vdd NAND2X1
X_1234_ _1214_/Y _1234_/B _1195_/C gnd _1314_/D vdd AOI21X1
X_1115_ sel_A[7] _1115_/B _1115_/C gnd _1116_/C vdd NAND3X1
X_766_ DATA_B[18] gnd _767_/B vdd INVX1
X_647_ _647_/A gnd NIBBLE_OUT[10] vdd BUFX2
X_986_ SEL[2] gnd _986_/Y vdd INVX2
X_867_ _835_/A _864_/Y _866_/Y gnd _867_/Y vdd NAND3X1
X_1216_ DATA_B[17] gnd _1217_/B vdd INVX1
X_748_ _737_/A _747_/Y gnd _748_/Y vdd NAND2X1
XBUFX2_insert15 sel_A[8] gnd _1075_/A vdd BUFX2
XFILL_5_1_1 gnd vdd FILL
X_1097_ _1016_/A DATA_B[2] gnd _1097_/Y vdd OR2X2
X_968_ sel_B[4] _968_/B _968_/C gnd _969_/C vdd NAND3X1
X_849_ _849_/A _848_/Y gnd _849_/Y vdd NAND2X1
X_1198_ _1235_/A _1197_/Y gnd _1198_/Y vdd NAND2X1
X_1079_ DATA_A[22] gnd _1079_/Y vdd INVX1
X_730_ DATA_B[13] gnd _732_/A vdd INVX1
X_950_ _831_/A _950_/B _950_/C gnd _950_/Y vdd NAND3X1
X_1299_ _1302_/A DATA_B[11] gnd _1300_/B vdd OR2X2
X_831_ _831_/A _826_/Y _830_/Y gnd _831_/Y vdd NAND3X1
X_1180_ DATA_B[24] gnd _1181_/B vdd INVX1
X_712_ _704_/A DATA_A[29] gnd _713_/C vdd NAND2X1
X_1061_ _1091_/A _1058_/Y _1061_/C gnd _1066_/B vdd NAND3X1
XFILL_12_1_0 gnd vdd FILL
X_932_ DATA_B[18] gnd _932_/Y vdd INVX1
X_1281_ sel_A[10] _1280_/Y _1281_/C gnd _1281_/Y vdd NAND3X1
X_1162_ sel_A[10] _1162_/B _1162_/C gnd _1163_/C vdd NAND3X1
X_813_ SEL[0] _803_/Y _813_/C gnd _814_/B vdd NAND3X1
X_694_ sel_B[1] _694_/B gnd _695_/C vdd NAND2X1
X_1043_ DATA_A[13] gnd _1045_/A vdd INVX1
XBUFX2_insert16 sel_A[8] gnd _1123_/B vdd BUFX2
X_914_ _957_/B _913_/Y gnd _914_/Y vdd NAND2X1
X_1263_ _1187_/A DATA_B[2] gnd _1266_/B vdd OR2X2
X_795_ _795_/A DATA_B[3] gnd _795_/Y vdd OR2X2
X_1144_ sel_B[6] _1144_/B _1144_/C gnd _1145_/C vdd NAND3X1
X_676_ sel_B[0] gnd _773_/A vdd INVX2
X_1025_ _1025_/A _1094_/A _1025_/C gnd _1026_/B vdd OAI21X1
X_896_ DATA_B[13] gnd _896_/Y vdd INVX1
X_1245_ DATA_A[22] gnd _1245_/Y vdd INVX1
X_777_ DATA_A[19] gnd _778_/B vdd INVX1
X_1126_ _986_/Y _1116_/Y _1126_/C gnd _1146_/A vdd NAND3X1
X_658_ DATA_A[16] gnd _658_/Y vdd INVX1
X_997_ _997_/A _997_/B _997_/C gnd _997_/Y vdd NAND3X1
X_1007_ _986_/Y _997_/Y _1007_/C gnd _1007_/Y vdd NAND3X1
X_878_ _944_/A DATA_A[29] gnd _878_/Y vdd NAND2X1
XFILL_12_1_1 gnd vdd FILL
X_1227_ _1188_/A _1227_/B _1227_/C gnd _1232_/B vdd NAND3X1
X_759_ _759_/A _759_/B _758_/Y gnd _764_/B vdd NAND3X1
X_1108_ _1030_/A DATA_A[3] gnd _1111_/B vdd OR2X2
XFILL_1_0_0 gnd vdd FILL
X_640_ _818_/Q gnd NIBBLE_OUT[3] vdd BUFX2
X_979_ SEL[1] _969_/Y _979_/C gnd _980_/B vdd NAND3X1
X_860_ sel_B[4] _860_/B gnd _861_/C vdd NAND2X1
XBUFX2_insert17 sel_A[8] gnd _991_/A vdd BUFX2
X_1209_ DATA_A[13] gnd _1211_/A vdd INVX1
X_741_ DATA_A[26] gnd _742_/B vdd INVX1
X_1090_ _1019_/A _1090_/B gnd _1091_/C vdd NAND2X1
XFILL_8_0_0 gnd vdd FILL
X_961_ _849_/A DATA_B[3] gnd _961_/Y vdd OR2X2
X_1310_ sel_B[9] _1310_/B _1310_/C gnd _1311_/C vdd NAND3X1
X_1191_ _1191_/A _1191_/B _1191_/C gnd _1192_/B vdd OAI21X1
X_842_ sel_B[3] gnd _939_/A vdd INVX2
X_723_ _723_/A DATA_B[9] gnd _724_/B vdd OR2X2
X_1072_ _992_/A _1072_/B _1072_/C gnd _1077_/B vdd NAND3X1
X_943_ DATA_A[19] gnd _943_/Y vdd INVX1
X_1292_ _1253_/A _1292_/B _1291_/Y gnd _1292_/Y vdd NAND3X1
X_824_ DATA_A[16] gnd _824_/Y vdd INVX1
X_1173_ _1253_/A _1163_/Y _1173_/C gnd _1173_/Y vdd NAND3X1
X_705_ sel_A[1] _705_/B _703_/Y gnd _705_/Y vdd NAND3X1
X_1054_ _1058_/A _1054_/B gnd _1056_/C vdd NAND2X1
X_925_ _856_/A _925_/B _925_/C gnd _930_/B vdd NAND3X1
XFILL_1_0_1 gnd vdd FILL
X_1274_ _1276_/A DATA_A[3] gnd _1277_/B vdd OR2X2
X_1155_ DATA_A[0] _1160_/A gnd _1158_/B vdd OR2X2
X_806_ _801_/A _805_/Y gnd _807_/C vdd NAND2X1
XBUFX2_insert18 sel_A[8] gnd _1074_/A vdd BUFX2
X_687_ _770_/A DATA_B[4] gnd _690_/B vdd OR2X2
X_1036_ _1074_/A DATA_A[9] gnd _1037_/B vdd OR2X2
XFILL_8_0_1 gnd vdd FILL
X_907_ DATA_A[26] gnd _907_/Y vdd INVX1
X_1256_ _1187_/A _1256_/B gnd _1257_/C vdd NAND2X1
X_788_ _669_/A _785_/Y _787_/Y gnd _788_/Y vdd NAND3X1
X_1137_ DATA_B[23] gnd _1138_/B vdd INVX1
X_669_ _669_/A _669_/B _668_/Y gnd _674_/B vdd NAND3X1
X_1018_ _1018_/A _1018_/B _1017_/Y gnd _1028_/B vdd NAND3X1
X_889_ _972_/A DATA_B[9] gnd _889_/Y vdd OR2X2
X_1238_ _1158_/A _1238_/B _1238_/C gnd _1243_/B vdd NAND3X1
X_1119_ _1123_/B _1118_/Y gnd _1120_/C vdd NAND2X1
X_770_ _770_/A DATA_B[26] gnd _771_/C vdd NAND2X1
X_990_ DATA_A[16] gnd _991_/B vdd INVX1
X_651_ _651_/A gnd NIBBLE_OUT[14] vdd BUFX2
X_1000_ _991_/A _999_/Y gnd _1001_/C vdd NAND2X1
X_871_ sel_A[4] _870_/Y _869_/Y gnd _872_/C vdd NAND3X1
X_1220_ _1304_/A _1219_/Y gnd _1222_/C vdd NAND2X1
X_752_ _750_/Y _751_/A _752_/C gnd _752_/Y vdd OAI21X1
X_1101_ DATA_B[10] gnd _1103_/A vdd INVX1
XFILL_2_1_0 gnd vdd FILL
XBUFX2_insert19 sel_A[8] gnd _1030_/A vdd BUFX2
X_972_ _972_/A _971_/Y gnd _973_/C vdd NAND2X1
X_853_ _853_/A DATA_B[4] gnd _853_/Y vdd OR2X2
X_1202_ _1169_/A DATA_A[9] gnd _1203_/B vdd OR2X2
X_1083_ _1075_/A DATA_A[30] gnd _1084_/C vdd NAND2X1
X_734_ sel_B[0] _729_/Y _734_/C gnd _735_/C vdd NAND3X1
XFILL_12_1 gnd vdd FILL
X_954_ _835_/A _951_/Y _953_/Y gnd _954_/Y vdd NAND3X1
XFILL_9_1_0 gnd vdd FILL
X_1303_ DATA_B[23] gnd _1303_/Y vdd INVX1
X_835_ _835_/A _832_/Y _834_/Y gnd _835_/Y vdd NAND3X1
X_1184_ _1271_/A _1179_/Y _1184_/C gnd _1194_/B vdd NAND3X1
X_716_ _755_/A _706_/Y _716_/C gnd _716_/Y vdd NAND3X1
X_1065_ sel_B[7] _1065_/B gnd _1066_/C vdd NAND2X1
X_1285_ _1276_/A _1284_/Y gnd _1285_/Y vdd NAND2X1
X_936_ _853_/A DATA_B[26] gnd _937_/C vdd NAND2X1
X_817_ _639_/A CLK _817_/D gnd vdd DFFPOSX1
X_1166_ _1169_/A _1165_/Y gnd _1167_/C vdd NAND2X1
X_698_ _704_/A DATA_A[1] gnd _698_/Y vdd OR2X2
X_1047_ sel_A[6] _1047_/B _1047_/C gnd _1047_/Y vdd NAND3X1
X_918_ _916_/Y _823_/B _918_/C gnd _918_/Y vdd OAI21X1
XBUFX2_insert20 sel_B[2] gnd _758_/A vdd BUFX2
X_1267_ DATA_B[10] gnd _1269_/A vdd INVX1
XFILL_2_1_1 gnd vdd FILL
X_1148_ _646_/A CLK _1068_/Y gnd vdd DFFPOSX1
X_799_ DATA_B[27] gnd _799_/Y vdd INVX1
X_680_ _723_/A _679_/Y gnd _681_/C vdd NAND2X1
X_1029_ _1007_/Y _1029_/B _985_/Y gnd _1147_/D vdd AOI21X1
XFILL_12_2 gnd vdd FILL
X_1249_ _1235_/A DATA_A[30] gnd _1250_/C vdd NAND2X1
X_900_ sel_B[3] _895_/Y _900_/C gnd _901_/C vdd NAND3X1
XFILL_9_1_1 gnd vdd FILL
X_781_ _781_/A _780_/Y gnd _781_/Y vdd NAND2X1
X_1130_ _1091_/A _1130_/B _1130_/C gnd _1135_/B vdd NAND3X1
X_662_ _662_/A _661_/Y gnd _662_/Y vdd NAND2X1
X_1011_ DATA_B[16] gnd _1012_/B vdd INVX1
X_882_ _841_/A _882_/B _882_/C gnd _882_/Y vdd NAND3X1
X_1231_ sel_B[10] _1231_/B gnd _1232_/C vdd NAND2X1
X_1112_ DATA_A[27] gnd _1113_/B vdd INVX1
X_763_ sel_B[1] _762_/Y _763_/C gnd _764_/C vdd NAND3X1
X_644_ _644_/A gnd NIBBLE_OUT[7] vdd BUFX2
X_983_ _983_/Q CLK _941_/Y gnd vdd DFFPOSX1
X_864_ _823_/B DATA_A[1] gnd _864_/Y vdd OR2X2
X_1213_ sel_A[9] _1213_/B _1213_/C gnd _1214_/C vdd NAND3X1
X_745_ _665_/A _740_/Y _744_/Y gnd _745_/Y vdd NAND3X1
XBUFX2_insert21 sel_B[2] gnd _801_/A vdd BUFX2
X_1094_ _1094_/A DATA_B[14] gnd _1095_/B vdd OR2X2
X_965_ DATA_B[27] gnd _965_/Y vdd INVX1
X_1314_ _650_/A CLK _1314_/D gnd vdd DFFPOSX1
X_1195_ _1173_/Y _1195_/B _1195_/C gnd _1195_/Y vdd AOI21X1
X_846_ _922_/A _845_/Y gnd _847_/C vdd NAND2X1
X_727_ DATA_B[21] gnd _728_/B vdd INVX1
X_1076_ sel_A[7] _1076_/B _1076_/C gnd _1077_/C vdd NAND3X1
X_947_ _905_/A _946_/Y gnd _949_/C vdd NAND2X1
X_1296_ _1188_/A _1296_/B _1296_/C gnd _1301_/B vdd NAND3X1
X_828_ _828_/A _827_/Y gnd _828_/Y vdd NAND2X1
X_1177_ DATA_B[16] gnd _1177_/Y vdd INVX1
X_709_ _781_/A _708_/Y gnd _710_/C vdd NAND2X1
X_1058_ _1058_/A DATA_B[5] gnd _1058_/Y vdd OR2X2
X_929_ sel_B[4] _928_/Y _927_/Y gnd _930_/C vdd NAND3X1
X_1278_ DATA_A[27] gnd _1278_/Y vdd INVX1
X_1159_ DATA_A[24] gnd _1159_/Y vdd INVX1
XFILL_3_1 gnd vdd FILL
X_810_ _808_/Y _795_/A _810_/C gnd _810_/Y vdd OAI21X1
XBUFX2_insert22 sel_B[2] gnd _770_/A vdd BUFX2
X_691_ DATA_B[12] gnd _693_/A vdd INVX1
X_1040_ DATA_A[21] gnd _1041_/B vdd INVX1
X_911_ _831_/A _906_/Y _910_/Y gnd _911_/Y vdd NAND3X1
X_1260_ _1191_/B DATA_B[14] gnd _1261_/B vdd OR2X2
X_792_ sel_A[1] _791_/Y gnd _793_/C vdd NAND2X1
XFILL_5_0_0 gnd vdd FILL
X_1141_ _1133_/A DATA_B[31] gnd _1142_/C vdd NAND2X1
X_673_ sel_A[1] _672_/Y gnd _674_/C vdd NAND2X1
X_1022_ _1091_/A _1022_/B _1022_/C gnd _1027_/B vdd NAND3X1
X_893_ DATA_B[21] gnd _893_/Y vdd INVX1
X_1242_ sel_A[10] _1242_/B _1242_/C gnd _1243_/C vdd NAND3X1
X_1123_ _1121_/Y _1123_/B _1123_/C gnd _1123_/Y vdd OAI21X1
X_774_ SEL[0] _774_/B _774_/C gnd _775_/B vdd NAND3X1
X_994_ _991_/A _993_/Y gnd _996_/C vdd NAND2X1
X_655_ sel_A[0] gnd _665_/A vdd INVX2
X_1004_ _1004_/A _1074_/A _1004_/C gnd _1005_/B vdd OAI21X1
X_875_ _905_/A _875_/B gnd _876_/C vdd NAND2X1
X_1224_ _1302_/A DATA_B[5] gnd _1227_/B vdd OR2X2
X_756_ _758_/A DATA_B[6] gnd _759_/B vdd OR2X2
XFILL_3_2 gnd vdd FILL
X_1105_ _1018_/A _1100_/Y _1105_/C gnd _1106_/C vdd NAND3X1
X_637_ _815_/Q gnd NIBBLE_OUT[0] vdd BUFX2
X_976_ _974_/Y _963_/A _975_/Y gnd _976_/Y vdd OAI21X1
XBUFX2_insert23 sel_B[2] gnd _723_/A vdd BUFX2
X_857_ DATA_B[12] gnd _859_/A vdd INVX1
X_1206_ DATA_A[21] gnd _1207_/B vdd INVX1
X_738_ DATA_A[18] gnd _738_/Y vdd INVX1
X_1087_ _986_/Y _1087_/B _1087_/C gnd _1087_/Y vdd NAND3X1
XFILL_5_0_1 gnd vdd FILL
X_958_ sel_A[4] _957_/Y gnd _959_/C vdd NAND2X1
X_1307_ _1304_/A DATA_B[31] gnd _1308_/C vdd NAND2X1
X_839_ sel_A[4] _838_/Y gnd _839_/Y vdd NAND2X1
X_1188_ _1188_/A _1188_/B _1187_/Y gnd _1193_/B vdd NAND3X1
X_720_ _759_/A _717_/Y _720_/C gnd _725_/B vdd NAND3X1
X_1069_ _1074_/A DATA_A[2] gnd _1072_/B vdd OR2X2
X_1289_ _1287_/Y _1250_/B _1289_/C gnd _1289_/Y vdd OAI21X1
X_940_ SEL[1] _940_/B _940_/C gnd _941_/B vdd NAND3X1
X_821_ sel_A[3] gnd _831_/A vdd INVX2
X_1170_ _1170_/A _1169_/A _1169_/Y gnd _1170_/Y vdd OAI21X1
X_702_ DATA_A[25] gnd _703_/B vdd INVX1
X_1051_ _1058_/A _1051_/B gnd _1052_/C vdd NAND2X1
XFILL_3_3 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
X_922_ _922_/A DATA_B[6] gnd _925_/B vdd OR2X2
X_1271_ _1271_/A _1271_/B _1271_/C gnd _1272_/C vdd NAND3X1
XBUFX2_insert24 sel_B[2] gnd _795_/A vdd BUFX2
X_803_ _773_/A _803_/B _802_/Y gnd _803_/Y vdd NAND3X1
X_1152_ SEL[3] gnd _1253_/A vdd INVX2
X_684_ _801_/A DATA_B[8] gnd _684_/Y vdd OR2X2
X_1033_ _992_/A _1033_/B _1033_/C gnd _1038_/B vdd NAND3X1
X_904_ DATA_A[18] gnd _904_/Y vdd INVX1
X_1253_ _1253_/A _1253_/B _1253_/C gnd _1253_/Y vdd NAND3X1
X_785_ _737_/A DATA_A[7] gnd _785_/Y vdd OR2X2
XFILL_6_1_0 gnd vdd FILL
X_1134_ sel_B[7] _1134_/B _1134_/C gnd _1134_/Y vdd NAND3X1
X_666_ _662_/A DATA_A[4] gnd _669_/B vdd OR2X2
X_1015_ _1016_/A _1014_/Y gnd _1017_/C vdd NAND2X1
X_886_ _856_/A _886_/B _885_/Y gnd _886_/Y vdd NAND3X1
X_1235_ _1235_/A DATA_A[2] gnd _1238_/B vdd OR2X2
X_1116_ _997_/A _1116_/B _1116_/C gnd _1116_/Y vdd NAND3X1
X_767_ _723_/A _767_/B gnd _768_/C vdd NAND2X1
X_987_ sel_A[6] gnd _997_/A vdd INVX2
X_648_ _648_/A gnd NIBBLE_OUT[11] vdd BUFX2
X_868_ DATA_A[25] gnd _868_/Y vdd INVX1
XFILL_12_0_1 gnd vdd FILL
X_1217_ _1302_/A _1217_/B gnd _1218_/C vdd NAND2X1
X_749_ _669_/A _746_/Y _748_/Y gnd _754_/B vdd NAND3X1
XBUFX2_insert25 sel_A[5] gnd _823_/B vdd BUFX2
X_1098_ DATA_B[18] gnd _1099_/B vdd INVX1
X_969_ _939_/A _964_/Y _969_/C gnd _969_/Y vdd NAND3X1
X_850_ _849_/A DATA_B[8] gnd _850_/Y vdd OR2X2
X_1199_ _1158_/A _1199_/B _1198_/Y gnd _1199_/Y vdd NAND3X1
XFILL_7_1 gnd vdd FILL
X_1080_ _1123_/B _1079_/Y gnd _1081_/C vdd NAND2X1
X_731_ _723_/A DATA_B[29] gnd _732_/C vdd NAND2X1
X_951_ _957_/B DATA_A[7] gnd _951_/Y vdd OR2X2
XFILL_6_1_1 gnd vdd FILL
X_1300_ sel_B[10] _1300_/B _1300_/C gnd _1301_/C vdd NAND3X1
X_832_ _944_/A DATA_A[4] gnd _832_/Y vdd OR2X2
X_1181_ _1293_/A _1181_/B gnd _1183_/C vdd NAND2X1
X_713_ _711_/Y _704_/A _713_/C gnd _713_/Y vdd OAI21X1
X_1062_ DATA_B[13] gnd _1064_/A vdd INVX1
X_933_ _849_/A _932_/Y gnd _934_/C vdd NAND2X1
X_1282_ _1282_/A _1277_/Y _1281_/Y gnd _1292_/B vdd NAND3X1
X_814_ _814_/A _814_/B _653_/Y gnd _814_/Y vdd AOI21X1
X_1163_ _1282_/A _1163_/B _1163_/C gnd _1163_/Y vdd NAND3X1
X_1044_ _1075_/A DATA_A[29] gnd _1045_/C vdd NAND2X1
X_695_ sel_B[0] _695_/B _695_/C gnd _696_/C vdd NAND3X1
XBUFX2_insert26 sel_A[5] gnd _905_/A vdd BUFX2
XFILL_13_1_0 gnd vdd FILL
X_915_ _835_/A _912_/Y _914_/Y gnd _920_/B vdd NAND3X1
X_1264_ DATA_B[18] gnd _1265_/B vdd INVX1
X_796_ DATA_B[19] gnd _797_/B vdd INVX1
X_1145_ SEL[2] _1145_/B _1145_/C gnd _1146_/B vdd NAND3X1
X_677_ sel_B[1] gnd _759_/A vdd INVX4
X_1026_ sel_B[7] _1026_/B gnd _1027_/C vdd NAND2X1
X_897_ _972_/A DATA_B[29] gnd _897_/Y vdd NAND2X1
X_1246_ _1250_/B _1245_/Y gnd _1247_/C vdd NAND2X1
X_778_ _781_/A _778_/B gnd _778_/Y vdd NAND2X1
X_1127_ _1133_/A DATA_B[3] gnd _1130_/B vdd OR2X2
X_998_ _991_/A DATA_A[4] gnd _998_/Y vdd OR2X2
X_659_ _704_/A _658_/Y gnd _660_/C vdd NAND2X1
X_1008_ sel_B[6] gnd _1018_/A vdd INVX2
X_879_ _879_/A _944_/A _878_/Y gnd _879_/Y vdd OAI21X1
X_1228_ DATA_B[13] gnd _1230_/A vdd INVX1
X_760_ DATA_B[30] gnd _761_/B vdd INVX1
X_1109_ DATA_A[19] gnd _1110_/B vdd INVX1
X_980_ _960_/Y _980_/B _980_/C gnd _984_/D vdd AOI21X1
X_641_ _981_/Q gnd NIBBLE_OUT[4] vdd BUFX2
XBUFX2_insert27 sel_A[5] gnd _957_/B vdd BUFX2
XFILL_13_1_1 gnd vdd FILL
X_861_ sel_B[3] _861_/B _861_/C gnd _862_/C vdd NAND3X1
X_1210_ _1169_/A DATA_A[29] gnd _1210_/Y vdd NAND2X1
X_742_ _751_/A _742_/B gnd _744_/C vdd NAND2X1
X_1091_ _1091_/A _1091_/B _1091_/C gnd _1096_/B vdd NAND3X1
X_962_ DATA_B[19] gnd _962_/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
X_1311_ SEL[3] _1311_/B _1311_/C gnd _1312_/B vdd NAND3X1
X_843_ sel_B[4] gnd _856_/A vdd INVX4
X_1192_ sel_B[10] _1192_/B gnd _1193_/C vdd NAND2X1
X_724_ sel_B[1] _724_/B _724_/C gnd _725_/C vdd NAND3X1
XFILL_11_1 gnd vdd FILL
X_1073_ DATA_A[26] gnd _1074_/B vdd INVX1
XFILL_9_0_0 gnd vdd FILL
X_944_ _944_/A _943_/Y gnd _945_/C vdd NAND2X1
X_1293_ _1293_/A DATA_B[3] gnd _1296_/B vdd OR2X2
X_825_ _823_/B _824_/Y gnd _826_/C vdd NAND2X1
X_1174_ sel_B[9] gnd _1271_/A vdd INVX2
X_706_ _665_/A _706_/B _705_/Y gnd _706_/Y vdd NAND3X1
X_1055_ _1058_/A DATA_B[9] gnd _1056_/B vdd OR2X2
X_926_ DATA_B[30] gnd _927_/B vdd INVX1
X_1275_ DATA_A[19] gnd _1275_/Y vdd INVX1
X_1156_ DATA_A[16] gnd _1156_/Y vdd INVX1
X_807_ _759_/A _804_/Y _807_/C gnd _807_/Y vdd NAND3X1
XBUFX2_insert28 sel_A[5] gnd _944_/A vdd BUFX2
X_688_ DATA_B[20] gnd _689_/B vdd INVX1
X_1037_ sel_A[7] _1037_/B _1037_/C gnd _1037_/Y vdd NAND3X1
X_908_ _905_/A _907_/Y gnd _910_/C vdd NAND2X1
X_1257_ _1188_/A _1257_/B _1257_/C gnd _1262_/B vdd NAND3X1
XFILL_2_0_1 gnd vdd FILL
X_789_ DATA_A[15] gnd _789_/Y vdd INVX1
X_1138_ _1016_/A _1138_/B gnd _1139_/C vdd NAND2X1
X_670_ DATA_A[12] gnd _670_/Y vdd INVX1
X_1019_ _1019_/A DATA_B[4] gnd _1022_/B vdd OR2X2
X_890_ sel_B[4] _889_/Y _890_/C gnd _891_/C vdd NAND3X1
XFILL_9_0_1 gnd vdd FILL
X_1239_ DATA_A[26] gnd _1240_/B vdd INVX1
X_1120_ _992_/A _1120_/B _1120_/C gnd _1120_/Y vdd NAND3X1
X_771_ _771_/A _770_/A _771_/C gnd _772_/B vdd OAI21X1
X_991_ _991_/A _991_/B gnd _992_/C vdd NAND2X1
X_652_ _652_/A gnd NIBBLE_OUT[15] vdd BUFX2
X_1001_ _992_/A _998_/Y _1001_/C gnd _1006_/B vdd NAND3X1
X_872_ _831_/A _867_/Y _872_/C gnd _882_/B vdd NAND3X1
X_1221_ _1304_/A DATA_B[9] gnd _1222_/B vdd OR2X2
X_753_ sel_A[1] _752_/Y gnd _754_/C vdd NAND2X1
X_1102_ _1094_/A DATA_B[26] gnd _1103_/C vdd NAND2X1
XBUFX2_insert29 sel_A[5] gnd _828_/A vdd BUFX2
X_973_ _856_/A _970_/Y _973_/C gnd _973_/Y vdd NAND3X1
X_854_ DATA_B[20] gnd _855_/B vdd INVX1
X_1203_ sel_A[10] _1203_/B _1201_/Y gnd _1204_/C vdd NAND3X1
X_1084_ _1084_/A _1075_/A _1084_/C gnd _1085_/B vdd OAI21X1
X_735_ SEL[0] _735_/B _735_/C gnd _736_/B vdd NAND3X1
X_955_ DATA_A[15] gnd _955_/Y vdd INVX1
XFILL_3_1_0 gnd vdd FILL
X_1304_ _1304_/A _1303_/Y gnd _1305_/C vdd NAND2X1
X_836_ DATA_A[12] gnd _836_/Y vdd INVX1
X_1185_ _1187_/A DATA_B[4] gnd _1188_/B vdd OR2X2
X_717_ _758_/A DATA_B[1] gnd _717_/Y vdd OR2X2
X_1066_ sel_B[6] _1066_/B _1066_/C gnd _1066_/Y vdd NAND3X1
X_1286_ _1158_/A _1283_/Y _1285_/Y gnd _1286_/Y vdd NAND3X1
X_937_ _935_/Y _853_/A _937_/C gnd _938_/B vdd OAI21X1
X_818_ _818_/Q CLK _814_/Y gnd vdd DFFPOSX1
X_1167_ _1158_/A _1164_/Y _1167_/C gnd _1167_/Y vdd NAND3X1
X_699_ DATA_A[17] gnd _700_/B vdd INVX1
X_1048_ _986_/Y _1048_/B _1047_/Y gnd _1048_/Y vdd NAND3X1
X_919_ sel_A[4] _918_/Y gnd _920_/C vdd NAND2X1
XBUFX2_insert30 sel_A[2] gnd _662_/A vdd BUFX2
X_1268_ _1191_/B DATA_B[26] gnd _1268_/Y vdd NAND2X1
XFILL_2_1 gnd vdd FILL
X_800_ _801_/A _799_/Y gnd _800_/Y vdd NAND2X1
X_1149_ _647_/A CLK _1107_/Y gnd vdd DFFPOSX1
X_681_ _759_/A _681_/B _681_/C gnd _686_/B vdd NAND3X1
X_1030_ _1030_/A DATA_A[1] gnd _1033_/B vdd OR2X2
X_1250_ _1248_/Y _1250_/B _1250_/C gnd _1250_/Y vdd OAI21X1
X_901_ SEL[1] _901_/B _901_/C gnd _902_/B vdd NAND3X1
XFILL_3_1_1 gnd vdd FILL
X_782_ _781_/A DATA_A[11] gnd _783_/B vdd OR2X2
X_1131_ DATA_B[27] gnd _1132_/B vdd INVX1
X_663_ _662_/A DATA_A[8] gnd _664_/B vdd OR2X2
X_1012_ _1019_/A _1012_/B gnd _1013_/C vdd NAND2X1
X_883_ _963_/A DATA_B[1] gnd _886_/B vdd OR2X2
X_1232_ sel_B[9] _1232_/B _1232_/C gnd _1233_/C vdd NAND3X1
X_1113_ _1123_/B _1113_/B gnd _1115_/C vdd NAND2X1
X_764_ sel_B[0] _764_/B _764_/C gnd _774_/B vdd NAND3X1
X_984_ _644_/A CLK _984_/D gnd vdd DFFPOSX1
X_645_ _645_/A gnd NIBBLE_OUT[8] vdd BUFX2
X_865_ DATA_A[17] gnd _865_/Y vdd INVX1
X_1214_ _1253_/A _1214_/B _1214_/C gnd _1214_/Y vdd NAND3X1
XBUFX2_insert31 sel_A[2] gnd _751_/A vdd BUFX2
X_746_ _737_/A DATA_A[6] gnd _746_/Y vdd OR2X2
XFILL_2_2 gnd vdd FILL
XFILL_10_1_0 gnd vdd FILL
X_1095_ sel_B[7] _1095_/B _1095_/C gnd _1096_/C vdd NAND3X1
X_966_ _972_/A _965_/Y gnd _968_/C vdd NAND2X1
X_1315_ _651_/A CLK _1273_/Y gnd vdd DFFPOSX1
X_1196_ _1235_/A DATA_A[1] gnd _1199_/B vdd OR2X2
X_847_ _856_/A _847_/B _847_/C gnd _852_/B vdd NAND3X1
X_728_ _795_/A _728_/B gnd _728_/Y vdd NAND2X1
X_1077_ _997_/A _1077_/B _1077_/C gnd _1087_/B vdd NAND3X1
X_948_ _905_/A DATA_A[11] gnd _948_/Y vdd OR2X2
X_1297_ DATA_B[27] gnd _1297_/Y vdd INVX1
X_829_ _828_/A DATA_A[8] gnd _830_/B vdd OR2X2
X_1178_ _1293_/A _1177_/Y gnd _1179_/C vdd NAND2X1
X_710_ _669_/A _710_/B _710_/C gnd _715_/B vdd NAND3X1
X_1059_ DATA_B[21] gnd _1059_/Y vdd INVX1
X_930_ sel_B[3] _930_/B _930_/C gnd _940_/B vdd NAND3X1
X_1279_ _1276_/A _1278_/Y gnd _1281_/C vdd NAND2X1
X_1160_ _1160_/A _1159_/Y gnd _1162_/C vdd NAND2X1
X_811_ sel_B[1] _810_/Y gnd _811_/Y vdd NAND2X1
XBUFX2_insert32 sel_A[2] gnd _704_/A vdd BUFX2
X_692_ _770_/A DATA_B[28] gnd _693_/C vdd NAND2X1
XFILL_2_3 gnd vdd FILL
X_1041_ _1030_/A _1041_/B gnd _1042_/C vdd NAND2X1
XFILL_10_1_1 gnd vdd FILL
X_912_ _957_/B DATA_A[6] gnd _912_/Y vdd OR2X2
X_1261_ sel_B[10] _1261_/B _1261_/C gnd _1262_/C vdd NAND3X1
X_793_ sel_A[0] _788_/Y _793_/C gnd _793_/Y vdd NAND3X1
X_1142_ _1142_/A _1133_/A _1142_/C gnd _1143_/B vdd OAI21X1
X_674_ sel_A[0] _674_/B _674_/C gnd _674_/Y vdd NAND3X1
X_1023_ DATA_B[12] gnd _1025_/A vdd INVX1
X_894_ _963_/A _893_/Y gnd _894_/Y vdd NAND2X1
X_1243_ _1282_/A _1243_/B _1243_/C gnd _1253_/B vdd NAND3X1
X_1124_ sel_A[7] _1123_/Y gnd _1124_/Y vdd NAND2X1
XFILL_6_0_0 gnd vdd FILL
X_775_ _775_/A _775_/B _653_/Y gnd _817_/D vdd AOI21X1
X_656_ sel_A[1] gnd _669_/A vdd INVX4
X_995_ _991_/A DATA_A[8] gnd _996_/B vdd OR2X2
X_1005_ sel_A[7] _1005_/B gnd _1005_/Y vdd NAND2X1
X_876_ _835_/A _876_/B _876_/C gnd _881_/B vdd NAND3X1
X_1225_ DATA_B[21] gnd _1226_/B vdd INVX1
X_757_ DATA_B[22] gnd _758_/B vdd INVX1
X_1106_ SEL[2] _1106_/B _1106_/C gnd _1107_/B vdd NAND3X1
X_977_ sel_B[4] _976_/Y gnd _978_/C vdd NAND2X1
X_638_ _638_/A gnd NIBBLE_OUT[1] vdd BUFX2
XBUFX2_insert33 sel_A[2] gnd _781_/A vdd BUFX2
X_858_ _853_/A DATA_B[28] gnd _859_/C vdd NAND2X1
X_1207_ _1250_/B _1207_/B gnd _1208_/C vdd NAND2X1
X_739_ _751_/A _738_/Y gnd _739_/Y vdd NAND2X1
X_1088_ _1019_/A DATA_B[6] gnd _1091_/B vdd OR2X2
X_959_ sel_A[3] _954_/Y _959_/C gnd _960_/C vdd NAND3X1
X_1308_ _1308_/A _1304_/A _1308_/C gnd _1309_/B vdd OAI21X1
X_840_ sel_A[3] _835_/Y _839_/Y gnd _841_/C vdd NAND3X1
XFILL_6_1 gnd vdd FILL
X_1189_ DATA_B[12] gnd _1191_/A vdd INVX1
X_721_ DATA_B[25] gnd _722_/B vdd INVX1
X_1070_ DATA_A[18] gnd _1071_/B vdd INVX1
XFILL_6_0_1 gnd vdd FILL
X_1290_ sel_A[10] _1289_/Y gnd _1291_/C vdd NAND2X1
X_941_ _941_/A _941_/B _980_/C gnd _941_/Y vdd AOI21X1
X_822_ sel_A[4] gnd _835_/A vdd INVX4
X_1171_ sel_A[10] _1170_/Y gnd _1172_/C vdd NAND2X1
X_703_ _662_/A _703_/B gnd _703_/Y vdd NAND2X1
X_1052_ _1091_/A _1052_/B _1052_/C gnd _1057_/B vdd NAND3X1
X_923_ DATA_B[22] gnd _923_/Y vdd INVX1
X_1272_ SEL[3] _1272_/B _1272_/C gnd _1273_/B vdd NAND3X1
X_1153_ sel_A[9] gnd _1282_/A vdd INVX2
XBUFX2_insert34 sel_A[2] gnd _737_/A vdd BUFX2
X_804_ _795_/A DATA_B[7] gnd _804_/Y vdd OR2X2
X_685_ sel_B[1] _684_/Y _683_/Y gnd _685_/Y vdd NAND3X1
X_1034_ DATA_A[25] gnd _1035_/B vdd INVX1
X_905_ _905_/A _904_/Y gnd _906_/C vdd NAND2X1
XFILL_13_0_0 gnd vdd FILL
X_1254_ _1187_/A DATA_B[6] gnd _1257_/B vdd OR2X2
X_786_ DATA_A[23] gnd _786_/Y vdd INVX1
XFILL_6_2 gnd vdd FILL
X_1135_ _1018_/A _1135_/B _1134_/Y gnd _1145_/B vdd NAND3X1
XFILL_0_1_0 gnd vdd FILL
X_667_ DATA_A[20] gnd _668_/B vdd INVX1
X_1016_ _1016_/A DATA_B[8] gnd _1017_/B vdd OR2X2
X_887_ DATA_B[25] gnd _887_/Y vdd INVX1
X_1236_ DATA_A[18] gnd _1236_/Y vdd INVX1
X_1117_ _1123_/B DATA_A[7] gnd _1120_/B vdd OR2X2
XFILL_7_1_0 gnd vdd FILL
X_768_ _759_/A _768_/B _768_/C gnd _768_/Y vdd NAND3X1
X_988_ sel_A[7] gnd _992_/A vdd INVX4
X_649_ _649_/A gnd NIBBLE_OUT[12] vdd BUFX2
X_869_ _828_/A _868_/Y gnd _869_/Y vdd NAND2X1
X_1218_ _1188_/A _1218_/B _1218_/C gnd _1223_/B vdd NAND3X1
X_750_ DATA_A[14] gnd _750_/Y vdd INVX1
XBUFX2_insert35 sel_B[11] gnd _1304_/A vdd BUFX2
X_1099_ _1016_/A _1099_/B gnd _1100_/C vdd NAND2X1
X_970_ _963_/A DATA_B[7] gnd _970_/Y vdd OR2X2
X_851_ sel_B[4] _850_/Y _849_/Y gnd _851_/Y vdd NAND3X1
X_1200_ DATA_A[25] gnd _1200_/Y vdd INVX1
XFILL_13_0_1 gnd vdd FILL
X_1081_ _992_/A _1081_/B _1081_/C gnd _1086_/B vdd NAND3X1
X_732_ _732_/A _801_/A _732_/C gnd _733_/B vdd OAI21X1
X_952_ DATA_A[23] gnd _952_/Y vdd INVX1
XFILL_0_1_1 gnd vdd FILL
X_1301_ _1271_/A _1301_/B _1301_/C gnd _1311_/B vdd NAND3X1
X_833_ DATA_A[20] gnd _833_/Y vdd INVX1
X_1182_ _1293_/A DATA_B[8] gnd _1182_/Y vdd OR2X2
X_714_ sel_A[1] _713_/Y gnd _715_/C vdd NAND2X1
XFILL_7_1_1 gnd vdd FILL
X_1063_ _1133_/A DATA_B[29] gnd _1064_/C vdd NAND2X1
XFILL_10_1 gnd vdd FILL
X_1283_ _1276_/A DATA_A[7] gnd _1283_/Y vdd OR2X2
X_934_ _856_/A _931_/Y _934_/C gnd _934_/Y vdd NAND3X1
X_815_ _815_/Q CLK _815_/D gnd vdd DFFPOSX1
X_1164_ _1235_/A DATA_A[4] gnd _1164_/Y vdd OR2X2
X_1045_ _1045_/A _1075_/A _1045_/C gnd _1046_/B vdd OAI21X1
X_696_ SEL[0] _696_/B _696_/C gnd _697_/B vdd NAND3X1
X_916_ DATA_A[14] gnd _916_/Y vdd INVX1
XBUFX2_insert36 sel_B[11] gnd _1293_/A vdd BUFX2
X_1265_ _1293_/A _1265_/B gnd _1266_/C vdd NAND2X1
X_1146_ _1146_/A _1146_/B _985_/Y gnd _1150_/D vdd AOI21X1
X_797_ _795_/A _797_/B gnd _798_/C vdd NAND2X1
X_678_ DATA_B[0] _723_/A gnd _681_/B vdd OR2X2
X_1027_ sel_B[6] _1027_/B _1027_/C gnd _1028_/C vdd NAND3X1
XBUFX2_insert0 sel_A[11] gnd _1250_/B vdd BUFX2
X_898_ _896_/Y _972_/A _897_/Y gnd _898_/Y vdd OAI21X1
X_779_ _669_/A _779_/B _778_/Y gnd _784_/B vdd NAND3X1
X_1247_ _1158_/A _1244_/Y _1247_/C gnd _1252_/B vdd NAND3X1
X_1128_ DATA_B[19] gnd _1128_/Y vdd INVX1
X_999_ DATA_A[20] gnd _999_/Y vdd INVX1
X_660_ _669_/A _657_/Y _660_/C gnd _660_/Y vdd NAND3X1
X_1009_ sel_B[7] gnd _1091_/A vdd INVX4
XFILL_10_2 gnd vdd FILL
X_880_ sel_A[4] _879_/Y gnd _881_/C vdd NAND2X1
X_1229_ _1304_/A DATA_B[29] gnd _1230_/C vdd NAND2X1
X_761_ _758_/A _761_/B gnd _763_/C vdd NAND2X1
X_1110_ _1030_/A _1110_/B gnd _1111_/C vdd NAND2X1
X_981_ _981_/Q CLK _863_/Y gnd vdd DFFPOSX1
X_642_ _982_/Q gnd NIBBLE_OUT[5] vdd BUFX2
XBUFX2_insert37 sel_B[11] gnd _1302_/A vdd BUFX2
X_862_ SEL[1] _862_/B _862_/C gnd _863_/B vdd NAND3X1
X_1211_ _1211_/A _1169_/A _1210_/Y gnd _1212_/B vdd OAI21X1
X_743_ _751_/A DATA_A[10] gnd _743_/Y vdd OR2X2
X_1092_ DATA_B[30] gnd _1093_/B vdd INVX1
X_963_ _963_/A _962_/Y gnd _964_/C vdd NAND2X1
X_1312_ _1292_/Y _1312_/B _1195_/C gnd _1316_/D vdd AOI21X1
XBUFX2_insert1 sel_A[11] gnd _1169_/A vdd BUFX2
X_844_ DATA_B[0] _922_/A gnd _847_/B vdd OR2X2
X_1193_ sel_B[9] _1193_/B _1193_/C gnd _1194_/C vdd NAND3X1
X_725_ _773_/A _725_/B _725_/C gnd _735_/B vdd NAND3X1
X_1074_ _1074_/A _1074_/B gnd _1076_/C vdd NAND2X1
X_945_ _835_/A _945_/B _945_/C gnd _950_/B vdd NAND3X1
XFILL_3_0_0 gnd vdd FILL
X_1294_ DATA_B[19] gnd _1295_/B vdd INVX1
X_826_ _835_/A _823_/Y _826_/C gnd _826_/Y vdd NAND3X1
X_1175_ sel_B[10] gnd _1188_/A vdd INVX4
X_707_ _781_/A DATA_A[5] gnd _710_/B vdd OR2X2
X_1056_ sel_B[7] _1056_/B _1056_/C gnd _1057_/C vdd NAND3X1
X_927_ _922_/A _927_/B gnd _927_/Y vdd NAND2X1
X_1276_ _1276_/A _1275_/Y gnd _1276_/Y vdd NAND2X1
X_1157_ _1160_/A _1156_/Y gnd _1157_/Y vdd NAND2X1
X_808_ DATA_B[15] gnd _808_/Y vdd INVX1
XBUFX2_insert38 sel_B[11] gnd _1191_/B vdd BUFX2
X_689_ _770_/A _689_/B gnd _690_/C vdd NAND2X1
X_1038_ _997_/A _1038_/B _1037_/Y gnd _1048_/B vdd NAND3X1
X_909_ _823_/B DATA_A[10] gnd _909_/Y vdd OR2X2
X_1258_ DATA_B[30] gnd _1259_/B vdd INVX1
XFILL_1_1 gnd vdd FILL
X_790_ _737_/A DATA_A[31] gnd _791_/C vdd NAND2X1
X_1139_ _1091_/A _1139_/B _1139_/C gnd _1144_/B vdd NAND3X1
X_671_ _662_/A DATA_A[28] gnd _672_/C vdd NAND2X1
XBUFX2_insert2 sel_A[11] gnd _1160_/A vdd BUFX2
X_1020_ DATA_B[20] gnd _1021_/B vdd INVX1
X_891_ _939_/A _886_/Y _891_/C gnd _901_/B vdd NAND3X1
X_1240_ _1160_/A _1240_/B gnd _1242_/C vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
X_1121_ DATA_A[15] gnd _1121_/Y vdd INVX1
X_772_ sel_B[1] _772_/B gnd _772_/Y vdd NAND2X1
X_992_ _992_/A _992_/B _992_/C gnd _997_/B vdd NAND3X1
X_653_ RESET_L gnd _653_/Y vdd INVX2
X_1002_ DATA_A[12] gnd _1004_/A vdd INVX1
X_873_ _905_/A DATA_A[5] gnd _876_/B vdd OR2X2
X_1222_ sel_B[10] _1222_/B _1222_/C gnd _1223_/C vdd NAND3X1
X_754_ sel_A[0] _754_/B _754_/C gnd _755_/C vdd NAND3X1
XFILL_14_1 gnd vdd FILL
X_1103_ _1103_/A _1094_/A _1103_/C gnd _1104_/B vdd OAI21X1
X_974_ DATA_B[15] gnd _974_/Y vdd INVX1
XBUFX2_insert39 sel_B[11] gnd _1187_/A vdd BUFX2
X_855_ _853_/A _855_/B gnd _855_/Y vdd NAND2X1
X_1204_ _1282_/A _1199_/Y _1204_/C gnd _1214_/B vdd NAND3X1
X_1085_ sel_A[7] _1085_/B gnd _1086_/C vdd NAND2X1
X_736_ _716_/Y _736_/B _653_/Y gnd _816_/D vdd AOI21X1
XFILL_10_0_0 gnd vdd FILL
XFILL_1_2 gnd vdd FILL
X_956_ _957_/B DATA_A[31] gnd _957_/C vdd NAND2X1
XBUFX2_insert3 sel_A[11] gnd _1276_/A vdd BUFX2
X_1305_ _1188_/A _1302_/Y _1305_/C gnd _1310_/B vdd NAND3X1
X_837_ _944_/A DATA_A[28] gnd _838_/C vdd NAND2X1
X_1186_ DATA_B[20] gnd _1187_/B vdd INVX1
X_718_ DATA_B[17] gnd _718_/Y vdd INVX1
X_1067_ SEL[2] _1067_/B _1066_/Y gnd _1068_/B vdd NAND3X1
X_1287_ DATA_A[15] gnd _1287_/Y vdd INVX1
X_938_ sel_B[4] _938_/B gnd _938_/Y vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
X_819_ RESET_L gnd _980_/C vdd INVX2
X_1168_ DATA_A[12] gnd _1170_/A vdd INVX1
X_700_ _704_/A _700_/B gnd _701_/C vdd NAND2X1
X_1049_ _1058_/A DATA_B[1] gnd _1052_/B vdd OR2X2
X_920_ sel_A[3] _920_/B _920_/C gnd _920_/Y vdd NAND3X1
XFILL_14_2 gnd vdd FILL
X_1269_ _1269_/A _1191_/B _1268_/Y gnd _1270_/B vdd OAI21X1
X_1150_ _648_/A CLK _1150_/D gnd vdd DFFPOSX1
X_801_ _801_/A DATA_B[11] gnd _801_/Y vdd OR2X2
X_682_ DATA_B[24] gnd _682_/Y vdd INVX1
X_1031_ DATA_A[17] gnd _1032_/B vdd INVX1
XFILL_1_3 gnd vdd FILL
X_1251_ sel_A[10] _1250_/Y gnd _1252_/C vdd NAND2X1
X_902_ _882_/Y _902_/B _980_/C gnd _982_/D vdd AOI21X1
XFILL_10_0_1 gnd vdd FILL
XBUFX2_insert4 sel_A[11] gnd _1235_/A vdd BUFX2
X_783_ sel_A[1] _783_/B _781_/Y gnd _783_/Y vdd NAND3X1
X_1132_ _1016_/A _1132_/B gnd _1134_/C vdd NAND2X1
X_664_ sel_A[1] _664_/B _662_/Y gnd _664_/Y vdd NAND3X1
X_1013_ _1091_/A _1013_/B _1013_/C gnd _1018_/B vdd NAND3X1
X_884_ DATA_B[17] gnd _884_/Y vdd INVX1
X_1233_ SEL[3] _1233_/B _1233_/C gnd _1234_/B vdd NAND3X1
XFILL_4_1_1 gnd vdd FILL
X_1114_ _1030_/A DATA_A[11] gnd _1115_/B vdd OR2X2
X_765_ _758_/A DATA_B[2] gnd _768_/B vdd OR2X2
X_646_ _646_/A gnd NIBBLE_OUT[9] vdd BUFX2
X_985_ RESET_L gnd _985_/Y vdd INVX2
X_866_ _828_/A _865_/Y gnd _866_/Y vdd NAND2X1
XFILL_14_3 gnd vdd FILL
X_1215_ _1293_/A DATA_B[1] gnd _1218_/B vdd OR2X2
X_747_ DATA_A[22] gnd _747_/Y vdd INVX1
X_1096_ sel_B[6] _1096_/B _1096_/C gnd _1106_/B vdd NAND3X1
X_967_ _972_/A DATA_B[11] gnd _968_/B vdd OR2X2
X_1316_ _652_/A CLK _1316_/D gnd vdd DFFPOSX1
X_848_ DATA_B[24] gnd _848_/Y vdd INVX1
X_1197_ DATA_A[17] gnd _1197_/Y vdd INVX1
X_1078_ _1123_/B DATA_A[6] gnd _1081_/B vdd OR2X2
X_729_ _759_/A _726_/Y _728_/Y gnd _729_/Y vdd NAND3X1
XBUFX2_insert5 sel_B[8] gnd _1016_/A vdd BUFX2
XFILL_11_1_0 gnd vdd FILL
X_949_ sel_A[4] _948_/Y _949_/C gnd _950_/C vdd NAND3X1
X_1298_ _1302_/A _1297_/Y gnd _1300_/C vdd NAND2X1
X_830_ sel_A[4] _830_/B _828_/Y gnd _830_/Y vdd NAND3X1
X_711_ DATA_A[13] gnd _711_/Y vdd INVX1
X_1179_ _1188_/A _1176_/Y _1179_/C gnd _1179_/Y vdd NAND3X1
X_1060_ _1058_/A _1059_/Y gnd _1061_/C vdd NAND2X1
X_931_ _849_/A DATA_B[2] gnd _931_/Y vdd OR2X2
X_1280_ _1276_/A DATA_A[11] gnd _1280_/Y vdd OR2X2
X_1161_ _1160_/A DATA_A[8] gnd _1162_/B vdd OR2X2
X_812_ sel_B[0] _807_/Y _811_/Y gnd _813_/C vdd NAND3X1
X_693_ _693_/A _770_/A _693_/C gnd _694_/B vdd OAI21X1
X_1042_ _992_/A _1042_/B _1042_/C gnd _1047_/B vdd NAND3X1
X_913_ DATA_A[22] gnd _913_/Y vdd INVX1
X_1262_ sel_B[9] _1262_/B _1262_/C gnd _1272_/B vdd NAND3X1
X_794_ _755_/A _794_/B _793_/Y gnd _814_/A vdd NAND3X1
X_1143_ sel_B[7] _1143_/B gnd _1144_/C vdd NAND2X1
X_675_ _755_/A _665_/Y _674_/Y gnd _697_/A vdd NAND3X1
XBUFX2_insert6 sel_B[8] gnd _1133_/A vdd BUFX2
X_1024_ _1094_/A DATA_B[28] gnd _1025_/C vdd NAND2X1
X_895_ _856_/A _892_/Y _894_/Y gnd _895_/Y vdd NAND3X1
XFILL_11_1_1 gnd vdd FILL
X_1244_ _1250_/B DATA_A[6] gnd _1244_/Y vdd OR2X2
X_1125_ sel_A[6] _1120_/Y _1124_/Y gnd _1126_/C vdd NAND3X1
X_776_ _781_/A DATA_A[3] gnd _779_/B vdd OR2X2
XFILL_0_0_0 gnd vdd FILL
X_996_ sel_A[7] _996_/B _996_/C gnd _997_/C vdd NAND3X1
X_657_ DATA_A[0] _751_/A gnd _657_/Y vdd OR2X2
X_1006_ sel_A[6] _1006_/B _1005_/Y gnd _1007_/C vdd NAND3X1
X_877_ DATA_A[13] gnd _879_/A vdd INVX1
X_1226_ _1302_/A _1226_/B gnd _1227_/C vdd NAND2X1
X_758_ _758_/A _758_/B gnd _758_/Y vdd NAND2X1
XFILL_7_0_0 gnd vdd FILL
X_1107_ _1087_/Y _1107_/B _985_/Y gnd _1107_/Y vdd AOI21X1
X_639_ _639_/A gnd NIBBLE_OUT[2] vdd BUFX2
X_978_ sel_B[3] _973_/Y _978_/C gnd _979_/C vdd NAND3X1
X_859_ _859_/A _853_/A _859_/C gnd _860_/B vdd OAI21X1
X_1208_ _1158_/A _1205_/Y _1208_/C gnd _1213_/B vdd NAND3X1
X_740_ _669_/A _737_/Y _739_/Y gnd _740_/Y vdd NAND3X1
X_1089_ DATA_B[22] gnd _1090_/B vdd INVX1
X_960_ _841_/A _950_/Y _960_/C gnd _960_/Y vdd NAND3X1
X_1309_ sel_B[10] _1309_/B gnd _1310_/C vdd NAND2X1
X_841_ _841_/A _831_/Y _841_/C gnd _841_/Y vdd NAND3X1
X_1190_ _1191_/B DATA_B[28] gnd _1191_/C vdd NAND2X1
XBUFX2_insert7 sel_B[8] gnd _1094_/A vdd BUFX2
X_722_ _723_/A _722_/B gnd _724_/C vdd NAND2X1
X_1071_ _1075_/A _1071_/B gnd _1072_/C vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
X_942_ _905_/A DATA_A[3] gnd _945_/B vdd OR2X2
X_1291_ sel_A[9] _1286_/Y _1291_/C gnd _1291_/Y vdd NAND3X1
X_823_ DATA_A[0] _823_/B gnd _823_/Y vdd OR2X2
X_1172_ sel_A[9] _1167_/Y _1172_/C gnd _1173_/C vdd NAND3X1
X_704_ _704_/A DATA_A[9] gnd _705_/B vdd OR2X2
X_1053_ DATA_B[25] gnd _1054_/B vdd INVX1
X_924_ _922_/A _923_/Y gnd _925_/C vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
X_1273_ _1253_/Y _1273_/B _1195_/C gnd _1273_/Y vdd AOI21X1
X_1154_ sel_A[10] gnd _1158_/A vdd INVX4
X_805_ DATA_B[23] gnd _805_/Y vdd INVX1
X_686_ _773_/A _686_/B _685_/Y gnd _696_/B vdd NAND3X1
X_1035_ _1074_/A _1035_/B gnd _1037_/C vdd NAND2X1
X_906_ _835_/A _903_/Y _906_/C gnd _906_/Y vdd NAND3X1
X_1255_ DATA_B[22] gnd _1256_/B vdd INVX1
X_787_ _737_/A _786_/Y gnd _787_/Y vdd NAND2X1
X_1136_ _1016_/A DATA_B[7] gnd _1139_/B vdd OR2X2
XBUFX2_insert8 sel_B[8] gnd _1019_/A vdd BUFX2
.ends

