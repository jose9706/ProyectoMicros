module selector4 (DATA_A, DATA_B, sel_A, sel_B, SEL, RESET_L, CLK, temp);

input RESET_L;
input CLK;
input [31:0] DATA_A;
input [31:0] DATA_B;
input [11:0] sel_A;
input [11:0] sel_B;
input [3:0] SEL;
output [15:0] temp;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(sel_A[11]), .Y(sel_A_11_bF_buf4_) );
BUFX4 BUFX4_2 ( .A(sel_A[11]), .Y(sel_A_11_bF_buf3_) );
BUFX4 BUFX4_3 ( .A(sel_A[11]), .Y(sel_A_11_bF_buf2_) );
BUFX4 BUFX4_4 ( .A(sel_A[11]), .Y(sel_A_11_bF_buf1_) );
BUFX4 BUFX4_5 ( .A(sel_A[11]), .Y(sel_A_11_bF_buf0_) );
BUFX4 BUFX4_6 ( .A(sel_B[8]), .Y(sel_B_8_bF_buf4_) );
BUFX4 BUFX4_7 ( .A(sel_B[8]), .Y(sel_B_8_bF_buf3_) );
BUFX4 BUFX4_8 ( .A(sel_B[8]), .Y(sel_B_8_bF_buf2_) );
BUFX4 BUFX4_9 ( .A(sel_B[8]), .Y(sel_B_8_bF_buf1_) );
BUFX4 BUFX4_10 ( .A(sel_B[8]), .Y(sel_B_8_bF_buf0_) );
BUFX4 BUFX4_11 ( .A(sel_B[5]), .Y(sel_B_5_bF_buf4_) );
BUFX4 BUFX4_12 ( .A(sel_B[5]), .Y(sel_B_5_bF_buf3_) );
BUFX4 BUFX4_13 ( .A(sel_B[5]), .Y(sel_B_5_bF_buf2_) );
BUFX4 BUFX4_14 ( .A(sel_B[5]), .Y(sel_B_5_bF_buf1_) );
BUFX4 BUFX4_15 ( .A(sel_B[5]), .Y(sel_B_5_bF_buf0_) );
BUFX4 BUFX4_16 ( .A(sel_A[8]), .Y(sel_A_8_bF_buf4_) );
BUFX4 BUFX4_17 ( .A(sel_A[8]), .Y(sel_A_8_bF_buf3_) );
BUFX4 BUFX4_18 ( .A(sel_A[8]), .Y(sel_A_8_bF_buf2_) );
BUFX4 BUFX4_19 ( .A(sel_A[8]), .Y(sel_A_8_bF_buf1_) );
BUFX4 BUFX4_20 ( .A(sel_A[8]), .Y(sel_A_8_bF_buf0_) );
BUFX4 BUFX4_21 ( .A(sel_B[2]), .Y(sel_B_2_bF_buf4_) );
BUFX4 BUFX4_22 ( .A(sel_B[2]), .Y(sel_B_2_bF_buf3_) );
BUFX4 BUFX4_23 ( .A(sel_B[2]), .Y(sel_B_2_bF_buf2_) );
BUFX4 BUFX4_24 ( .A(sel_B[2]), .Y(sel_B_2_bF_buf1_) );
BUFX4 BUFX4_25 ( .A(sel_B[2]), .Y(sel_B_2_bF_buf0_) );
BUFX4 BUFX4_26 ( .A(sel_A[5]), .Y(sel_A_5_bF_buf4_) );
BUFX4 BUFX4_27 ( .A(sel_A[5]), .Y(sel_A_5_bF_buf3_) );
BUFX4 BUFX4_28 ( .A(sel_A[5]), .Y(sel_A_5_bF_buf2_) );
BUFX4 BUFX4_29 ( .A(sel_A[5]), .Y(sel_A_5_bF_buf1_) );
BUFX4 BUFX4_30 ( .A(sel_A[5]), .Y(sel_A_5_bF_buf0_) );
BUFX4 BUFX4_31 ( .A(sel_A[2]), .Y(sel_A_2_bF_buf4_) );
BUFX4 BUFX4_32 ( .A(sel_A[2]), .Y(sel_A_2_bF_buf3_) );
BUFX4 BUFX4_33 ( .A(sel_A[2]), .Y(sel_A_2_bF_buf2_) );
BUFX4 BUFX4_34 ( .A(sel_A[2]), .Y(sel_A_2_bF_buf1_) );
BUFX4 BUFX4_35 ( .A(sel_A[2]), .Y(sel_A_2_bF_buf0_) );
BUFX4 BUFX4_36 ( .A(sel_B[11]), .Y(sel_B_11_bF_buf4_) );
BUFX4 BUFX4_37 ( .A(sel_B[11]), .Y(sel_B_11_bF_buf3_) );
BUFX4 BUFX4_38 ( .A(sel_B[11]), .Y(sel_B_11_bF_buf2_) );
BUFX4 BUFX4_39 ( .A(sel_B[11]), .Y(sel_B_11_bF_buf1_) );
BUFX4 BUFX4_40 ( .A(sel_B[11]), .Y(sel_B_11_bF_buf0_) );
NAND2X1 NAND2X1_1 ( .A(sel_B_8_bF_buf4_), .B(_469_), .Y(_470_) );
NAND3X1 NAND3X1_1 ( .A(_458_), .B(_468_), .C(_470_), .Y(_471_) );
INVX1 INVX1_1 ( .A(DATA_B[12]), .Y(_472_) );
NAND2X1 NAND2X1_2 ( .A(sel_B_8_bF_buf3_), .B(DATA_B[28]), .Y(_473_) );
OAI21X1 OAI21X1_1 ( .A(_472_), .B(sel_B_8_bF_buf2_), .C(_473_), .Y(_474_) );
NAND2X1 NAND2X1_3 ( .A(sel_B[7]), .B(_474_), .Y(_475_) );
NAND3X1 NAND3X1_2 ( .A(sel_B[6]), .B(_471_), .C(_475_), .Y(_476_) );
NAND3X1 NAND3X1_3 ( .A(_456_), .B(_467_), .C(_476_), .Y(_477_) );
INVX2 INVX2_1 ( .A(sel_A[6]), .Y(_320_) );
INVX4 INVX4_1 ( .A(sel_A[7]), .Y(_321_) );
OR2X2 OR2X2_1 ( .A(DATA_A[0]), .B(sel_A_8_bF_buf4_), .Y(_322_) );
INVX1 INVX1_2 ( .A(DATA_A[16]), .Y(_323_) );
NAND2X1 NAND2X1_4 ( .A(sel_A_8_bF_buf3_), .B(_323_), .Y(_324_) );
NAND3X1 NAND3X1_4 ( .A(_321_), .B(_322_), .C(_324_), .Y(_325_) );
INVX1 INVX1_3 ( .A(DATA_A[24]), .Y(_326_) );
NAND2X1 NAND2X1_5 ( .A(sel_A_8_bF_buf2_), .B(_326_), .Y(_327_) );
OR2X2 OR2X2_2 ( .A(sel_A_8_bF_buf1_), .B(DATA_A[8]), .Y(_328_) );
NAND3X1 NAND3X1_5 ( .A(sel_A[7]), .B(_328_), .C(_327_), .Y(_329_) );
NAND3X1 NAND3X1_6 ( .A(_320_), .B(_325_), .C(_329_), .Y(_330_) );
OR2X2 OR2X2_3 ( .A(sel_A_8_bF_buf0_), .B(DATA_A[4]), .Y(_331_) );
INVX1 INVX1_4 ( .A(DATA_A[20]), .Y(_332_) );
NAND2X1 NAND2X1_6 ( .A(sel_A_8_bF_buf4_), .B(_332_), .Y(_333_) );
NAND3X1 NAND3X1_7 ( .A(_321_), .B(_331_), .C(_333_), .Y(_334_) );
INVX1 INVX1_5 ( .A(DATA_A[12]), .Y(_335_) );
NAND2X1 NAND2X1_7 ( .A(sel_A_8_bF_buf3_), .B(DATA_A[28]), .Y(_336_) );
OAI21X1 OAI21X1_2 ( .A(_335_), .B(sel_A_8_bF_buf2_), .C(_336_), .Y(_337_) );
NAND2X1 NAND2X1_8 ( .A(sel_A[7]), .B(_337_), .Y(_338_) );
NAND3X1 NAND3X1_8 ( .A(sel_A[6]), .B(_334_), .C(_338_), .Y(_339_) );
NAND3X1 NAND3X1_9 ( .A(SEL[2]), .B(_330_), .C(_339_), .Y(_340_) );
AOI21X1 AOI21X1_1 ( .A(_477_), .B(_340_), .C(_455_), .Y(_319__0_) );
OR2X2 OR2X2_4 ( .A(sel_B_8_bF_buf1_), .B(DATA_B[1]), .Y(_341_) );
INVX1 INVX1_6 ( .A(DATA_B[17]), .Y(_342_) );
NAND2X1 NAND2X1_9 ( .A(sel_B_8_bF_buf0_), .B(_342_), .Y(_343_) );
NAND3X1 NAND3X1_10 ( .A(_458_), .B(_341_), .C(_343_), .Y(_344_) );
INVX1 INVX1_7 ( .A(DATA_B[25]), .Y(_345_) );
NAND2X1 NAND2X1_10 ( .A(sel_B_8_bF_buf4_), .B(_345_), .Y(_346_) );
OR2X2 OR2X2_5 ( .A(sel_B_8_bF_buf3_), .B(DATA_B[9]), .Y(_347_) );
NAND3X1 NAND3X1_11 ( .A(sel_B[7]), .B(_347_), .C(_346_), .Y(_348_) );
NAND3X1 NAND3X1_12 ( .A(_457_), .B(_344_), .C(_348_), .Y(_349_) );
OR2X2 OR2X2_6 ( .A(sel_B_8_bF_buf2_), .B(DATA_B[5]), .Y(_350_) );
INVX1 INVX1_8 ( .A(DATA_B[21]), .Y(_351_) );
NAND2X1 NAND2X1_11 ( .A(sel_B_8_bF_buf1_), .B(_351_), .Y(_352_) );
NAND3X1 NAND3X1_13 ( .A(_458_), .B(_350_), .C(_352_), .Y(_353_) );
INVX1 INVX1_9 ( .A(DATA_B[13]), .Y(_354_) );
NAND2X1 NAND2X1_12 ( .A(sel_B_8_bF_buf0_), .B(DATA_B[29]), .Y(_355_) );
OAI21X1 OAI21X1_3 ( .A(_354_), .B(sel_B_8_bF_buf4_), .C(_355_), .Y(_356_) );
NAND2X1 NAND2X1_13 ( .A(sel_B[7]), .B(_356_), .Y(_357_) );
NAND3X1 NAND3X1_14 ( .A(sel_B[6]), .B(_353_), .C(_357_), .Y(_358_) );
NAND3X1 NAND3X1_15 ( .A(_456_), .B(_349_), .C(_358_), .Y(_359_) );
OR2X2 OR2X2_7 ( .A(sel_A_8_bF_buf1_), .B(DATA_A[1]), .Y(_360_) );
INVX1 INVX1_10 ( .A(DATA_A[17]), .Y(_361_) );
NAND2X1 NAND2X1_14 ( .A(sel_A_8_bF_buf0_), .B(_361_), .Y(_362_) );
NAND3X1 NAND3X1_16 ( .A(_321_), .B(_360_), .C(_362_), .Y(_363_) );
INVX1 INVX1_11 ( .A(DATA_A[25]), .Y(_364_) );
NAND2X1 NAND2X1_15 ( .A(sel_A_8_bF_buf4_), .B(_364_), .Y(_365_) );
OR2X2 OR2X2_8 ( .A(sel_A_8_bF_buf3_), .B(DATA_A[9]), .Y(_366_) );
NAND3X1 NAND3X1_17 ( .A(sel_A[7]), .B(_366_), .C(_365_), .Y(_367_) );
NAND3X1 NAND3X1_18 ( .A(_320_), .B(_363_), .C(_367_), .Y(_368_) );
OR2X2 OR2X2_9 ( .A(sel_A_8_bF_buf2_), .B(DATA_A[5]), .Y(_369_) );
INVX1 INVX1_12 ( .A(DATA_A[21]), .Y(_370_) );
NAND2X1 NAND2X1_16 ( .A(sel_A_8_bF_buf1_), .B(_370_), .Y(_371_) );
NAND3X1 NAND3X1_19 ( .A(_321_), .B(_369_), .C(_371_), .Y(_372_) );
INVX1 INVX1_13 ( .A(DATA_A[13]), .Y(_373_) );
NAND2X1 NAND2X1_17 ( .A(sel_A_8_bF_buf0_), .B(DATA_A[29]), .Y(_374_) );
OAI21X1 OAI21X1_4 ( .A(_373_), .B(sel_A_8_bF_buf4_), .C(_374_), .Y(_375_) );
NAND2X1 NAND2X1_18 ( .A(sel_A[7]), .B(_375_), .Y(_376_) );
NAND3X1 NAND3X1_20 ( .A(sel_A[6]), .B(_372_), .C(_376_), .Y(_377_) );
NAND3X1 NAND3X1_21 ( .A(SEL[2]), .B(_368_), .C(_377_), .Y(_378_) );
AOI21X1 AOI21X1_2 ( .A(_359_), .B(_378_), .C(_455_), .Y(_319__1_) );
OR2X2 OR2X2_10 ( .A(sel_B_8_bF_buf3_), .B(DATA_B[2]), .Y(_379_) );
INVX1 INVX1_14 ( .A(DATA_B[18]), .Y(_380_) );
NAND2X1 NAND2X1_19 ( .A(sel_B_8_bF_buf2_), .B(_380_), .Y(_381_) );
NAND3X1 NAND3X1_22 ( .A(_458_), .B(_379_), .C(_381_), .Y(_382_) );
INVX1 INVX1_15 ( .A(DATA_B[26]), .Y(_383_) );
NAND2X1 NAND2X1_20 ( .A(sel_B_8_bF_buf1_), .B(_383_), .Y(_384_) );
OR2X2 OR2X2_11 ( .A(sel_B_8_bF_buf0_), .B(DATA_B[10]), .Y(_385_) );
NAND3X1 NAND3X1_23 ( .A(sel_B[7]), .B(_385_), .C(_384_), .Y(_386_) );
NAND3X1 NAND3X1_24 ( .A(_457_), .B(_382_), .C(_386_), .Y(_387_) );
OR2X2 OR2X2_12 ( .A(sel_B_8_bF_buf4_), .B(DATA_B[6]), .Y(_388_) );
INVX1 INVX1_16 ( .A(DATA_B[22]), .Y(_389_) );
NAND2X1 NAND2X1_21 ( .A(sel_B_8_bF_buf3_), .B(_389_), .Y(_390_) );
NAND3X1 NAND3X1_25 ( .A(_458_), .B(_388_), .C(_390_), .Y(_391_) );
INVX1 INVX1_17 ( .A(DATA_B[14]), .Y(_392_) );
NAND2X1 NAND2X1_22 ( .A(sel_B_8_bF_buf2_), .B(DATA_B[30]), .Y(_393_) );
OAI21X1 OAI21X1_5 ( .A(_392_), .B(sel_B_8_bF_buf1_), .C(_393_), .Y(_394_) );
NAND2X1 NAND2X1_23 ( .A(sel_B[7]), .B(_394_), .Y(_395_) );
NAND3X1 NAND3X1_26 ( .A(sel_B[6]), .B(_391_), .C(_395_), .Y(_396_) );
NAND3X1 NAND3X1_27 ( .A(_456_), .B(_387_), .C(_396_), .Y(_397_) );
OR2X2 OR2X2_13 ( .A(sel_A_8_bF_buf3_), .B(DATA_A[6]), .Y(_398_) );
INVX1 INVX1_18 ( .A(DATA_A[22]), .Y(_399_) );
NAND2X1 NAND2X1_24 ( .A(sel_A_8_bF_buf2_), .B(_399_), .Y(_400_) );
NAND3X1 NAND3X1_28 ( .A(_321_), .B(_398_), .C(_400_), .Y(_401_) );
INVX1 INVX1_19 ( .A(DATA_A[30]), .Y(_402_) );
NAND2X1 NAND2X1_25 ( .A(sel_A_8_bF_buf1_), .B(_402_), .Y(_403_) );
OR2X2 OR2X2_14 ( .A(sel_A_8_bF_buf0_), .B(DATA_A[14]), .Y(_404_) );
NAND3X1 NAND3X1_29 ( .A(sel_A[7]), .B(_404_), .C(_403_), .Y(_405_) );
NAND3X1 NAND3X1_30 ( .A(sel_A[6]), .B(_401_), .C(_405_), .Y(_406_) );
OR2X2 OR2X2_15 ( .A(sel_A_8_bF_buf4_), .B(DATA_A[2]), .Y(_407_) );
INVX1 INVX1_20 ( .A(DATA_A[18]), .Y(_408_) );
NAND2X1 NAND2X1_26 ( .A(sel_A_8_bF_buf3_), .B(_408_), .Y(_409_) );
NAND3X1 NAND3X1_31 ( .A(_321_), .B(_407_), .C(_409_), .Y(_410_) );
INVX1 INVX1_21 ( .A(DATA_A[10]), .Y(_411_) );
NAND2X1 NAND2X1_27 ( .A(sel_A_8_bF_buf2_), .B(DATA_A[26]), .Y(_412_) );
OAI21X1 OAI21X1_6 ( .A(_411_), .B(sel_A_8_bF_buf1_), .C(_412_), .Y(_413_) );
NAND2X1 NAND2X1_28 ( .A(sel_A[7]), .B(_413_), .Y(_414_) );
NAND3X1 NAND3X1_32 ( .A(_320_), .B(_410_), .C(_414_), .Y(_415_) );
NAND3X1 NAND3X1_33 ( .A(SEL[2]), .B(_406_), .C(_415_), .Y(_416_) );
AOI21X1 AOI21X1_3 ( .A(_397_), .B(_416_), .C(_455_), .Y(_319__2_) );
OR2X2 OR2X2_16 ( .A(sel_B_8_bF_buf0_), .B(DATA_B[3]), .Y(_417_) );
INVX1 INVX1_22 ( .A(DATA_B[19]), .Y(_418_) );
NAND2X1 NAND2X1_29 ( .A(sel_B_8_bF_buf4_), .B(_418_), .Y(_419_) );
NAND3X1 NAND3X1_34 ( .A(_458_), .B(_417_), .C(_419_), .Y(_420_) );
INVX1 INVX1_23 ( .A(DATA_B[27]), .Y(_421_) );
NAND2X1 NAND2X1_30 ( .A(sel_B_8_bF_buf3_), .B(_421_), .Y(_422_) );
OR2X2 OR2X2_17 ( .A(sel_B_8_bF_buf2_), .B(DATA_B[11]), .Y(_423_) );
NAND3X1 NAND3X1_35 ( .A(sel_B[7]), .B(_423_), .C(_422_), .Y(_424_) );
NAND3X1 NAND3X1_36 ( .A(_457_), .B(_420_), .C(_424_), .Y(_425_) );
OR2X2 OR2X2_18 ( .A(sel_B_8_bF_buf1_), .B(DATA_B[7]), .Y(_426_) );
INVX1 INVX1_24 ( .A(DATA_B[23]), .Y(_427_) );
NAND2X1 NAND2X1_31 ( .A(sel_B_8_bF_buf0_), .B(_427_), .Y(_428_) );
NAND3X1 NAND3X1_37 ( .A(_458_), .B(_426_), .C(_428_), .Y(_429_) );
INVX1 INVX1_25 ( .A(DATA_B[15]), .Y(_430_) );
NAND2X1 NAND2X1_32 ( .A(sel_B_8_bF_buf4_), .B(DATA_B[31]), .Y(_431_) );
OAI21X1 OAI21X1_7 ( .A(_430_), .B(sel_B_8_bF_buf3_), .C(_431_), .Y(_432_) );
NAND2X1 NAND2X1_33 ( .A(sel_B[7]), .B(_432_), .Y(_433_) );
NAND3X1 NAND3X1_38 ( .A(sel_B[6]), .B(_429_), .C(_433_), .Y(_434_) );
NAND3X1 NAND3X1_39 ( .A(_456_), .B(_425_), .C(_434_), .Y(_435_) );
OR2X2 OR2X2_19 ( .A(sel_A_8_bF_buf0_), .B(DATA_A[3]), .Y(_436_) );
INVX1 INVX1_26 ( .A(DATA_A[19]), .Y(_437_) );
NAND2X1 NAND2X1_34 ( .A(sel_A_8_bF_buf4_), .B(_437_), .Y(_438_) );
NAND3X1 NAND3X1_40 ( .A(_321_), .B(_436_), .C(_438_), .Y(_439_) );
INVX1 INVX1_27 ( .A(DATA_A[27]), .Y(_440_) );
NAND2X1 NAND2X1_35 ( .A(sel_A_8_bF_buf3_), .B(_440_), .Y(_441_) );
OR2X2 OR2X2_20 ( .A(sel_A_8_bF_buf2_), .B(DATA_A[11]), .Y(_442_) );
NAND3X1 NAND3X1_41 ( .A(sel_A[7]), .B(_442_), .C(_441_), .Y(_443_) );
NAND3X1 NAND3X1_42 ( .A(_320_), .B(_439_), .C(_443_), .Y(_444_) );
OR2X2 OR2X2_21 ( .A(sel_A_8_bF_buf1_), .B(DATA_A[7]), .Y(_445_) );
INVX1 INVX1_28 ( .A(DATA_A[23]), .Y(_446_) );
NAND2X1 NAND2X1_36 ( .A(sel_A_8_bF_buf0_), .B(_446_), .Y(_447_) );
NAND3X1 NAND3X1_43 ( .A(_321_), .B(_445_), .C(_447_), .Y(_448_) );
INVX1 INVX1_29 ( .A(DATA_A[15]), .Y(_449_) );
NAND2X1 NAND2X1_37 ( .A(sel_A_8_bF_buf4_), .B(DATA_A[31]), .Y(_450_) );
OAI21X1 OAI21X1_8 ( .A(_449_), .B(sel_A_8_bF_buf3_), .C(_450_), .Y(_451_) );
NAND2X1 NAND2X1_38 ( .A(sel_A[7]), .B(_451_), .Y(_452_) );
NAND3X1 NAND3X1_44 ( .A(sel_A[6]), .B(_448_), .C(_452_), .Y(_453_) );
NAND3X1 NAND3X1_45 ( .A(SEL[2]), .B(_444_), .C(_453_), .Y(_454_) );
AOI21X1 AOI21X1_4 ( .A(_435_), .B(_454_), .C(_455_), .Y(_319__3_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(CLK), .D(_319__0_), .Q(_0__8_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(CLK), .D(_319__1_), .Q(_0__9_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(CLK), .D(_319__2_), .Q(_0__10_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(CLK), .D(_319__3_), .Q(_0__11_) );
INVX2 INVX2_2 ( .A(RESET_L), .Y(_614_) );
INVX2 INVX2_3 ( .A(SEL[3]), .Y(_615_) );
INVX2 INVX2_4 ( .A(sel_B[9]), .Y(_616_) );
INVX4 INVX4_2 ( .A(sel_B[10]), .Y(_617_) );
OR2X2 OR2X2_22 ( .A(DATA_B[0]), .B(sel_B_11_bF_buf4_), .Y(_618_) );
INVX1 INVX1_30 ( .A(DATA_B[16]), .Y(_619_) );
NAND2X1 NAND2X1_39 ( .A(sel_B_11_bF_buf3_), .B(_619_), .Y(_620_) );
NAND3X1 NAND3X1_46 ( .A(_617_), .B(_618_), .C(_620_), .Y(_621_) );
INVX1 INVX1_31 ( .A(DATA_B[24]), .Y(_622_) );
NAND2X1 NAND2X1_40 ( .A(sel_B_11_bF_buf2_), .B(_622_), .Y(_623_) );
OR2X2 OR2X2_23 ( .A(sel_B_11_bF_buf1_), .B(DATA_B[8]), .Y(_624_) );
NAND3X1 NAND3X1_47 ( .A(sel_B[10]), .B(_624_), .C(_623_), .Y(_625_) );
NAND3X1 NAND3X1_48 ( .A(_616_), .B(_621_), .C(_625_), .Y(_626_) );
OR2X2 OR2X2_24 ( .A(sel_B_11_bF_buf0_), .B(DATA_B[4]), .Y(_627_) );
INVX1 INVX1_32 ( .A(DATA_B[20]), .Y(_628_) );
NAND2X1 NAND2X1_41 ( .A(sel_B_11_bF_buf4_), .B(_628_), .Y(_629_) );
NAND3X1 NAND3X1_49 ( .A(_617_), .B(_627_), .C(_629_), .Y(_630_) );
INVX1 INVX1_33 ( .A(DATA_B[12]), .Y(_631_) );
NAND2X1 NAND2X1_42 ( .A(sel_B_11_bF_buf3_), .B(DATA_B[28]), .Y(_632_) );
OAI21X1 OAI21X1_9 ( .A(_631_), .B(sel_B_11_bF_buf2_), .C(_632_), .Y(_633_) );
NAND2X1 NAND2X1_43 ( .A(sel_B[10]), .B(_633_), .Y(_634_) );
NAND3X1 NAND3X1_50 ( .A(sel_B[9]), .B(_630_), .C(_634_), .Y(_635_) );
NAND3X1 NAND3X1_51 ( .A(_615_), .B(_626_), .C(_635_), .Y(_636_) );
INVX2 INVX2_5 ( .A(sel_A[9]), .Y(_479_) );
INVX4 INVX4_3 ( .A(sel_A[10]), .Y(_480_) );
OR2X2 OR2X2_25 ( .A(DATA_A[0]), .B(sel_A_11_bF_buf4_), .Y(_481_) );
INVX1 INVX1_34 ( .A(DATA_A[16]), .Y(_482_) );
NAND2X1 NAND2X1_44 ( .A(sel_A_11_bF_buf3_), .B(_482_), .Y(_483_) );
NAND3X1 NAND3X1_52 ( .A(_480_), .B(_481_), .C(_483_), .Y(_484_) );
INVX1 INVX1_35 ( .A(DATA_A[24]), .Y(_485_) );
NAND2X1 NAND2X1_45 ( .A(sel_A_11_bF_buf2_), .B(_485_), .Y(_486_) );
OR2X2 OR2X2_26 ( .A(sel_A_11_bF_buf1_), .B(DATA_A[8]), .Y(_487_) );
NAND3X1 NAND3X1_53 ( .A(sel_A[10]), .B(_487_), .C(_486_), .Y(_488_) );
NAND3X1 NAND3X1_54 ( .A(_479_), .B(_484_), .C(_488_), .Y(_489_) );
OR2X2 OR2X2_27 ( .A(sel_A_11_bF_buf0_), .B(DATA_A[4]), .Y(_490_) );
INVX1 INVX1_36 ( .A(DATA_A[20]), .Y(_491_) );
NAND2X1 NAND2X1_46 ( .A(sel_A_11_bF_buf4_), .B(_491_), .Y(_492_) );
NAND3X1 NAND3X1_55 ( .A(_480_), .B(_490_), .C(_492_), .Y(_493_) );
INVX1 INVX1_37 ( .A(DATA_A[12]), .Y(_494_) );
NAND2X1 NAND2X1_47 ( .A(sel_A_11_bF_buf3_), .B(DATA_A[28]), .Y(_495_) );
OAI21X1 OAI21X1_10 ( .A(_494_), .B(sel_A_11_bF_buf2_), .C(_495_), .Y(_496_) );
NAND2X1 NAND2X1_48 ( .A(sel_A[10]), .B(_496_), .Y(_497_) );
NAND3X1 NAND3X1_56 ( .A(sel_A[9]), .B(_493_), .C(_497_), .Y(_498_) );
NAND3X1 NAND3X1_57 ( .A(SEL[3]), .B(_489_), .C(_498_), .Y(_499_) );
AOI21X1 AOI21X1_5 ( .A(_636_), .B(_499_), .C(_614_), .Y(_478__0_) );
OR2X2 OR2X2_28 ( .A(sel_B_11_bF_buf1_), .B(DATA_B[1]), .Y(_500_) );
INVX1 INVX1_38 ( .A(DATA_B[17]), .Y(_501_) );
NAND2X1 NAND2X1_49 ( .A(sel_B_11_bF_buf0_), .B(_501_), .Y(_502_) );
NAND3X1 NAND3X1_58 ( .A(_617_), .B(_500_), .C(_502_), .Y(_503_) );
INVX1 INVX1_39 ( .A(DATA_B[25]), .Y(_504_) );
NAND2X1 NAND2X1_50 ( .A(sel_B_11_bF_buf4_), .B(_504_), .Y(_505_) );
OR2X2 OR2X2_29 ( .A(sel_B_11_bF_buf3_), .B(DATA_B[9]), .Y(_506_) );
NAND3X1 NAND3X1_59 ( .A(sel_B[10]), .B(_506_), .C(_505_), .Y(_507_) );
NAND3X1 NAND3X1_60 ( .A(_616_), .B(_503_), .C(_507_), .Y(_508_) );
OR2X2 OR2X2_30 ( .A(sel_B_11_bF_buf2_), .B(DATA_B[5]), .Y(_509_) );
INVX1 INVX1_40 ( .A(DATA_B[21]), .Y(_510_) );
NAND2X1 NAND2X1_51 ( .A(sel_B_11_bF_buf1_), .B(_510_), .Y(_511_) );
NAND3X1 NAND3X1_61 ( .A(_617_), .B(_509_), .C(_511_), .Y(_512_) );
INVX1 INVX1_41 ( .A(DATA_B[13]), .Y(_513_) );
NAND2X1 NAND2X1_52 ( .A(sel_B_11_bF_buf0_), .B(DATA_B[29]), .Y(_514_) );
OAI21X1 OAI21X1_11 ( .A(_513_), .B(sel_B_11_bF_buf4_), .C(_514_), .Y(_515_) );
NAND2X1 NAND2X1_53 ( .A(sel_B[10]), .B(_515_), .Y(_516_) );
NAND3X1 NAND3X1_62 ( .A(sel_B[9]), .B(_512_), .C(_516_), .Y(_517_) );
NAND3X1 NAND3X1_63 ( .A(_615_), .B(_508_), .C(_517_), .Y(_518_) );
OR2X2 OR2X2_31 ( .A(sel_A_11_bF_buf1_), .B(DATA_A[1]), .Y(_519_) );
INVX1 INVX1_42 ( .A(DATA_A[17]), .Y(_520_) );
NAND2X1 NAND2X1_54 ( .A(sel_A_11_bF_buf0_), .B(_520_), .Y(_521_) );
NAND3X1 NAND3X1_64 ( .A(_480_), .B(_519_), .C(_521_), .Y(_522_) );
INVX1 INVX1_43 ( .A(DATA_A[25]), .Y(_523_) );
NAND2X1 NAND2X1_55 ( .A(sel_A_11_bF_buf4_), .B(_523_), .Y(_524_) );
OR2X2 OR2X2_32 ( .A(sel_A_11_bF_buf3_), .B(DATA_A[9]), .Y(_525_) );
NAND3X1 NAND3X1_65 ( .A(sel_A[10]), .B(_525_), .C(_524_), .Y(_526_) );
NAND3X1 NAND3X1_66 ( .A(_479_), .B(_522_), .C(_526_), .Y(_527_) );
OR2X2 OR2X2_33 ( .A(sel_A_11_bF_buf2_), .B(DATA_A[5]), .Y(_528_) );
INVX1 INVX1_44 ( .A(DATA_A[21]), .Y(_529_) );
NAND2X1 NAND2X1_56 ( .A(sel_A_11_bF_buf1_), .B(_529_), .Y(_530_) );
NAND3X1 NAND3X1_67 ( .A(_480_), .B(_528_), .C(_530_), .Y(_531_) );
INVX1 INVX1_45 ( .A(DATA_A[13]), .Y(_532_) );
NAND2X1 NAND2X1_57 ( .A(sel_A_11_bF_buf0_), .B(DATA_A[29]), .Y(_533_) );
OAI21X1 OAI21X1_12 ( .A(_532_), .B(sel_A_11_bF_buf4_), .C(_533_), .Y(_534_) );
NAND2X1 NAND2X1_58 ( .A(sel_A[10]), .B(_534_), .Y(_535_) );
NAND3X1 NAND3X1_68 ( .A(sel_A[9]), .B(_531_), .C(_535_), .Y(_536_) );
NAND3X1 NAND3X1_69 ( .A(SEL[3]), .B(_527_), .C(_536_), .Y(_537_) );
AOI21X1 AOI21X1_6 ( .A(_518_), .B(_537_), .C(_614_), .Y(_478__1_) );
OR2X2 OR2X2_34 ( .A(sel_B_11_bF_buf3_), .B(DATA_B[2]), .Y(_538_) );
INVX1 INVX1_46 ( .A(DATA_B[18]), .Y(_539_) );
NAND2X1 NAND2X1_59 ( .A(sel_B_11_bF_buf2_), .B(_539_), .Y(_540_) );
NAND3X1 NAND3X1_70 ( .A(_617_), .B(_538_), .C(_540_), .Y(_541_) );
INVX1 INVX1_47 ( .A(DATA_B[26]), .Y(_542_) );
NAND2X1 NAND2X1_60 ( .A(sel_B_11_bF_buf1_), .B(_542_), .Y(_543_) );
OR2X2 OR2X2_35 ( .A(sel_B_11_bF_buf0_), .B(DATA_B[10]), .Y(_544_) );
NAND3X1 NAND3X1_71 ( .A(sel_B[10]), .B(_544_), .C(_543_), .Y(_545_) );
NAND3X1 NAND3X1_72 ( .A(_616_), .B(_541_), .C(_545_), .Y(_546_) );
OR2X2 OR2X2_36 ( .A(sel_B_11_bF_buf4_), .B(DATA_B[6]), .Y(_547_) );
INVX1 INVX1_48 ( .A(DATA_B[22]), .Y(_548_) );
NAND2X1 NAND2X1_61 ( .A(sel_B_11_bF_buf3_), .B(_548_), .Y(_549_) );
NAND3X1 NAND3X1_73 ( .A(_617_), .B(_547_), .C(_549_), .Y(_550_) );
INVX1 INVX1_49 ( .A(DATA_B[14]), .Y(_551_) );
NAND2X1 NAND2X1_62 ( .A(sel_B_11_bF_buf2_), .B(DATA_B[30]), .Y(_552_) );
OAI21X1 OAI21X1_13 ( .A(_551_), .B(sel_B_11_bF_buf1_), .C(_552_), .Y(_553_) );
NAND2X1 NAND2X1_63 ( .A(sel_B[10]), .B(_553_), .Y(_554_) );
NAND3X1 NAND3X1_74 ( .A(sel_B[9]), .B(_550_), .C(_554_), .Y(_555_) );
NAND3X1 NAND3X1_75 ( .A(_615_), .B(_546_), .C(_555_), .Y(_556_) );
OR2X2 OR2X2_37 ( .A(sel_A_11_bF_buf3_), .B(DATA_A[6]), .Y(_557_) );
INVX1 INVX1_50 ( .A(DATA_A[22]), .Y(_558_) );
NAND2X1 NAND2X1_64 ( .A(sel_A_11_bF_buf2_), .B(_558_), .Y(_559_) );
NAND3X1 NAND3X1_76 ( .A(_480_), .B(_557_), .C(_559_), .Y(_560_) );
INVX1 INVX1_51 ( .A(DATA_A[30]), .Y(_561_) );
NAND2X1 NAND2X1_65 ( .A(sel_A_11_bF_buf1_), .B(_561_), .Y(_562_) );
OR2X2 OR2X2_38 ( .A(sel_A_11_bF_buf0_), .B(DATA_A[14]), .Y(_563_) );
NAND3X1 NAND3X1_77 ( .A(sel_A[10]), .B(_563_), .C(_562_), .Y(_564_) );
NAND3X1 NAND3X1_78 ( .A(sel_A[9]), .B(_560_), .C(_564_), .Y(_565_) );
OR2X2 OR2X2_39 ( .A(sel_A_11_bF_buf4_), .B(DATA_A[2]), .Y(_566_) );
INVX1 INVX1_52 ( .A(DATA_A[18]), .Y(_567_) );
NAND2X1 NAND2X1_66 ( .A(sel_A_11_bF_buf3_), .B(_567_), .Y(_568_) );
NAND3X1 NAND3X1_79 ( .A(_480_), .B(_566_), .C(_568_), .Y(_569_) );
INVX1 INVX1_53 ( .A(DATA_A[10]), .Y(_570_) );
NAND2X1 NAND2X1_67 ( .A(sel_A_11_bF_buf2_), .B(DATA_A[26]), .Y(_571_) );
OAI21X1 OAI21X1_14 ( .A(_570_), .B(sel_A_11_bF_buf1_), .C(_571_), .Y(_572_) );
NAND2X1 NAND2X1_68 ( .A(sel_A[10]), .B(_572_), .Y(_573_) );
NAND3X1 NAND3X1_80 ( .A(_479_), .B(_569_), .C(_573_), .Y(_574_) );
NAND3X1 NAND3X1_81 ( .A(SEL[3]), .B(_565_), .C(_574_), .Y(_575_) );
AOI21X1 AOI21X1_7 ( .A(_556_), .B(_575_), .C(_614_), .Y(_478__2_) );
OR2X2 OR2X2_40 ( .A(sel_B_11_bF_buf0_), .B(DATA_B[3]), .Y(_576_) );
INVX1 INVX1_54 ( .A(DATA_B[19]), .Y(_577_) );
NAND2X1 NAND2X1_69 ( .A(sel_B_11_bF_buf4_), .B(_577_), .Y(_578_) );
NAND3X1 NAND3X1_82 ( .A(_617_), .B(_576_), .C(_578_), .Y(_579_) );
INVX1 INVX1_55 ( .A(DATA_B[27]), .Y(_580_) );
NAND2X1 NAND2X1_70 ( .A(sel_B_11_bF_buf3_), .B(_580_), .Y(_581_) );
OR2X2 OR2X2_41 ( .A(sel_B_11_bF_buf2_), .B(DATA_B[11]), .Y(_582_) );
NAND3X1 NAND3X1_83 ( .A(sel_B[10]), .B(_582_), .C(_581_), .Y(_583_) );
NAND3X1 NAND3X1_84 ( .A(_616_), .B(_579_), .C(_583_), .Y(_584_) );
OR2X2 OR2X2_42 ( .A(sel_B_11_bF_buf1_), .B(DATA_B[7]), .Y(_585_) );
INVX1 INVX1_56 ( .A(DATA_B[23]), .Y(_586_) );
NAND2X1 NAND2X1_71 ( .A(sel_B_11_bF_buf0_), .B(_586_), .Y(_587_) );
NAND3X1 NAND3X1_85 ( .A(_617_), .B(_585_), .C(_587_), .Y(_588_) );
INVX1 INVX1_57 ( .A(DATA_B[15]), .Y(_589_) );
NAND2X1 NAND2X1_72 ( .A(sel_B_11_bF_buf4_), .B(DATA_B[31]), .Y(_590_) );
OAI21X1 OAI21X1_15 ( .A(_589_), .B(sel_B_11_bF_buf3_), .C(_590_), .Y(_591_) );
NAND2X1 NAND2X1_73 ( .A(sel_B[10]), .B(_591_), .Y(_592_) );
NAND3X1 NAND3X1_86 ( .A(sel_B[9]), .B(_588_), .C(_592_), .Y(_593_) );
NAND3X1 NAND3X1_87 ( .A(_615_), .B(_584_), .C(_593_), .Y(_594_) );
OR2X2 OR2X2_43 ( .A(sel_A_11_bF_buf0_), .B(DATA_A[3]), .Y(_595_) );
INVX1 INVX1_58 ( .A(DATA_A[19]), .Y(_596_) );
NAND2X1 NAND2X1_74 ( .A(sel_A_11_bF_buf4_), .B(_596_), .Y(_597_) );
NAND3X1 NAND3X1_88 ( .A(_480_), .B(_595_), .C(_597_), .Y(_598_) );
INVX1 INVX1_59 ( .A(DATA_A[27]), .Y(_599_) );
NAND2X1 NAND2X1_75 ( .A(sel_A_11_bF_buf3_), .B(_599_), .Y(_600_) );
OR2X2 OR2X2_44 ( .A(sel_A_11_bF_buf2_), .B(DATA_A[11]), .Y(_601_) );
NAND3X1 NAND3X1_89 ( .A(sel_A[10]), .B(_601_), .C(_600_), .Y(_602_) );
NAND3X1 NAND3X1_90 ( .A(_479_), .B(_598_), .C(_602_), .Y(_603_) );
OR2X2 OR2X2_45 ( .A(sel_A_11_bF_buf1_), .B(DATA_A[7]), .Y(_604_) );
INVX1 INVX1_60 ( .A(DATA_A[23]), .Y(_605_) );
NAND2X1 NAND2X1_76 ( .A(sel_A_11_bF_buf0_), .B(_605_), .Y(_606_) );
NAND3X1 NAND3X1_91 ( .A(_480_), .B(_604_), .C(_606_), .Y(_607_) );
INVX1 INVX1_61 ( .A(DATA_A[15]), .Y(_608_) );
NAND2X1 NAND2X1_77 ( .A(sel_A_11_bF_buf4_), .B(DATA_A[31]), .Y(_609_) );
OAI21X1 OAI21X1_16 ( .A(_608_), .B(sel_A_11_bF_buf3_), .C(_609_), .Y(_610_) );
NAND2X1 NAND2X1_78 ( .A(sel_A[10]), .B(_610_), .Y(_611_) );
NAND3X1 NAND3X1_92 ( .A(sel_A[9]), .B(_607_), .C(_611_), .Y(_612_) );
NAND3X1 NAND3X1_93 ( .A(SEL[3]), .B(_603_), .C(_612_), .Y(_613_) );
AOI21X1 AOI21X1_8 ( .A(_594_), .B(_613_), .C(_614_), .Y(_478__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(CLK), .D(_478__0_), .Q(_0__12_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(CLK), .D(_478__1_), .Q(_0__13_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(CLK), .D(_478__2_), .Q(_0__14_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(CLK), .D(_478__3_), .Q(_0__15_) );
BUFX2 BUFX2_1 ( .A(_0__0_), .Y(temp[0]) );
BUFX2 BUFX2_2 ( .A(_0__1_), .Y(temp[1]) );
BUFX2 BUFX2_3 ( .A(_0__2_), .Y(temp[2]) );
BUFX2 BUFX2_4 ( .A(_0__3_), .Y(temp[3]) );
BUFX2 BUFX2_5 ( .A(_0__4_), .Y(temp[4]) );
BUFX2 BUFX2_6 ( .A(_0__5_), .Y(temp[5]) );
BUFX2 BUFX2_7 ( .A(_0__6_), .Y(temp[6]) );
BUFX2 BUFX2_8 ( .A(_0__7_), .Y(temp[7]) );
BUFX2 BUFX2_9 ( .A(_0__8_), .Y(temp[8]) );
BUFX2 BUFX2_10 ( .A(_0__9_), .Y(temp[9]) );
BUFX2 BUFX2_11 ( .A(_0__10_), .Y(temp[10]) );
BUFX2 BUFX2_12 ( .A(_0__11_), .Y(temp[11]) );
BUFX2 BUFX2_13 ( .A(_0__12_), .Y(temp[12]) );
BUFX2 BUFX2_14 ( .A(_0__13_), .Y(temp[13]) );
BUFX2 BUFX2_15 ( .A(_0__14_), .Y(temp[14]) );
BUFX2 BUFX2_16 ( .A(_0__15_), .Y(temp[15]) );
INVX2 INVX2_6 ( .A(RESET_L), .Y(_137_) );
INVX2 INVX2_7 ( .A(SEL[0]), .Y(_138_) );
INVX2 INVX2_8 ( .A(sel_B[0]), .Y(_139_) );
INVX4 INVX4_4 ( .A(sel_B[1]), .Y(_140_) );
OR2X2 OR2X2_46 ( .A(DATA_B[0]), .B(sel_B_2_bF_buf4_), .Y(_141_) );
INVX1 INVX1_62 ( .A(DATA_B[16]), .Y(_142_) );
NAND2X1 NAND2X1_79 ( .A(sel_B_2_bF_buf3_), .B(_142_), .Y(_143_) );
NAND3X1 NAND3X1_94 ( .A(_140_), .B(_141_), .C(_143_), .Y(_144_) );
INVX1 INVX1_63 ( .A(DATA_B[24]), .Y(_145_) );
NAND2X1 NAND2X1_80 ( .A(sel_B_2_bF_buf2_), .B(_145_), .Y(_146_) );
OR2X2 OR2X2_47 ( .A(sel_B_2_bF_buf1_), .B(DATA_B[8]), .Y(_147_) );
NAND3X1 NAND3X1_95 ( .A(sel_B[1]), .B(_147_), .C(_146_), .Y(_148_) );
NAND3X1 NAND3X1_96 ( .A(_139_), .B(_144_), .C(_148_), .Y(_149_) );
OR2X2 OR2X2_48 ( .A(sel_B_2_bF_buf0_), .B(DATA_B[4]), .Y(_150_) );
INVX1 INVX1_64 ( .A(DATA_B[20]), .Y(_151_) );
NAND2X1 NAND2X1_81 ( .A(sel_B_2_bF_buf4_), .B(_151_), .Y(_152_) );
NAND3X1 NAND3X1_97 ( .A(_140_), .B(_150_), .C(_152_), .Y(_153_) );
INVX1 INVX1_65 ( .A(DATA_B[12]), .Y(_154_) );
NAND2X1 NAND2X1_82 ( .A(sel_B_2_bF_buf3_), .B(DATA_B[28]), .Y(_155_) );
OAI21X1 OAI21X1_17 ( .A(_154_), .B(sel_B_2_bF_buf2_), .C(_155_), .Y(_156_) );
NAND2X1 NAND2X1_83 ( .A(sel_B[1]), .B(_156_), .Y(_157_) );
NAND3X1 NAND3X1_98 ( .A(sel_B[0]), .B(_153_), .C(_157_), .Y(_158_) );
NAND3X1 NAND3X1_99 ( .A(_138_), .B(_149_), .C(_158_), .Y(_159_) );
INVX2 INVX2_9 ( .A(sel_A[0]), .Y(_2_) );
INVX4 INVX4_5 ( .A(sel_A[1]), .Y(_3_) );
OR2X2 OR2X2_49 ( .A(DATA_A[0]), .B(sel_A_2_bF_buf4_), .Y(_4_) );
INVX1 INVX1_66 ( .A(DATA_A[16]), .Y(_5_) );
NAND2X1 NAND2X1_84 ( .A(sel_A_2_bF_buf3_), .B(_5_), .Y(_6_) );
NAND3X1 NAND3X1_100 ( .A(_3_), .B(_4_), .C(_6_), .Y(_7_) );
INVX1 INVX1_67 ( .A(DATA_A[24]), .Y(_8_) );
NAND2X1 NAND2X1_85 ( .A(sel_A_2_bF_buf2_), .B(_8_), .Y(_9_) );
OR2X2 OR2X2_50 ( .A(sel_A_2_bF_buf1_), .B(DATA_A[8]), .Y(_10_) );
NAND3X1 NAND3X1_101 ( .A(sel_A[1]), .B(_10_), .C(_9_), .Y(_11_) );
NAND3X1 NAND3X1_102 ( .A(_2_), .B(_7_), .C(_11_), .Y(_12_) );
OR2X2 OR2X2_51 ( .A(sel_A_2_bF_buf0_), .B(DATA_A[4]), .Y(_13_) );
INVX1 INVX1_68 ( .A(DATA_A[20]), .Y(_14_) );
NAND2X1 NAND2X1_86 ( .A(sel_A_2_bF_buf4_), .B(_14_), .Y(_15_) );
NAND3X1 NAND3X1_103 ( .A(_3_), .B(_13_), .C(_15_), .Y(_16_) );
INVX1 INVX1_69 ( .A(DATA_A[12]), .Y(_17_) );
NAND2X1 NAND2X1_87 ( .A(sel_A_2_bF_buf3_), .B(DATA_A[28]), .Y(_18_) );
OAI21X1 OAI21X1_18 ( .A(_17_), .B(sel_A_2_bF_buf2_), .C(_18_), .Y(_19_) );
NAND2X1 NAND2X1_88 ( .A(sel_A[1]), .B(_19_), .Y(_20_) );
NAND3X1 NAND3X1_104 ( .A(sel_A[0]), .B(_16_), .C(_20_), .Y(_21_) );
NAND3X1 NAND3X1_105 ( .A(SEL[0]), .B(_12_), .C(_21_), .Y(_22_) );
AOI21X1 AOI21X1_9 ( .A(_159_), .B(_22_), .C(_137_), .Y(_1__0_) );
OR2X2 OR2X2_52 ( .A(sel_B_2_bF_buf1_), .B(DATA_B[1]), .Y(_23_) );
INVX1 INVX1_70 ( .A(DATA_B[17]), .Y(_24_) );
NAND2X1 NAND2X1_89 ( .A(sel_B_2_bF_buf0_), .B(_24_), .Y(_25_) );
NAND3X1 NAND3X1_106 ( .A(_140_), .B(_23_), .C(_25_), .Y(_26_) );
INVX1 INVX1_71 ( .A(DATA_B[25]), .Y(_27_) );
NAND2X1 NAND2X1_90 ( .A(sel_B_2_bF_buf4_), .B(_27_), .Y(_28_) );
OR2X2 OR2X2_53 ( .A(sel_B_2_bF_buf3_), .B(DATA_B[9]), .Y(_29_) );
NAND3X1 NAND3X1_107 ( .A(sel_B[1]), .B(_29_), .C(_28_), .Y(_30_) );
NAND3X1 NAND3X1_108 ( .A(_139_), .B(_26_), .C(_30_), .Y(_31_) );
OR2X2 OR2X2_54 ( .A(sel_B_2_bF_buf2_), .B(DATA_B[5]), .Y(_32_) );
INVX1 INVX1_72 ( .A(DATA_B[21]), .Y(_33_) );
NAND2X1 NAND2X1_91 ( .A(sel_B_2_bF_buf1_), .B(_33_), .Y(_34_) );
NAND3X1 NAND3X1_109 ( .A(_140_), .B(_32_), .C(_34_), .Y(_35_) );
INVX1 INVX1_73 ( .A(DATA_B[13]), .Y(_36_) );
NAND2X1 NAND2X1_92 ( .A(sel_B_2_bF_buf0_), .B(DATA_B[29]), .Y(_37_) );
OAI21X1 OAI21X1_19 ( .A(_36_), .B(sel_B_2_bF_buf4_), .C(_37_), .Y(_38_) );
NAND2X1 NAND2X1_93 ( .A(sel_B[1]), .B(_38_), .Y(_39_) );
NAND3X1 NAND3X1_110 ( .A(sel_B[0]), .B(_35_), .C(_39_), .Y(_40_) );
NAND3X1 NAND3X1_111 ( .A(_138_), .B(_31_), .C(_40_), .Y(_41_) );
OR2X2 OR2X2_55 ( .A(sel_A_2_bF_buf1_), .B(DATA_A[1]), .Y(_42_) );
INVX1 INVX1_74 ( .A(DATA_A[17]), .Y(_43_) );
NAND2X1 NAND2X1_94 ( .A(sel_A_2_bF_buf0_), .B(_43_), .Y(_44_) );
NAND3X1 NAND3X1_112 ( .A(_3_), .B(_42_), .C(_44_), .Y(_45_) );
INVX1 INVX1_75 ( .A(DATA_A[25]), .Y(_46_) );
NAND2X1 NAND2X1_95 ( .A(sel_A_2_bF_buf4_), .B(_46_), .Y(_47_) );
OR2X2 OR2X2_56 ( .A(sel_A_2_bF_buf3_), .B(DATA_A[9]), .Y(_48_) );
NAND3X1 NAND3X1_113 ( .A(sel_A[1]), .B(_48_), .C(_47_), .Y(_49_) );
NAND3X1 NAND3X1_114 ( .A(_2_), .B(_45_), .C(_49_), .Y(_50_) );
OR2X2 OR2X2_57 ( .A(sel_A_2_bF_buf2_), .B(DATA_A[5]), .Y(_51_) );
INVX1 INVX1_76 ( .A(DATA_A[21]), .Y(_52_) );
NAND2X1 NAND2X1_96 ( .A(sel_A_2_bF_buf1_), .B(_52_), .Y(_53_) );
NAND3X1 NAND3X1_115 ( .A(_3_), .B(_51_), .C(_53_), .Y(_54_) );
INVX1 INVX1_77 ( .A(DATA_A[13]), .Y(_55_) );
NAND2X1 NAND2X1_97 ( .A(sel_A_2_bF_buf0_), .B(DATA_A[29]), .Y(_56_) );
OAI21X1 OAI21X1_20 ( .A(_55_), .B(sel_A_2_bF_buf4_), .C(_56_), .Y(_57_) );
NAND2X1 NAND2X1_98 ( .A(sel_A[1]), .B(_57_), .Y(_58_) );
NAND3X1 NAND3X1_116 ( .A(sel_A[0]), .B(_54_), .C(_58_), .Y(_59_) );
NAND3X1 NAND3X1_117 ( .A(SEL[0]), .B(_50_), .C(_59_), .Y(_60_) );
AOI21X1 AOI21X1_10 ( .A(_41_), .B(_60_), .C(_137_), .Y(_1__1_) );
OR2X2 OR2X2_58 ( .A(sel_B_2_bF_buf3_), .B(DATA_B[2]), .Y(_61_) );
INVX1 INVX1_78 ( .A(DATA_B[18]), .Y(_62_) );
NAND2X1 NAND2X1_99 ( .A(sel_B_2_bF_buf2_), .B(_62_), .Y(_63_) );
NAND3X1 NAND3X1_118 ( .A(_140_), .B(_61_), .C(_63_), .Y(_64_) );
INVX1 INVX1_79 ( .A(DATA_B[26]), .Y(_65_) );
NAND2X1 NAND2X1_100 ( .A(sel_B_2_bF_buf1_), .B(_65_), .Y(_66_) );
OR2X2 OR2X2_59 ( .A(sel_B_2_bF_buf0_), .B(DATA_B[10]), .Y(_67_) );
NAND3X1 NAND3X1_119 ( .A(sel_B[1]), .B(_67_), .C(_66_), .Y(_68_) );
NAND3X1 NAND3X1_120 ( .A(_139_), .B(_64_), .C(_68_), .Y(_69_) );
OR2X2 OR2X2_60 ( .A(sel_B_2_bF_buf4_), .B(DATA_B[6]), .Y(_70_) );
INVX1 INVX1_80 ( .A(DATA_B[22]), .Y(_71_) );
NAND2X1 NAND2X1_101 ( .A(sel_B_2_bF_buf3_), .B(_71_), .Y(_72_) );
NAND3X1 NAND3X1_121 ( .A(_140_), .B(_70_), .C(_72_), .Y(_73_) );
INVX1 INVX1_81 ( .A(DATA_B[14]), .Y(_74_) );
NAND2X1 NAND2X1_102 ( .A(sel_B_2_bF_buf2_), .B(DATA_B[30]), .Y(_75_) );
OAI21X1 OAI21X1_21 ( .A(_74_), .B(sel_B_2_bF_buf1_), .C(_75_), .Y(_76_) );
NAND2X1 NAND2X1_103 ( .A(sel_B[1]), .B(_76_), .Y(_77_) );
NAND3X1 NAND3X1_122 ( .A(sel_B[0]), .B(_73_), .C(_77_), .Y(_78_) );
NAND3X1 NAND3X1_123 ( .A(_138_), .B(_69_), .C(_78_), .Y(_79_) );
OR2X2 OR2X2_61 ( .A(sel_A_2_bF_buf3_), .B(DATA_A[6]), .Y(_80_) );
INVX1 INVX1_82 ( .A(DATA_A[22]), .Y(_81_) );
NAND2X1 NAND2X1_104 ( .A(sel_A_2_bF_buf2_), .B(_81_), .Y(_82_) );
NAND3X1 NAND3X1_124 ( .A(_3_), .B(_80_), .C(_82_), .Y(_83_) );
INVX1 INVX1_83 ( .A(DATA_A[30]), .Y(_84_) );
NAND2X1 NAND2X1_105 ( .A(sel_A_2_bF_buf1_), .B(_84_), .Y(_85_) );
OR2X2 OR2X2_62 ( .A(sel_A_2_bF_buf0_), .B(DATA_A[14]), .Y(_86_) );
NAND3X1 NAND3X1_125 ( .A(sel_A[1]), .B(_86_), .C(_85_), .Y(_87_) );
NAND3X1 NAND3X1_126 ( .A(sel_A[0]), .B(_83_), .C(_87_), .Y(_88_) );
OR2X2 OR2X2_63 ( .A(sel_A_2_bF_buf4_), .B(DATA_A[2]), .Y(_89_) );
INVX1 INVX1_84 ( .A(DATA_A[18]), .Y(_90_) );
NAND2X1 NAND2X1_106 ( .A(sel_A_2_bF_buf3_), .B(_90_), .Y(_91_) );
NAND3X1 NAND3X1_127 ( .A(_3_), .B(_89_), .C(_91_), .Y(_92_) );
INVX1 INVX1_85 ( .A(DATA_A[10]), .Y(_93_) );
NAND2X1 NAND2X1_107 ( .A(sel_A_2_bF_buf2_), .B(DATA_A[26]), .Y(_94_) );
OAI21X1 OAI21X1_22 ( .A(_93_), .B(sel_A_2_bF_buf1_), .C(_94_), .Y(_95_) );
NAND2X1 NAND2X1_108 ( .A(sel_A[1]), .B(_95_), .Y(_96_) );
NAND3X1 NAND3X1_128 ( .A(_2_), .B(_92_), .C(_96_), .Y(_97_) );
NAND3X1 NAND3X1_129 ( .A(SEL[0]), .B(_88_), .C(_97_), .Y(_98_) );
AOI21X1 AOI21X1_11 ( .A(_79_), .B(_98_), .C(_137_), .Y(_1__2_) );
OR2X2 OR2X2_64 ( .A(sel_B_2_bF_buf0_), .B(DATA_B[3]), .Y(_99_) );
INVX1 INVX1_86 ( .A(DATA_B[19]), .Y(_100_) );
NAND2X1 NAND2X1_109 ( .A(sel_B_2_bF_buf4_), .B(_100_), .Y(_101_) );
NAND3X1 NAND3X1_130 ( .A(_140_), .B(_99_), .C(_101_), .Y(_102_) );
INVX1 INVX1_87 ( .A(DATA_B[27]), .Y(_103_) );
NAND2X1 NAND2X1_110 ( .A(sel_B_2_bF_buf3_), .B(_103_), .Y(_104_) );
OR2X2 OR2X2_65 ( .A(sel_B_2_bF_buf2_), .B(DATA_B[11]), .Y(_105_) );
NAND3X1 NAND3X1_131 ( .A(sel_B[1]), .B(_105_), .C(_104_), .Y(_106_) );
NAND3X1 NAND3X1_132 ( .A(_139_), .B(_102_), .C(_106_), .Y(_107_) );
OR2X2 OR2X2_66 ( .A(sel_B_2_bF_buf1_), .B(DATA_B[7]), .Y(_108_) );
INVX1 INVX1_88 ( .A(DATA_B[23]), .Y(_109_) );
NAND2X1 NAND2X1_111 ( .A(sel_B_2_bF_buf0_), .B(_109_), .Y(_110_) );
NAND3X1 NAND3X1_133 ( .A(_140_), .B(_108_), .C(_110_), .Y(_111_) );
INVX1 INVX1_89 ( .A(DATA_B[15]), .Y(_112_) );
NAND2X1 NAND2X1_112 ( .A(sel_B_2_bF_buf4_), .B(DATA_B[31]), .Y(_113_) );
OAI21X1 OAI21X1_23 ( .A(_112_), .B(sel_B_2_bF_buf3_), .C(_113_), .Y(_114_) );
NAND2X1 NAND2X1_113 ( .A(sel_B[1]), .B(_114_), .Y(_115_) );
NAND3X1 NAND3X1_134 ( .A(sel_B[0]), .B(_111_), .C(_115_), .Y(_116_) );
NAND3X1 NAND3X1_135 ( .A(_138_), .B(_107_), .C(_116_), .Y(_117_) );
OR2X2 OR2X2_67 ( .A(sel_A_2_bF_buf0_), .B(DATA_A[3]), .Y(_118_) );
INVX1 INVX1_90 ( .A(DATA_A[19]), .Y(_119_) );
NAND2X1 NAND2X1_114 ( .A(sel_A_2_bF_buf4_), .B(_119_), .Y(_120_) );
NAND3X1 NAND3X1_136 ( .A(_3_), .B(_118_), .C(_120_), .Y(_121_) );
INVX1 INVX1_91 ( .A(DATA_A[27]), .Y(_122_) );
NAND2X1 NAND2X1_115 ( .A(sel_A_2_bF_buf3_), .B(_122_), .Y(_123_) );
OR2X2 OR2X2_68 ( .A(sel_A_2_bF_buf2_), .B(DATA_A[11]), .Y(_124_) );
NAND3X1 NAND3X1_137 ( .A(sel_A[1]), .B(_124_), .C(_123_), .Y(_125_) );
NAND3X1 NAND3X1_138 ( .A(_2_), .B(_121_), .C(_125_), .Y(_126_) );
OR2X2 OR2X2_69 ( .A(sel_A_2_bF_buf1_), .B(DATA_A[7]), .Y(_127_) );
INVX1 INVX1_92 ( .A(DATA_A[23]), .Y(_128_) );
NAND2X1 NAND2X1_116 ( .A(sel_A_2_bF_buf0_), .B(_128_), .Y(_129_) );
NAND3X1 NAND3X1_139 ( .A(_3_), .B(_127_), .C(_129_), .Y(_130_) );
INVX1 INVX1_93 ( .A(DATA_A[15]), .Y(_131_) );
NAND2X1 NAND2X1_117 ( .A(sel_A_2_bF_buf4_), .B(DATA_A[31]), .Y(_132_) );
OAI21X1 OAI21X1_24 ( .A(_131_), .B(sel_A_2_bF_buf3_), .C(_132_), .Y(_133_) );
NAND2X1 NAND2X1_118 ( .A(sel_A[1]), .B(_133_), .Y(_134_) );
NAND3X1 NAND3X1_140 ( .A(sel_A[0]), .B(_130_), .C(_134_), .Y(_135_) );
NAND3X1 NAND3X1_141 ( .A(SEL[0]), .B(_126_), .C(_135_), .Y(_136_) );
AOI21X1 AOI21X1_12 ( .A(_117_), .B(_136_), .C(_137_), .Y(_1__3_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(CLK), .D(_1__0_), .Q(_0__0_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(CLK), .D(_1__1_), .Q(_0__1_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(CLK), .D(_1__2_), .Q(_0__2_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(CLK), .D(_1__3_), .Q(_0__3_) );
INVX2 INVX2_10 ( .A(RESET_L), .Y(_296_) );
INVX2 INVX2_11 ( .A(SEL[1]), .Y(_297_) );
INVX2 INVX2_12 ( .A(sel_B[3]), .Y(_298_) );
INVX4 INVX4_6 ( .A(sel_B[4]), .Y(_299_) );
OR2X2 OR2X2_70 ( .A(DATA_B[0]), .B(sel_B_5_bF_buf4_), .Y(_300_) );
INVX1 INVX1_94 ( .A(DATA_B[16]), .Y(_301_) );
NAND2X1 NAND2X1_119 ( .A(sel_B_5_bF_buf3_), .B(_301_), .Y(_302_) );
NAND3X1 NAND3X1_142 ( .A(_299_), .B(_300_), .C(_302_), .Y(_303_) );
INVX1 INVX1_95 ( .A(DATA_B[24]), .Y(_304_) );
NAND2X1 NAND2X1_120 ( .A(sel_B_5_bF_buf2_), .B(_304_), .Y(_305_) );
OR2X2 OR2X2_71 ( .A(sel_B_5_bF_buf1_), .B(DATA_B[8]), .Y(_306_) );
NAND3X1 NAND3X1_143 ( .A(sel_B[4]), .B(_306_), .C(_305_), .Y(_307_) );
NAND3X1 NAND3X1_144 ( .A(_298_), .B(_303_), .C(_307_), .Y(_308_) );
OR2X2 OR2X2_72 ( .A(sel_B_5_bF_buf0_), .B(DATA_B[4]), .Y(_309_) );
INVX1 INVX1_96 ( .A(DATA_B[20]), .Y(_310_) );
NAND2X1 NAND2X1_121 ( .A(sel_B_5_bF_buf4_), .B(_310_), .Y(_311_) );
NAND3X1 NAND3X1_145 ( .A(_299_), .B(_309_), .C(_311_), .Y(_312_) );
INVX1 INVX1_97 ( .A(DATA_B[12]), .Y(_313_) );
NAND2X1 NAND2X1_122 ( .A(sel_B_5_bF_buf3_), .B(DATA_B[28]), .Y(_314_) );
OAI21X1 OAI21X1_25 ( .A(_313_), .B(sel_B_5_bF_buf2_), .C(_314_), .Y(_315_) );
NAND2X1 NAND2X1_123 ( .A(sel_B[4]), .B(_315_), .Y(_316_) );
NAND3X1 NAND3X1_146 ( .A(sel_B[3]), .B(_312_), .C(_316_), .Y(_317_) );
NAND3X1 NAND3X1_147 ( .A(_297_), .B(_308_), .C(_317_), .Y(_318_) );
INVX2 INVX2_13 ( .A(sel_A[3]), .Y(_161_) );
INVX4 INVX4_7 ( .A(sel_A[4]), .Y(_162_) );
OR2X2 OR2X2_73 ( .A(DATA_A[0]), .B(sel_A_5_bF_buf4_), .Y(_163_) );
INVX1 INVX1_98 ( .A(DATA_A[16]), .Y(_164_) );
NAND2X1 NAND2X1_124 ( .A(sel_A_5_bF_buf3_), .B(_164_), .Y(_165_) );
NAND3X1 NAND3X1_148 ( .A(_162_), .B(_163_), .C(_165_), .Y(_166_) );
INVX1 INVX1_99 ( .A(DATA_A[24]), .Y(_167_) );
NAND2X1 NAND2X1_125 ( .A(sel_A_5_bF_buf2_), .B(_167_), .Y(_168_) );
OR2X2 OR2X2_74 ( .A(sel_A_5_bF_buf1_), .B(DATA_A[8]), .Y(_169_) );
NAND3X1 NAND3X1_149 ( .A(sel_A[4]), .B(_169_), .C(_168_), .Y(_170_) );
NAND3X1 NAND3X1_150 ( .A(_161_), .B(_166_), .C(_170_), .Y(_171_) );
OR2X2 OR2X2_75 ( .A(sel_A_5_bF_buf0_), .B(DATA_A[4]), .Y(_172_) );
INVX1 INVX1_100 ( .A(DATA_A[20]), .Y(_173_) );
NAND2X1 NAND2X1_126 ( .A(sel_A_5_bF_buf4_), .B(_173_), .Y(_174_) );
NAND3X1 NAND3X1_151 ( .A(_162_), .B(_172_), .C(_174_), .Y(_175_) );
INVX1 INVX1_101 ( .A(DATA_A[12]), .Y(_176_) );
NAND2X1 NAND2X1_127 ( .A(sel_A_5_bF_buf3_), .B(DATA_A[28]), .Y(_177_) );
OAI21X1 OAI21X1_26 ( .A(_176_), .B(sel_A_5_bF_buf2_), .C(_177_), .Y(_178_) );
NAND2X1 NAND2X1_128 ( .A(sel_A[4]), .B(_178_), .Y(_179_) );
NAND3X1 NAND3X1_152 ( .A(sel_A[3]), .B(_175_), .C(_179_), .Y(_180_) );
NAND3X1 NAND3X1_153 ( .A(SEL[1]), .B(_171_), .C(_180_), .Y(_181_) );
AOI21X1 AOI21X1_13 ( .A(_318_), .B(_181_), .C(_296_), .Y(_160__0_) );
OR2X2 OR2X2_76 ( .A(sel_B_5_bF_buf1_), .B(DATA_B[1]), .Y(_182_) );
INVX1 INVX1_102 ( .A(DATA_B[17]), .Y(_183_) );
NAND2X1 NAND2X1_129 ( .A(sel_B_5_bF_buf0_), .B(_183_), .Y(_184_) );
NAND3X1 NAND3X1_154 ( .A(_299_), .B(_182_), .C(_184_), .Y(_185_) );
INVX1 INVX1_103 ( .A(DATA_B[25]), .Y(_186_) );
NAND2X1 NAND2X1_130 ( .A(sel_B_5_bF_buf4_), .B(_186_), .Y(_187_) );
OR2X2 OR2X2_77 ( .A(sel_B_5_bF_buf3_), .B(DATA_B[9]), .Y(_188_) );
NAND3X1 NAND3X1_155 ( .A(sel_B[4]), .B(_188_), .C(_187_), .Y(_189_) );
NAND3X1 NAND3X1_156 ( .A(_298_), .B(_185_), .C(_189_), .Y(_190_) );
OR2X2 OR2X2_78 ( .A(sel_B_5_bF_buf2_), .B(DATA_B[5]), .Y(_191_) );
INVX1 INVX1_104 ( .A(DATA_B[21]), .Y(_192_) );
NAND2X1 NAND2X1_131 ( .A(sel_B_5_bF_buf1_), .B(_192_), .Y(_193_) );
NAND3X1 NAND3X1_157 ( .A(_299_), .B(_191_), .C(_193_), .Y(_194_) );
INVX1 INVX1_105 ( .A(DATA_B[13]), .Y(_195_) );
NAND2X1 NAND2X1_132 ( .A(sel_B_5_bF_buf0_), .B(DATA_B[29]), .Y(_196_) );
OAI21X1 OAI21X1_27 ( .A(_195_), .B(sel_B_5_bF_buf4_), .C(_196_), .Y(_197_) );
NAND2X1 NAND2X1_133 ( .A(sel_B[4]), .B(_197_), .Y(_198_) );
NAND3X1 NAND3X1_158 ( .A(sel_B[3]), .B(_194_), .C(_198_), .Y(_199_) );
NAND3X1 NAND3X1_159 ( .A(_297_), .B(_190_), .C(_199_), .Y(_200_) );
OR2X2 OR2X2_79 ( .A(sel_A_5_bF_buf1_), .B(DATA_A[1]), .Y(_201_) );
INVX1 INVX1_106 ( .A(DATA_A[17]), .Y(_202_) );
NAND2X1 NAND2X1_134 ( .A(sel_A_5_bF_buf0_), .B(_202_), .Y(_203_) );
NAND3X1 NAND3X1_160 ( .A(_162_), .B(_201_), .C(_203_), .Y(_204_) );
INVX1 INVX1_107 ( .A(DATA_A[25]), .Y(_205_) );
NAND2X1 NAND2X1_135 ( .A(sel_A_5_bF_buf4_), .B(_205_), .Y(_206_) );
OR2X2 OR2X2_80 ( .A(sel_A_5_bF_buf3_), .B(DATA_A[9]), .Y(_207_) );
NAND3X1 NAND3X1_161 ( .A(sel_A[4]), .B(_207_), .C(_206_), .Y(_208_) );
NAND3X1 NAND3X1_162 ( .A(_161_), .B(_204_), .C(_208_), .Y(_209_) );
OR2X2 OR2X2_81 ( .A(sel_A_5_bF_buf2_), .B(DATA_A[5]), .Y(_210_) );
INVX1 INVX1_108 ( .A(DATA_A[21]), .Y(_211_) );
NAND2X1 NAND2X1_136 ( .A(sel_A_5_bF_buf1_), .B(_211_), .Y(_212_) );
NAND3X1 NAND3X1_163 ( .A(_162_), .B(_210_), .C(_212_), .Y(_213_) );
INVX1 INVX1_109 ( .A(DATA_A[13]), .Y(_214_) );
NAND2X1 NAND2X1_137 ( .A(sel_A_5_bF_buf0_), .B(DATA_A[29]), .Y(_215_) );
OAI21X1 OAI21X1_28 ( .A(_214_), .B(sel_A_5_bF_buf4_), .C(_215_), .Y(_216_) );
NAND2X1 NAND2X1_138 ( .A(sel_A[4]), .B(_216_), .Y(_217_) );
NAND3X1 NAND3X1_164 ( .A(sel_A[3]), .B(_213_), .C(_217_), .Y(_218_) );
NAND3X1 NAND3X1_165 ( .A(SEL[1]), .B(_209_), .C(_218_), .Y(_219_) );
AOI21X1 AOI21X1_14 ( .A(_200_), .B(_219_), .C(_296_), .Y(_160__1_) );
OR2X2 OR2X2_82 ( .A(sel_B_5_bF_buf3_), .B(DATA_B[2]), .Y(_220_) );
INVX1 INVX1_110 ( .A(DATA_B[18]), .Y(_221_) );
NAND2X1 NAND2X1_139 ( .A(sel_B_5_bF_buf2_), .B(_221_), .Y(_222_) );
NAND3X1 NAND3X1_166 ( .A(_299_), .B(_220_), .C(_222_), .Y(_223_) );
INVX1 INVX1_111 ( .A(DATA_B[26]), .Y(_224_) );
NAND2X1 NAND2X1_140 ( .A(sel_B_5_bF_buf1_), .B(_224_), .Y(_225_) );
OR2X2 OR2X2_83 ( .A(sel_B_5_bF_buf0_), .B(DATA_B[10]), .Y(_226_) );
NAND3X1 NAND3X1_167 ( .A(sel_B[4]), .B(_226_), .C(_225_), .Y(_227_) );
NAND3X1 NAND3X1_168 ( .A(_298_), .B(_223_), .C(_227_), .Y(_228_) );
OR2X2 OR2X2_84 ( .A(sel_B_5_bF_buf4_), .B(DATA_B[6]), .Y(_229_) );
INVX1 INVX1_112 ( .A(DATA_B[22]), .Y(_230_) );
NAND2X1 NAND2X1_141 ( .A(sel_B_5_bF_buf3_), .B(_230_), .Y(_231_) );
NAND3X1 NAND3X1_169 ( .A(_299_), .B(_229_), .C(_231_), .Y(_232_) );
INVX1 INVX1_113 ( .A(DATA_B[14]), .Y(_233_) );
NAND2X1 NAND2X1_142 ( .A(sel_B_5_bF_buf2_), .B(DATA_B[30]), .Y(_234_) );
OAI21X1 OAI21X1_29 ( .A(_233_), .B(sel_B_5_bF_buf1_), .C(_234_), .Y(_235_) );
NAND2X1 NAND2X1_143 ( .A(sel_B[4]), .B(_235_), .Y(_236_) );
NAND3X1 NAND3X1_170 ( .A(sel_B[3]), .B(_232_), .C(_236_), .Y(_237_) );
NAND3X1 NAND3X1_171 ( .A(_297_), .B(_228_), .C(_237_), .Y(_238_) );
OR2X2 OR2X2_85 ( .A(sel_A_5_bF_buf3_), .B(DATA_A[6]), .Y(_239_) );
INVX1 INVX1_114 ( .A(DATA_A[22]), .Y(_240_) );
NAND2X1 NAND2X1_144 ( .A(sel_A_5_bF_buf2_), .B(_240_), .Y(_241_) );
NAND3X1 NAND3X1_172 ( .A(_162_), .B(_239_), .C(_241_), .Y(_242_) );
INVX1 INVX1_115 ( .A(DATA_A[30]), .Y(_243_) );
NAND2X1 NAND2X1_145 ( .A(sel_A_5_bF_buf1_), .B(_243_), .Y(_244_) );
OR2X2 OR2X2_86 ( .A(sel_A_5_bF_buf0_), .B(DATA_A[14]), .Y(_245_) );
NAND3X1 NAND3X1_173 ( .A(sel_A[4]), .B(_245_), .C(_244_), .Y(_246_) );
NAND3X1 NAND3X1_174 ( .A(sel_A[3]), .B(_242_), .C(_246_), .Y(_247_) );
OR2X2 OR2X2_87 ( .A(sel_A_5_bF_buf4_), .B(DATA_A[2]), .Y(_248_) );
INVX1 INVX1_116 ( .A(DATA_A[18]), .Y(_249_) );
NAND2X1 NAND2X1_146 ( .A(sel_A_5_bF_buf3_), .B(_249_), .Y(_250_) );
NAND3X1 NAND3X1_175 ( .A(_162_), .B(_248_), .C(_250_), .Y(_251_) );
INVX1 INVX1_117 ( .A(DATA_A[10]), .Y(_252_) );
NAND2X1 NAND2X1_147 ( .A(sel_A_5_bF_buf2_), .B(DATA_A[26]), .Y(_253_) );
OAI21X1 OAI21X1_30 ( .A(_252_), .B(sel_A_5_bF_buf1_), .C(_253_), .Y(_254_) );
NAND2X1 NAND2X1_148 ( .A(sel_A[4]), .B(_254_), .Y(_255_) );
NAND3X1 NAND3X1_176 ( .A(_161_), .B(_251_), .C(_255_), .Y(_256_) );
NAND3X1 NAND3X1_177 ( .A(SEL[1]), .B(_247_), .C(_256_), .Y(_257_) );
AOI21X1 AOI21X1_15 ( .A(_238_), .B(_257_), .C(_296_), .Y(_160__2_) );
OR2X2 OR2X2_88 ( .A(sel_B_5_bF_buf0_), .B(DATA_B[3]), .Y(_258_) );
INVX1 INVX1_118 ( .A(DATA_B[19]), .Y(_259_) );
NAND2X1 NAND2X1_149 ( .A(sel_B_5_bF_buf4_), .B(_259_), .Y(_260_) );
NAND3X1 NAND3X1_178 ( .A(_299_), .B(_258_), .C(_260_), .Y(_261_) );
INVX1 INVX1_119 ( .A(DATA_B[27]), .Y(_262_) );
NAND2X1 NAND2X1_150 ( .A(sel_B_5_bF_buf3_), .B(_262_), .Y(_263_) );
OR2X2 OR2X2_89 ( .A(sel_B_5_bF_buf2_), .B(DATA_B[11]), .Y(_264_) );
NAND3X1 NAND3X1_179 ( .A(sel_B[4]), .B(_264_), .C(_263_), .Y(_265_) );
NAND3X1 NAND3X1_180 ( .A(_298_), .B(_261_), .C(_265_), .Y(_266_) );
OR2X2 OR2X2_90 ( .A(sel_B_5_bF_buf1_), .B(DATA_B[7]), .Y(_267_) );
INVX1 INVX1_120 ( .A(DATA_B[23]), .Y(_268_) );
NAND2X1 NAND2X1_151 ( .A(sel_B_5_bF_buf0_), .B(_268_), .Y(_269_) );
NAND3X1 NAND3X1_181 ( .A(_299_), .B(_267_), .C(_269_), .Y(_270_) );
INVX1 INVX1_121 ( .A(DATA_B[15]), .Y(_271_) );
NAND2X1 NAND2X1_152 ( .A(sel_B_5_bF_buf4_), .B(DATA_B[31]), .Y(_272_) );
OAI21X1 OAI21X1_31 ( .A(_271_), .B(sel_B_5_bF_buf3_), .C(_272_), .Y(_273_) );
NAND2X1 NAND2X1_153 ( .A(sel_B[4]), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_182 ( .A(sel_B[3]), .B(_270_), .C(_274_), .Y(_275_) );
NAND3X1 NAND3X1_183 ( .A(_297_), .B(_266_), .C(_275_), .Y(_276_) );
OR2X2 OR2X2_91 ( .A(sel_A_5_bF_buf0_), .B(DATA_A[3]), .Y(_277_) );
INVX1 INVX1_122 ( .A(DATA_A[19]), .Y(_278_) );
NAND2X1 NAND2X1_154 ( .A(sel_A_5_bF_buf4_), .B(_278_), .Y(_279_) );
NAND3X1 NAND3X1_184 ( .A(_162_), .B(_277_), .C(_279_), .Y(_280_) );
INVX1 INVX1_123 ( .A(DATA_A[27]), .Y(_281_) );
NAND2X1 NAND2X1_155 ( .A(sel_A_5_bF_buf3_), .B(_281_), .Y(_282_) );
OR2X2 OR2X2_92 ( .A(sel_A_5_bF_buf2_), .B(DATA_A[11]), .Y(_283_) );
NAND3X1 NAND3X1_185 ( .A(sel_A[4]), .B(_283_), .C(_282_), .Y(_284_) );
NAND3X1 NAND3X1_186 ( .A(_161_), .B(_280_), .C(_284_), .Y(_285_) );
OR2X2 OR2X2_93 ( .A(sel_A_5_bF_buf1_), .B(DATA_A[7]), .Y(_286_) );
INVX1 INVX1_124 ( .A(DATA_A[23]), .Y(_287_) );
NAND2X1 NAND2X1_156 ( .A(sel_A_5_bF_buf0_), .B(_287_), .Y(_288_) );
NAND3X1 NAND3X1_187 ( .A(_162_), .B(_286_), .C(_288_), .Y(_289_) );
INVX1 INVX1_125 ( .A(DATA_A[15]), .Y(_290_) );
NAND2X1 NAND2X1_157 ( .A(sel_A_5_bF_buf4_), .B(DATA_A[31]), .Y(_291_) );
OAI21X1 OAI21X1_32 ( .A(_290_), .B(sel_A_5_bF_buf3_), .C(_291_), .Y(_292_) );
NAND2X1 NAND2X1_158 ( .A(sel_A[4]), .B(_292_), .Y(_293_) );
NAND3X1 NAND3X1_188 ( .A(sel_A[3]), .B(_289_), .C(_293_), .Y(_294_) );
NAND3X1 NAND3X1_189 ( .A(SEL[1]), .B(_285_), .C(_294_), .Y(_295_) );
AOI21X1 AOI21X1_16 ( .A(_276_), .B(_295_), .C(_296_), .Y(_160__3_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(CLK), .D(_160__0_), .Q(_0__4_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(CLK), .D(_160__1_), .Q(_0__5_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(CLK), .D(_160__2_), .Q(_0__6_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(CLK), .D(_160__3_), .Q(_0__7_) );
INVX2 INVX2_14 ( .A(RESET_L), .Y(_455_) );
INVX2 INVX2_15 ( .A(SEL[2]), .Y(_456_) );
INVX2 INVX2_16 ( .A(sel_B[6]), .Y(_457_) );
INVX4 INVX4_8 ( .A(sel_B[7]), .Y(_458_) );
OR2X2 OR2X2_94 ( .A(DATA_B[0]), .B(sel_B_8_bF_buf2_), .Y(_459_) );
INVX1 INVX1_126 ( .A(DATA_B[16]), .Y(_460_) );
NAND2X1 NAND2X1_159 ( .A(sel_B_8_bF_buf1_), .B(_460_), .Y(_461_) );
NAND3X1 NAND3X1_190 ( .A(_458_), .B(_459_), .C(_461_), .Y(_462_) );
INVX1 INVX1_127 ( .A(DATA_B[24]), .Y(_463_) );
NAND2X1 NAND2X1_160 ( .A(sel_B_8_bF_buf0_), .B(_463_), .Y(_464_) );
OR2X2 OR2X2_95 ( .A(sel_B_8_bF_buf4_), .B(DATA_B[8]), .Y(_465_) );
NAND3X1 NAND3X1_191 ( .A(sel_B[7]), .B(_465_), .C(_464_), .Y(_466_) );
NAND3X1 NAND3X1_192 ( .A(_457_), .B(_462_), .C(_466_), .Y(_467_) );
OR2X2 OR2X2_96 ( .A(sel_B_8_bF_buf3_), .B(DATA_B[4]), .Y(_468_) );
INVX1 INVX1_128 ( .A(DATA_B[20]), .Y(_469_) );
endmodule
