magic
tech scmos
timestamp 1563080643
<< metal1 >>
rect 600 1603 602 1607
rect 606 1603 609 1607
rect 613 1603 616 1607
rect 270 1568 278 1571
rect 1405 1568 1406 1572
rect 1474 1568 1497 1571
rect 270 1566 274 1568
rect 14 1558 25 1561
rect 110 1551 113 1561
rect 158 1552 161 1561
rect 230 1558 241 1561
rect 110 1548 129 1551
rect 350 1551 353 1561
rect 374 1561 377 1568
rect 374 1558 385 1561
rect 470 1558 481 1561
rect 606 1558 614 1561
rect 670 1558 681 1561
rect 734 1558 745 1561
rect 977 1558 982 1562
rect 1038 1558 1049 1561
rect 1158 1561 1161 1568
rect 1150 1558 1161 1561
rect 350 1548 369 1551
rect 598 1548 622 1551
rect 902 1548 921 1551
rect 1094 1551 1097 1558
rect 1070 1548 1089 1551
rect 1094 1548 1105 1551
rect 1162 1548 1169 1551
rect 1214 1548 1222 1551
rect 1294 1548 1302 1551
rect 1358 1548 1377 1551
rect 1390 1548 1401 1551
rect 1470 1551 1473 1558
rect 1462 1548 1473 1551
rect 1582 1548 1590 1551
rect 38 1538 46 1541
rect 70 1538 89 1541
rect 110 1538 118 1541
rect 162 1538 169 1541
rect 282 1538 289 1541
rect 350 1538 358 1541
rect 574 1538 585 1541
rect 618 1538 641 1541
rect 650 1538 657 1541
rect 798 1538 810 1541
rect 918 1538 921 1548
rect 1390 1542 1393 1548
rect 990 1538 998 1541
rect 1006 1538 1025 1541
rect 1110 1538 1134 1541
rect 1178 1538 1193 1541
rect 1206 1538 1214 1541
rect 1550 1538 1566 1541
rect 310 1528 313 1538
rect 806 1536 810 1538
rect 762 1528 769 1531
rect 822 1531 826 1536
rect 822 1528 838 1531
rect 1138 1528 1145 1531
rect 1250 1528 1257 1531
rect 1694 1531 1698 1536
rect 1682 1528 1698 1531
rect 154 1518 155 1522
rect 226 1518 227 1522
rect 389 1518 390 1522
rect 442 1518 443 1522
rect 501 1518 502 1522
rect 666 1518 667 1522
rect 789 1518 790 1522
rect 1034 1518 1035 1522
rect 1205 1518 1206 1522
rect 1112 1503 1114 1507
rect 1118 1503 1121 1507
rect 1125 1503 1128 1507
rect 1014 1488 1025 1491
rect 1022 1482 1025 1488
rect 610 1478 617 1481
rect 70 1462 73 1471
rect 94 1468 105 1471
rect 182 1468 193 1471
rect 342 1468 353 1471
rect 362 1468 369 1471
rect 430 1468 441 1471
rect 534 1471 537 1478
rect 524 1468 537 1471
rect 668 1468 670 1472
rect 754 1468 769 1471
rect 966 1468 982 1471
rect 182 1462 185 1468
rect 502 1461 505 1468
rect 1206 1462 1209 1471
rect 1286 1468 1294 1471
rect 1382 1471 1385 1481
rect 494 1458 505 1461
rect 790 1458 810 1461
rect 842 1458 849 1461
rect 1046 1458 1054 1461
rect 1110 1458 1134 1461
rect 1294 1458 1313 1461
rect 1374 1461 1377 1471
rect 1382 1468 1398 1471
rect 1422 1468 1430 1471
rect 1458 1468 1481 1471
rect 1374 1458 1406 1461
rect 1466 1458 1473 1461
rect 806 1456 810 1458
rect 202 1448 209 1451
rect 542 1448 550 1451
rect 1077 1438 1078 1442
rect 1534 1441 1537 1451
rect 1526 1438 1537 1441
rect 157 1418 158 1422
rect 285 1418 286 1422
rect 333 1418 334 1422
rect 378 1418 379 1422
rect 450 1418 451 1422
rect 1578 1418 1579 1422
rect 600 1403 602 1407
rect 606 1403 609 1407
rect 613 1403 616 1407
rect 1110 1388 1126 1391
rect 1290 1388 1291 1392
rect 1357 1388 1358 1392
rect 1533 1388 1534 1392
rect 1674 1388 1675 1392
rect 1389 1378 1390 1382
rect 118 1368 129 1371
rect 565 1368 566 1372
rect 1586 1368 1598 1371
rect 118 1362 121 1368
rect 410 1358 414 1362
rect 422 1358 441 1361
rect 234 1348 241 1351
rect 494 1351 497 1361
rect 522 1358 529 1361
rect 494 1348 513 1351
rect 886 1348 894 1351
rect 1054 1348 1065 1351
rect 1246 1351 1250 1354
rect 1182 1348 1193 1351
rect 1230 1348 1250 1351
rect 1394 1348 1417 1351
rect 1486 1351 1490 1354
rect 1486 1348 1505 1351
rect 1678 1348 1705 1351
rect 50 1338 65 1341
rect 390 1338 401 1341
rect 462 1338 473 1341
rect 670 1338 678 1341
rect 854 1338 873 1341
rect 902 1338 905 1348
rect 1206 1338 1225 1341
rect 1438 1338 1449 1341
rect 1622 1338 1630 1341
rect 1078 1328 1081 1338
rect 1114 1328 1137 1331
rect 1182 1331 1185 1338
rect 1438 1332 1441 1338
rect 1174 1328 1185 1331
rect 42 1318 43 1322
rect 98 1318 105 1321
rect 226 1318 227 1322
rect 285 1318 286 1322
rect 370 1318 371 1322
rect 533 1318 534 1322
rect 589 1318 590 1322
rect 629 1318 630 1322
rect 685 1318 686 1322
rect 766 1318 774 1321
rect 1112 1303 1114 1307
rect 1118 1303 1121 1307
rect 1125 1303 1128 1307
rect 978 1288 979 1292
rect 1162 1288 1163 1292
rect 1597 1288 1598 1292
rect 238 1278 246 1281
rect 1426 1278 1430 1282
rect 1614 1278 1622 1282
rect 78 1262 81 1271
rect 286 1271 290 1272
rect 294 1271 297 1278
rect 286 1268 297 1271
rect 438 1271 441 1278
rect 1614 1272 1617 1278
rect 430 1268 441 1271
rect 958 1268 969 1271
rect 1214 1268 1225 1271
rect 1274 1268 1289 1271
rect 1430 1268 1438 1271
rect 734 1258 745 1261
rect 1310 1258 1313 1268
rect 1334 1258 1342 1261
rect 1358 1261 1361 1268
rect 1358 1258 1369 1261
rect 1398 1258 1409 1261
rect 1438 1258 1457 1261
rect 1510 1258 1529 1261
rect 1558 1258 1577 1261
rect 390 1251 393 1258
rect 734 1252 737 1258
rect 1398 1252 1401 1258
rect 390 1248 401 1251
rect 702 1248 710 1251
rect 750 1248 761 1251
rect 770 1248 777 1251
rect 958 1248 966 1251
rect 382 1238 390 1241
rect 430 1241 433 1248
rect 422 1238 433 1241
rect 1058 1238 1061 1242
rect 1218 1238 1225 1241
rect 550 1228 553 1238
rect 1349 1218 1350 1222
rect 600 1203 602 1207
rect 606 1203 609 1207
rect 613 1203 616 1207
rect 1458 1188 1459 1192
rect 102 1168 113 1171
rect 270 1168 286 1171
rect 334 1168 342 1171
rect 382 1168 393 1171
rect 883 1168 886 1172
rect 930 1168 933 1172
rect 1526 1168 1537 1171
rect 110 1162 113 1168
rect 390 1162 393 1168
rect 1526 1162 1529 1168
rect 54 1158 65 1161
rect 86 1158 97 1161
rect 138 1158 145 1161
rect 214 1158 225 1161
rect 534 1158 545 1161
rect 610 1148 633 1151
rect 1150 1148 1158 1151
rect 1230 1148 1238 1151
rect 1342 1148 1350 1151
rect 1378 1148 1393 1151
rect 1450 1148 1457 1151
rect 1474 1148 1489 1151
rect 1662 1148 1670 1151
rect 10 1138 17 1141
rect 806 1138 818 1141
rect 1094 1138 1122 1141
rect 1310 1138 1326 1141
rect 1374 1138 1382 1141
rect 1542 1138 1545 1148
rect 1582 1138 1593 1141
rect 74 1128 81 1131
rect 414 1128 422 1131
rect 122 1118 124 1122
rect 229 1118 230 1122
rect 354 1118 361 1121
rect 462 1118 470 1121
rect 662 1118 670 1121
rect 694 1118 702 1121
rect 1112 1103 1114 1107
rect 1118 1103 1121 1107
rect 1125 1103 1128 1107
rect 322 1088 323 1092
rect 150 1071 154 1072
rect 158 1071 161 1078
rect 150 1068 161 1071
rect 418 1068 425 1071
rect 738 1068 745 1071
rect 1054 1068 1062 1071
rect 1350 1068 1358 1071
rect 302 1058 313 1061
rect 574 1058 582 1061
rect 726 1058 734 1061
rect 1086 1058 1094 1061
rect 1270 1061 1274 1064
rect 1262 1058 1274 1061
rect 1318 1058 1329 1061
rect 1358 1058 1377 1061
rect 310 1052 313 1058
rect 10 1048 17 1051
rect 22 1048 30 1051
rect 326 1048 337 1051
rect 446 1048 465 1051
rect 550 1048 558 1051
rect 1406 1048 1417 1051
rect 70 1041 73 1048
rect 62 1038 73 1041
rect 162 1038 177 1041
rect 478 1041 481 1048
rect 470 1038 481 1041
rect 582 1041 585 1048
rect 582 1038 593 1041
rect 502 1028 505 1038
rect 670 1028 673 1038
rect 600 1003 602 1007
rect 606 1003 609 1007
rect 613 1003 616 1007
rect 602 988 617 991
rect 170 968 177 971
rect 414 968 425 971
rect 518 968 529 971
rect 590 968 598 971
rect 914 968 921 971
rect 422 962 425 968
rect 526 962 529 968
rect 38 958 49 961
rect 182 958 201 961
rect 398 958 409 961
rect 502 958 513 961
rect 662 961 665 968
rect 638 958 649 961
rect 654 958 665 961
rect 754 958 761 961
rect 802 958 809 961
rect 790 948 801 951
rect 798 942 801 948
rect 1022 942 1025 951
rect 1630 948 1646 951
rect 62 938 78 941
rect 364 938 377 941
rect 422 938 430 941
rect 530 938 537 941
rect 666 938 673 941
rect 1158 938 1166 941
rect 374 932 377 938
rect 534 928 537 938
rect 670 928 673 938
rect 1026 928 1033 931
rect 1118 928 1134 931
rect 110 918 118 921
rect 742 918 750 921
rect 974 918 982 921
rect 1112 903 1114 907
rect 1118 903 1121 907
rect 1125 903 1128 907
rect 901 888 902 892
rect 1717 888 1718 892
rect 302 878 313 881
rect 310 872 313 878
rect 66 868 73 871
rect 182 868 190 871
rect 578 868 585 871
rect 654 868 662 871
rect 718 871 722 872
rect 726 871 729 878
rect 718 868 729 871
rect 828 868 830 872
rect 842 868 849 871
rect 1134 868 1142 871
rect 342 858 353 861
rect 598 858 614 861
rect 1102 858 1110 861
rect 1578 858 1585 861
rect 38 848 49 851
rect 114 848 121 851
rect 174 851 177 858
rect 342 852 345 858
rect 166 848 177 851
rect 486 851 489 858
rect 1102 857 1106 858
rect 478 848 489 851
rect 802 848 809 851
rect 10 838 17 841
rect 430 838 457 841
rect 490 838 497 841
rect 626 838 633 841
rect 818 838 825 841
rect 1114 818 1129 821
rect 600 803 602 807
rect 606 803 609 807
rect 613 803 616 807
rect 378 788 379 792
rect 950 772 953 781
rect 438 768 449 771
rect 446 762 449 768
rect 110 758 129 761
rect 198 758 209 761
rect 238 758 249 761
rect 270 758 281 761
rect 422 758 433 761
rect 598 758 606 761
rect 1230 758 1238 761
rect 1230 756 1234 758
rect 282 748 289 751
rect 362 748 374 751
rect 146 738 153 741
rect 350 738 369 741
rect 446 738 462 741
rect 778 738 785 741
rect 898 738 905 741
rect 1414 738 1422 741
rect 1442 738 1449 741
rect 150 728 153 738
rect 214 728 217 738
rect 770 728 777 731
rect 1498 728 1505 731
rect 13 718 14 722
rect 194 718 195 722
rect 1112 703 1114 707
rect 1118 703 1121 707
rect 1125 703 1128 707
rect 589 688 590 692
rect 645 688 646 692
rect 757 688 758 692
rect 1102 688 1110 691
rect 214 678 222 682
rect 1718 678 1726 681
rect 214 672 217 678
rect 910 674 914 678
rect 1470 672 1474 677
rect 430 668 441 671
rect 498 668 505 671
rect 598 668 606 671
rect 654 668 662 671
rect 1114 668 1129 671
rect 118 656 122 658
rect 126 641 129 661
rect 890 658 897 661
rect 1286 657 1290 658
rect 258 648 265 651
rect 350 648 361 651
rect 394 648 401 651
rect 478 648 486 651
rect 522 648 526 652
rect 630 648 641 651
rect 678 648 689 651
rect 742 648 753 651
rect 1414 651 1418 654
rect 1414 648 1422 651
rect 246 646 250 648
rect 214 642 218 644
rect 110 638 129 641
rect 194 638 201 641
rect 406 638 414 641
rect 546 638 553 641
rect 310 628 313 638
rect 600 603 602 607
rect 606 603 609 607
rect 613 603 616 607
rect 1718 588 1734 591
rect 1422 572 1425 581
rect 1454 572 1457 581
rect 174 568 190 571
rect 770 558 777 561
rect 1106 558 1113 561
rect 1198 558 1209 561
rect 1270 558 1281 561
rect 1310 558 1321 561
rect 1414 558 1422 561
rect 1494 558 1505 561
rect 1534 558 1542 561
rect 1558 558 1577 561
rect 1610 558 1614 562
rect 1670 558 1681 561
rect 190 552 194 554
rect 934 548 950 551
rect 1602 548 1609 551
rect 14 538 25 541
rect 86 538 105 541
rect 170 538 172 542
rect 1130 538 1137 541
rect 1250 538 1257 541
rect 1386 538 1393 541
rect 1590 538 1601 541
rect 22 532 25 538
rect 220 528 222 532
rect 414 528 417 538
rect 450 528 457 531
rect 1530 518 1531 522
rect 1112 503 1114 507
rect 1118 503 1121 507
rect 1125 503 1128 507
rect 18 488 25 491
rect 122 488 123 492
rect 260 488 262 492
rect 700 488 702 492
rect 1012 488 1014 492
rect 1234 488 1241 491
rect 1426 488 1433 491
rect 470 472 473 481
rect 386 468 393 471
rect 454 468 465 471
rect 526 468 534 471
rect 538 468 545 471
rect 766 471 769 481
rect 1342 478 1350 481
rect 766 468 774 471
rect 898 468 905 471
rect 918 468 929 471
rect 1022 468 1033 471
rect 1094 468 1105 471
rect 1582 471 1585 478
rect 1538 468 1545 471
rect 1572 468 1585 471
rect 454 462 457 468
rect 918 462 921 468
rect 1022 462 1025 468
rect 82 458 97 461
rect 1054 458 1073 461
rect 70 448 89 451
rect 142 448 153 451
rect 326 448 334 451
rect 430 448 438 451
rect 470 451 473 458
rect 470 448 481 451
rect 502 448 513 451
rect 678 448 686 451
rect 790 448 809 451
rect 834 448 841 451
rect 934 451 937 458
rect 934 448 945 451
rect 1070 448 1073 458
rect 1222 448 1230 451
rect 150 442 153 448
rect 442 438 449 441
rect 582 438 606 441
rect 902 441 905 448
rect 902 438 913 441
rect 974 438 1009 441
rect 1085 438 1086 442
rect 1506 438 1513 441
rect 582 428 585 438
rect 974 428 977 438
rect 1510 428 1513 438
rect 600 403 602 407
rect 606 403 609 407
rect 613 403 616 407
rect 174 371 177 381
rect 230 372 233 381
rect 142 368 177 371
rect 1330 368 1337 371
rect 1406 368 1417 371
rect 1438 371 1441 381
rect 1438 368 1462 371
rect 198 361 201 368
rect 198 358 209 361
rect 286 358 294 361
rect 366 358 377 361
rect 510 358 521 361
rect 886 361 889 368
rect 1414 362 1417 368
rect 838 358 849 361
rect 878 358 889 361
rect 1086 358 1094 361
rect 1238 358 1249 361
rect 1686 358 1697 361
rect 1702 358 1710 361
rect 166 352 170 354
rect 762 348 769 351
rect 1042 348 1049 351
rect 1534 351 1538 354
rect 1522 348 1538 351
rect 44 338 46 342
rect 270 338 278 341
rect 342 338 353 341
rect 390 338 393 348
rect 414 338 425 341
rect 476 338 489 341
rect 590 338 598 341
rect 782 338 793 341
rect 822 338 830 341
rect 980 338 982 342
rect 1138 338 1145 341
rect 1326 341 1329 348
rect 1318 338 1329 341
rect 342 332 345 338
rect 382 328 385 338
rect 486 332 489 338
rect 578 328 582 332
rect 1130 328 1137 331
rect 1174 328 1182 331
rect 1278 328 1281 338
rect 1349 318 1350 322
rect 1112 303 1114 307
rect 1118 303 1121 307
rect 1125 303 1128 307
rect 637 288 638 292
rect 661 288 662 292
rect 826 288 833 291
rect 974 288 982 291
rect 1053 288 1054 292
rect 1082 288 1089 291
rect 1173 288 1174 292
rect 1266 288 1267 292
rect 1364 288 1366 292
rect 1386 288 1387 292
rect 1498 288 1499 292
rect 1522 288 1529 291
rect 1554 288 1555 292
rect 1710 288 1718 291
rect 302 268 313 271
rect 382 268 390 271
rect 494 271 497 278
rect 486 268 497 271
rect 950 271 953 278
rect 940 268 953 271
rect 1478 268 1489 271
rect 1486 262 1489 268
rect 606 258 622 261
rect 1118 258 1126 261
rect 1454 258 1473 261
rect 14 248 25 251
rect 422 248 433 251
rect 438 248 446 251
rect 462 248 473 251
rect 618 248 633 251
rect 910 248 921 251
rect 990 248 998 251
rect 1038 248 1049 251
rect 1070 248 1078 251
rect 1158 251 1161 258
rect 1454 256 1458 258
rect 1150 248 1161 251
rect 310 241 313 248
rect 234 238 241 241
rect 310 238 321 241
rect 726 238 742 241
rect 974 238 998 241
rect 1438 238 1446 241
rect 342 228 345 238
rect 542 228 545 238
rect 600 203 602 207
rect 606 203 609 207
rect 613 203 616 207
rect 573 188 574 192
rect 749 188 750 192
rect 1122 188 1129 191
rect 1405 188 1406 192
rect 458 168 459 172
rect 974 168 985 171
rect 1437 168 1438 172
rect 974 162 977 168
rect 118 158 126 161
rect 174 158 182 161
rect 514 158 521 161
rect 990 158 1001 161
rect 1102 158 1110 161
rect 574 148 582 151
rect 642 148 649 151
rect 750 148 758 151
rect 1406 148 1422 151
rect 1538 148 1545 151
rect 1714 148 1734 151
rect 38 138 49 141
rect 366 138 374 141
rect 398 138 406 141
rect 430 138 438 141
rect 582 138 593 141
rect 630 138 641 141
rect 758 138 769 141
rect 966 138 977 141
rect 1378 138 1385 141
rect 1446 138 1457 141
rect 1558 138 1577 141
rect 1670 138 1681 141
rect 46 132 49 138
rect 486 128 489 138
rect 966 132 969 138
rect 1112 103 1114 107
rect 1118 103 1121 107
rect 1125 103 1128 107
rect 18 88 19 92
rect 234 88 235 92
rect 274 88 275 92
rect 362 88 363 92
rect 474 88 475 92
rect 573 88 574 92
rect 693 88 694 92
rect 762 88 763 92
rect 837 88 838 92
rect 877 88 878 92
rect 1042 88 1043 92
rect 1093 88 1094 92
rect 1365 88 1366 92
rect 1389 88 1390 92
rect 1413 88 1414 92
rect 1477 88 1478 92
rect 1501 88 1502 92
rect 606 78 614 81
rect 50 68 57 71
rect 102 68 113 71
rect 214 68 225 71
rect 370 68 377 71
rect 222 62 225 68
rect 422 62 425 71
rect 478 68 489 71
rect 534 68 542 71
rect 606 68 633 71
rect 702 68 710 71
rect 890 68 897 71
rect 962 68 969 71
rect 1174 68 1185 71
rect 1350 68 1358 71
rect 1374 68 1382 71
rect 1518 71 1521 78
rect 1510 68 1521 71
rect 478 62 481 68
rect 70 58 89 61
rect 158 58 166 61
rect 382 58 401 61
rect 942 58 958 61
rect 978 58 985 61
rect 1134 58 1153 61
rect 1214 58 1222 61
rect 1290 58 1297 61
rect 34 48 41 51
rect 70 48 73 58
rect 238 48 249 51
rect 302 48 313 51
rect 366 48 374 51
rect 398 48 401 58
rect 502 48 521 51
rect 646 48 665 51
rect 726 48 737 51
rect 766 48 777 51
rect 822 48 833 51
rect 862 48 873 51
rect 910 48 921 51
rect 1046 48 1057 51
rect 1078 48 1089 51
rect 1150 48 1153 58
rect 1262 48 1273 51
rect 1310 48 1321 51
rect 1438 48 1449 51
rect 413 38 414 42
rect 1382 41 1386 44
rect 1378 38 1386 41
rect 600 3 602 7
rect 606 3 609 7
rect 613 3 616 7
<< m2contact >>
rect 602 1603 606 1607
rect 609 1603 613 1607
rect 278 1568 282 1572
rect 374 1568 378 1572
rect 806 1568 810 1572
rect 1158 1568 1162 1572
rect 1406 1568 1410 1572
rect 1470 1568 1474 1572
rect 1502 1568 1506 1572
rect 1518 1568 1522 1572
rect 62 1558 66 1562
rect 94 1548 98 1552
rect 118 1558 122 1562
rect 206 1558 210 1562
rect 158 1548 162 1552
rect 182 1548 186 1552
rect 334 1548 338 1552
rect 358 1558 362 1562
rect 446 1558 450 1562
rect 494 1558 498 1562
rect 534 1558 538 1562
rect 614 1558 618 1562
rect 630 1558 634 1562
rect 694 1558 698 1562
rect 782 1558 786 1562
rect 902 1558 906 1562
rect 982 1558 986 1562
rect 1078 1558 1082 1562
rect 1094 1558 1098 1562
rect 1174 1558 1178 1562
rect 1302 1558 1306 1562
rect 1366 1558 1370 1562
rect 1454 1558 1458 1562
rect 1470 1558 1474 1562
rect 1478 1558 1482 1562
rect 1534 1558 1538 1562
rect 1558 1558 1562 1562
rect 1590 1558 1594 1562
rect 1614 1558 1618 1562
rect 422 1548 426 1552
rect 542 1548 546 1552
rect 590 1548 594 1552
rect 622 1548 626 1552
rect 758 1548 762 1552
rect 870 1547 874 1551
rect 926 1548 930 1552
rect 942 1548 946 1552
rect 966 1548 970 1552
rect 982 1548 986 1552
rect 998 1548 1002 1552
rect 1158 1548 1162 1552
rect 1182 1548 1186 1552
rect 1222 1548 1226 1552
rect 1246 1548 1250 1552
rect 1302 1548 1306 1552
rect 1318 1548 1322 1552
rect 1382 1548 1386 1552
rect 1430 1548 1434 1552
rect 1446 1548 1450 1552
rect 1486 1548 1490 1552
rect 1526 1548 1530 1552
rect 1574 1548 1578 1552
rect 1590 1548 1594 1552
rect 46 1538 50 1542
rect 118 1538 122 1542
rect 134 1538 138 1542
rect 142 1538 146 1542
rect 158 1538 162 1542
rect 190 1538 194 1542
rect 214 1538 218 1542
rect 254 1538 258 1542
rect 278 1538 282 1542
rect 310 1538 314 1542
rect 326 1538 330 1542
rect 358 1538 362 1542
rect 374 1538 378 1542
rect 398 1538 402 1542
rect 406 1538 410 1542
rect 430 1538 434 1542
rect 454 1538 458 1542
rect 510 1538 514 1542
rect 518 1538 522 1542
rect 558 1538 562 1542
rect 614 1538 618 1542
rect 646 1538 650 1542
rect 710 1538 714 1542
rect 718 1538 722 1542
rect 886 1538 890 1542
rect 910 1538 914 1542
rect 1646 1547 1650 1551
rect 950 1538 954 1542
rect 958 1538 962 1542
rect 998 1538 1002 1542
rect 1062 1538 1066 1542
rect 1094 1538 1098 1542
rect 1134 1538 1138 1542
rect 1158 1538 1162 1542
rect 1174 1538 1178 1542
rect 1214 1538 1218 1542
rect 1238 1538 1242 1542
rect 1310 1538 1314 1542
rect 1326 1538 1330 1542
rect 1350 1538 1354 1542
rect 1390 1538 1394 1542
rect 1438 1538 1442 1542
rect 1470 1538 1474 1542
rect 1518 1538 1522 1542
rect 1542 1538 1546 1542
rect 1566 1538 1570 1542
rect 1598 1538 1602 1542
rect 1654 1538 1658 1542
rect 6 1528 10 1532
rect 78 1528 82 1532
rect 246 1528 250 1532
rect 278 1528 282 1532
rect 302 1528 306 1532
rect 486 1528 490 1532
rect 566 1528 570 1532
rect 686 1528 690 1532
rect 750 1528 754 1532
rect 758 1528 762 1532
rect 774 1528 778 1532
rect 838 1528 842 1532
rect 1014 1528 1018 1532
rect 1046 1528 1050 1532
rect 1118 1528 1122 1532
rect 1134 1528 1138 1532
rect 1230 1528 1234 1532
rect 1246 1528 1250 1532
rect 1286 1528 1290 1532
rect 1334 1528 1338 1532
rect 1342 1528 1346 1532
rect 1414 1528 1418 1532
rect 1422 1528 1426 1532
rect 1678 1528 1682 1532
rect 22 1518 26 1522
rect 62 1518 66 1522
rect 150 1518 154 1522
rect 206 1518 210 1522
rect 222 1518 226 1522
rect 270 1518 274 1522
rect 294 1518 298 1522
rect 318 1518 322 1522
rect 390 1518 394 1522
rect 438 1518 442 1522
rect 470 1518 474 1522
rect 502 1518 506 1522
rect 534 1518 538 1522
rect 662 1518 666 1522
rect 694 1518 698 1522
rect 734 1518 738 1522
rect 790 1518 794 1522
rect 942 1518 946 1522
rect 1030 1518 1034 1522
rect 1206 1518 1210 1522
rect 1614 1518 1618 1522
rect 1114 1503 1118 1507
rect 1121 1503 1125 1507
rect 398 1488 402 1492
rect 990 1488 994 1492
rect 1198 1488 1202 1492
rect 1374 1488 1378 1492
rect 1446 1488 1450 1492
rect 1486 1488 1490 1492
rect 1606 1488 1610 1492
rect 62 1478 66 1482
rect 110 1478 114 1482
rect 182 1478 186 1482
rect 198 1478 202 1482
rect 262 1478 266 1482
rect 310 1478 314 1482
rect 358 1478 362 1482
rect 422 1478 426 1482
rect 470 1478 474 1482
rect 502 1478 506 1482
rect 534 1478 538 1482
rect 550 1478 554 1482
rect 606 1478 610 1482
rect 710 1478 714 1482
rect 750 1478 754 1482
rect 758 1478 762 1482
rect 838 1478 842 1482
rect 910 1478 914 1482
rect 998 1478 1002 1482
rect 1022 1478 1026 1482
rect 1270 1478 1274 1482
rect 54 1468 58 1472
rect 134 1468 138 1472
rect 166 1468 170 1472
rect 238 1468 242 1472
rect 254 1468 258 1472
rect 294 1468 298 1472
rect 358 1468 362 1472
rect 478 1468 482 1472
rect 502 1468 506 1472
rect 622 1468 626 1472
rect 638 1468 642 1472
rect 670 1468 674 1472
rect 734 1468 738 1472
rect 750 1468 754 1472
rect 782 1468 786 1472
rect 854 1468 858 1472
rect 862 1468 866 1472
rect 878 1468 882 1472
rect 894 1468 898 1472
rect 918 1468 922 1472
rect 958 1468 962 1472
rect 982 1468 986 1472
rect 1038 1468 1042 1472
rect 1086 1468 1090 1472
rect 1102 1468 1106 1472
rect 1118 1468 1122 1472
rect 1174 1468 1178 1472
rect 22 1458 26 1462
rect 38 1458 42 1462
rect 70 1458 74 1462
rect 86 1458 90 1462
rect 118 1458 122 1462
rect 158 1458 162 1462
rect 182 1458 186 1462
rect 214 1458 218 1462
rect 286 1458 290 1462
rect 334 1458 338 1462
rect 374 1458 378 1462
rect 414 1458 418 1462
rect 446 1458 450 1462
rect 1230 1468 1234 1472
rect 1254 1468 1258 1472
rect 1294 1468 1298 1472
rect 1326 1468 1330 1472
rect 1510 1478 1514 1482
rect 1598 1478 1602 1482
rect 534 1458 538 1462
rect 582 1458 586 1462
rect 654 1458 658 1462
rect 686 1458 690 1462
rect 726 1458 730 1462
rect 774 1458 778 1462
rect 814 1458 818 1462
rect 838 1458 842 1462
rect 870 1458 874 1462
rect 902 1458 906 1462
rect 942 1458 946 1462
rect 982 1458 986 1462
rect 1022 1458 1026 1462
rect 1054 1458 1058 1462
rect 1078 1458 1082 1462
rect 1134 1458 1138 1462
rect 1158 1458 1162 1462
rect 1182 1458 1186 1462
rect 1206 1458 1210 1462
rect 1222 1458 1226 1462
rect 1246 1458 1250 1462
rect 1318 1458 1322 1462
rect 1366 1458 1370 1462
rect 1398 1468 1402 1472
rect 1430 1468 1434 1472
rect 1438 1468 1442 1472
rect 1454 1468 1458 1472
rect 1494 1468 1498 1472
rect 1566 1468 1570 1472
rect 1654 1468 1658 1472
rect 1406 1458 1410 1462
rect 1430 1458 1434 1462
rect 1462 1458 1466 1462
rect 1502 1458 1506 1462
rect 1526 1458 1530 1462
rect 1542 1458 1546 1462
rect 1574 1458 1578 1462
rect 1614 1458 1618 1462
rect 1654 1458 1658 1462
rect 30 1448 34 1452
rect 70 1448 74 1452
rect 142 1448 146 1452
rect 198 1448 202 1452
rect 270 1448 274 1452
rect 318 1448 322 1452
rect 390 1448 394 1452
rect 462 1448 466 1452
rect 550 1448 554 1452
rect 590 1448 594 1452
rect 646 1448 650 1452
rect 678 1448 682 1452
rect 798 1448 802 1452
rect 950 1448 954 1452
rect 974 1448 978 1452
rect 1030 1448 1034 1452
rect 1062 1448 1066 1452
rect 1094 1448 1098 1452
rect 1166 1448 1170 1452
rect 1198 1448 1202 1452
rect 1206 1448 1210 1452
rect 1238 1448 1242 1452
rect 1270 1448 1274 1452
rect 1302 1448 1306 1452
rect 1422 1448 1426 1452
rect 14 1438 18 1442
rect 222 1438 226 1442
rect 526 1438 530 1442
rect 574 1438 578 1442
rect 662 1438 666 1442
rect 694 1438 698 1442
rect 822 1438 826 1442
rect 934 1438 938 1442
rect 1014 1438 1018 1442
rect 1078 1438 1082 1442
rect 1150 1438 1154 1442
rect 1254 1438 1258 1442
rect 1558 1448 1562 1452
rect 1590 1448 1594 1452
rect 1550 1438 1554 1442
rect 942 1428 946 1432
rect 1158 1428 1162 1432
rect 22 1418 26 1422
rect 158 1418 162 1422
rect 174 1418 178 1422
rect 214 1418 218 1422
rect 286 1418 290 1422
rect 302 1418 306 1422
rect 334 1418 338 1422
rect 374 1418 378 1422
rect 446 1418 450 1422
rect 510 1418 514 1422
rect 558 1418 562 1422
rect 582 1418 586 1422
rect 702 1418 706 1422
rect 718 1418 722 1422
rect 750 1418 754 1422
rect 830 1418 834 1422
rect 894 1418 898 1422
rect 1574 1418 1578 1422
rect 1710 1418 1714 1422
rect 602 1403 606 1407
rect 609 1403 613 1407
rect 910 1388 914 1392
rect 998 1388 1002 1392
rect 1030 1388 1034 1392
rect 1062 1388 1066 1392
rect 1126 1388 1130 1392
rect 1134 1388 1138 1392
rect 1270 1388 1274 1392
rect 1286 1388 1290 1392
rect 1326 1388 1330 1392
rect 1358 1388 1362 1392
rect 1462 1388 1466 1392
rect 1534 1388 1538 1392
rect 1550 1388 1554 1392
rect 1590 1388 1594 1392
rect 1670 1388 1674 1392
rect 22 1378 26 1382
rect 262 1378 266 1382
rect 1390 1378 1394 1382
rect 102 1368 106 1372
rect 566 1368 570 1372
rect 766 1368 770 1372
rect 934 1368 938 1372
rect 966 1368 970 1372
rect 990 1368 994 1372
rect 1022 1368 1026 1372
rect 1262 1368 1266 1372
rect 1470 1368 1474 1372
rect 1582 1368 1586 1372
rect 1598 1368 1602 1372
rect 46 1358 50 1362
rect 86 1358 90 1362
rect 118 1358 122 1362
rect 134 1358 138 1362
rect 142 1358 146 1362
rect 166 1358 170 1362
rect 190 1358 194 1362
rect 230 1358 234 1362
rect 278 1358 282 1362
rect 318 1358 322 1362
rect 374 1358 378 1362
rect 406 1358 410 1362
rect 446 1358 450 1362
rect 6 1348 10 1352
rect 94 1348 98 1352
rect 230 1348 234 1352
rect 406 1348 410 1352
rect 478 1348 482 1352
rect 502 1358 506 1362
rect 518 1358 522 1362
rect 550 1358 554 1362
rect 582 1358 586 1362
rect 622 1358 626 1362
rect 678 1358 682 1362
rect 718 1358 722 1362
rect 782 1358 786 1362
rect 790 1358 794 1362
rect 814 1358 818 1362
rect 894 1358 898 1362
rect 918 1358 922 1362
rect 950 1358 954 1362
rect 1006 1358 1010 1362
rect 1038 1358 1042 1362
rect 1238 1358 1242 1362
rect 1246 1358 1250 1362
rect 1302 1358 1306 1362
rect 1374 1358 1378 1362
rect 1406 1358 1410 1362
rect 1494 1358 1498 1362
rect 1518 1358 1522 1362
rect 1582 1358 1586 1362
rect 1630 1358 1634 1362
rect 1686 1358 1690 1362
rect 1718 1358 1722 1362
rect 566 1348 570 1352
rect 774 1348 778 1352
rect 830 1348 834 1352
rect 862 1348 866 1352
rect 878 1348 882 1352
rect 894 1348 898 1352
rect 902 1348 906 1352
rect 926 1348 930 1352
rect 942 1348 946 1352
rect 958 1348 962 1352
rect 974 1348 978 1352
rect 998 1348 1002 1352
rect 1022 1348 1026 1352
rect 1086 1348 1090 1352
rect 1158 1348 1162 1352
rect 1254 1348 1258 1352
rect 1286 1348 1290 1352
rect 1326 1348 1330 1352
rect 1342 1348 1346 1352
rect 1358 1348 1362 1352
rect 1390 1348 1394 1352
rect 1422 1348 1426 1352
rect 1438 1348 1442 1352
rect 1478 1348 1482 1352
rect 1534 1348 1538 1352
rect 1590 1348 1594 1352
rect 1654 1348 1658 1352
rect 1670 1348 1674 1352
rect 30 1338 34 1342
rect 46 1338 50 1342
rect 78 1338 82 1342
rect 118 1338 122 1342
rect 158 1338 162 1342
rect 182 1338 186 1342
rect 206 1338 210 1342
rect 214 1338 218 1342
rect 294 1338 298 1342
rect 302 1338 306 1342
rect 334 1338 338 1342
rect 358 1338 362 1342
rect 430 1338 434 1342
rect 494 1338 498 1342
rect 518 1338 522 1342
rect 542 1338 546 1342
rect 574 1338 578 1342
rect 598 1338 602 1342
rect 638 1338 642 1342
rect 654 1338 658 1342
rect 678 1338 682 1342
rect 694 1338 698 1342
rect 702 1338 706 1342
rect 734 1338 738 1342
rect 750 1338 754 1342
rect 806 1338 810 1342
rect 838 1338 842 1342
rect 1078 1338 1082 1342
rect 1094 1338 1098 1342
rect 1150 1338 1154 1342
rect 1182 1338 1186 1342
rect 1278 1338 1282 1342
rect 1334 1338 1338 1342
rect 1366 1338 1370 1342
rect 1398 1338 1402 1342
rect 1430 1338 1434 1342
rect 1510 1338 1514 1342
rect 1542 1338 1546 1342
rect 1566 1340 1570 1344
rect 1574 1338 1578 1342
rect 1630 1338 1634 1342
rect 1646 1338 1650 1342
rect 1662 1338 1666 1342
rect 1694 1338 1698 1342
rect 54 1328 58 1332
rect 270 1328 274 1332
rect 326 1328 330 1332
rect 382 1328 386 1332
rect 454 1328 458 1332
rect 646 1328 650 1332
rect 726 1328 730 1332
rect 846 1328 850 1332
rect 1046 1328 1050 1332
rect 1110 1328 1114 1332
rect 1166 1328 1170 1332
rect 1198 1328 1202 1332
rect 1214 1328 1218 1332
rect 1310 1328 1314 1332
rect 1438 1328 1442 1332
rect 1454 1328 1458 1332
rect 1614 1328 1618 1332
rect 1630 1328 1634 1332
rect 38 1318 42 1322
rect 94 1318 98 1322
rect 142 1318 146 1322
rect 166 1318 170 1322
rect 190 1318 194 1322
rect 222 1318 226 1322
rect 254 1318 258 1322
rect 286 1318 290 1322
rect 318 1318 322 1322
rect 350 1318 354 1322
rect 366 1318 370 1322
rect 534 1318 538 1322
rect 590 1318 594 1322
rect 630 1318 634 1322
rect 686 1318 690 1322
rect 718 1318 722 1322
rect 774 1318 778 1322
rect 790 1318 794 1322
rect 814 1318 818 1322
rect 1718 1318 1722 1322
rect 1114 1303 1118 1307
rect 1121 1303 1125 1307
rect 14 1288 18 1292
rect 566 1288 570 1292
rect 814 1288 818 1292
rect 830 1288 834 1292
rect 854 1288 858 1292
rect 974 1288 978 1292
rect 990 1288 994 1292
rect 1030 1288 1034 1292
rect 1038 1288 1042 1292
rect 1158 1288 1162 1292
rect 1246 1288 1250 1292
rect 1294 1288 1298 1292
rect 1478 1288 1482 1292
rect 1542 1288 1546 1292
rect 1598 1288 1602 1292
rect 246 1278 250 1282
rect 294 1278 298 1282
rect 406 1278 410 1282
rect 438 1278 442 1282
rect 502 1278 506 1282
rect 638 1278 642 1282
rect 766 1278 770 1282
rect 950 1278 954 1282
rect 1174 1278 1178 1282
rect 1182 1278 1186 1282
rect 1302 1278 1306 1282
rect 1310 1278 1314 1282
rect 1358 1278 1362 1282
rect 1374 1278 1378 1282
rect 1430 1278 1434 1282
rect 1470 1278 1474 1282
rect 22 1268 26 1272
rect 230 1268 234 1272
rect 254 1268 258 1272
rect 390 1268 394 1272
rect 446 1268 450 1272
rect 510 1268 514 1272
rect 646 1268 650 1272
rect 662 1268 666 1272
rect 734 1268 738 1272
rect 806 1268 810 1272
rect 846 1268 850 1272
rect 1006 1268 1010 1272
rect 1014 1268 1018 1272
rect 1118 1268 1122 1272
rect 1150 1268 1154 1272
rect 1270 1268 1274 1272
rect 1310 1268 1314 1272
rect 1326 1268 1330 1272
rect 1358 1268 1362 1272
rect 1382 1268 1386 1272
rect 1414 1268 1418 1272
rect 1438 1268 1442 1272
rect 1462 1268 1466 1272
rect 1486 1268 1490 1272
rect 1502 1268 1506 1272
rect 1534 1268 1538 1272
rect 1550 1268 1554 1272
rect 1582 1268 1586 1272
rect 1606 1268 1610 1272
rect 1614 1268 1618 1272
rect 1630 1268 1634 1272
rect 1662 1268 1666 1272
rect 46 1258 50 1262
rect 78 1258 82 1262
rect 94 1258 98 1262
rect 126 1258 130 1262
rect 166 1258 170 1262
rect 198 1258 202 1262
rect 214 1258 218 1262
rect 270 1258 274 1262
rect 294 1258 298 1262
rect 326 1258 330 1262
rect 350 1258 354 1262
rect 390 1258 394 1262
rect 462 1258 466 1262
rect 486 1258 490 1262
rect 526 1258 530 1262
rect 550 1258 554 1262
rect 582 1258 586 1262
rect 622 1258 626 1262
rect 678 1258 682 1262
rect 710 1258 714 1262
rect 782 1258 786 1262
rect 886 1258 890 1262
rect 918 1259 922 1263
rect 1102 1259 1106 1263
rect 1190 1258 1194 1262
rect 1206 1258 1210 1262
rect 1238 1258 1242 1262
rect 1262 1258 1266 1262
rect 1278 1258 1282 1262
rect 1342 1258 1346 1262
rect 1494 1258 1498 1262
rect 1670 1258 1674 1262
rect 54 1248 58 1252
rect 86 1248 90 1252
rect 118 1248 122 1252
rect 174 1248 178 1252
rect 206 1248 210 1252
rect 302 1248 306 1252
rect 334 1248 338 1252
rect 342 1248 346 1252
rect 374 1248 378 1252
rect 414 1248 418 1252
rect 430 1248 434 1252
rect 494 1248 498 1252
rect 558 1248 562 1252
rect 630 1248 634 1252
rect 670 1248 674 1252
rect 710 1248 714 1252
rect 734 1248 738 1252
rect 766 1248 770 1252
rect 830 1248 834 1252
rect 966 1248 970 1252
rect 982 1248 986 1252
rect 990 1248 994 1252
rect 1030 1248 1034 1252
rect 1166 1248 1170 1252
rect 1246 1248 1250 1252
rect 1398 1248 1402 1252
rect 1446 1248 1450 1252
rect 1518 1248 1522 1252
rect 1566 1248 1570 1252
rect 1590 1248 1594 1252
rect 1614 1248 1618 1252
rect 38 1238 42 1242
rect 102 1238 106 1242
rect 134 1238 138 1242
rect 158 1238 162 1242
rect 190 1238 194 1242
rect 286 1238 290 1242
rect 318 1238 322 1242
rect 358 1238 362 1242
rect 390 1238 394 1242
rect 478 1238 482 1242
rect 542 1238 546 1242
rect 550 1238 554 1242
rect 614 1238 618 1242
rect 686 1238 690 1242
rect 718 1238 722 1242
rect 790 1238 794 1242
rect 1054 1238 1058 1242
rect 1214 1238 1218 1242
rect 166 1228 170 1232
rect 14 1218 18 1222
rect 46 1218 50 1222
rect 70 1218 74 1222
rect 110 1218 114 1222
rect 142 1218 146 1222
rect 198 1218 202 1222
rect 326 1218 330 1222
rect 350 1218 354 1222
rect 486 1218 490 1222
rect 622 1218 626 1222
rect 678 1218 682 1222
rect 710 1218 714 1222
rect 798 1218 802 1222
rect 1350 1218 1354 1222
rect 1390 1218 1394 1222
rect 1726 1218 1730 1222
rect 602 1203 606 1207
rect 609 1203 613 1207
rect 318 1188 322 1192
rect 718 1188 722 1192
rect 902 1188 906 1192
rect 910 1188 914 1192
rect 1206 1188 1210 1192
rect 1438 1188 1442 1192
rect 1454 1188 1458 1192
rect 1558 1188 1562 1192
rect 526 1178 530 1182
rect 126 1168 130 1172
rect 286 1168 290 1172
rect 294 1168 298 1172
rect 342 1168 346 1172
rect 358 1168 362 1172
rect 462 1168 466 1172
rect 574 1168 578 1172
rect 662 1168 666 1172
rect 694 1168 698 1172
rect 886 1168 890 1172
rect 926 1168 930 1172
rect 110 1158 114 1162
rect 134 1158 138 1162
rect 278 1158 282 1162
rect 342 1158 346 1162
rect 374 1158 378 1162
rect 390 1158 394 1162
rect 478 1158 482 1162
rect 558 1158 562 1162
rect 678 1158 682 1162
rect 710 1158 714 1162
rect 1214 1158 1218 1162
rect 1350 1158 1354 1162
rect 1358 1158 1362 1162
rect 1406 1158 1410 1162
rect 1470 1158 1474 1162
rect 1478 1158 1482 1162
rect 1510 1158 1514 1162
rect 1526 1158 1530 1162
rect 1566 1158 1570 1162
rect 1582 1158 1586 1162
rect 134 1148 138 1152
rect 150 1148 154 1152
rect 182 1148 186 1152
rect 286 1148 290 1152
rect 350 1148 354 1152
rect 398 1148 402 1152
rect 470 1148 474 1152
rect 566 1148 570 1152
rect 606 1148 610 1152
rect 670 1148 674 1152
rect 702 1148 706 1152
rect 782 1147 786 1151
rect 838 1147 842 1151
rect 870 1148 874 1152
rect 974 1147 978 1151
rect 1070 1147 1074 1151
rect 1158 1148 1162 1152
rect 1222 1148 1226 1152
rect 1238 1148 1242 1152
rect 1246 1148 1250 1152
rect 1278 1148 1282 1152
rect 1302 1148 1306 1152
rect 1334 1148 1338 1152
rect 1350 1148 1354 1152
rect 1374 1148 1378 1152
rect 1446 1148 1450 1152
rect 1470 1148 1474 1152
rect 1494 1148 1498 1152
rect 1542 1148 1546 1152
rect 1598 1148 1602 1152
rect 1606 1148 1610 1152
rect 1614 1148 1618 1152
rect 1670 1148 1674 1152
rect 6 1138 10 1142
rect 38 1138 42 1142
rect 110 1138 114 1142
rect 166 1138 170 1142
rect 238 1138 242 1142
rect 254 1138 258 1142
rect 390 1138 394 1142
rect 430 1138 434 1142
rect 446 1138 450 1142
rect 494 1138 498 1142
rect 510 1138 514 1142
rect 518 1138 522 1142
rect 990 1138 994 1142
rect 1238 1138 1242 1142
rect 1270 1138 1274 1142
rect 1326 1138 1330 1142
rect 1382 1138 1386 1142
rect 1406 1138 1410 1142
rect 1414 1138 1418 1142
rect 1422 1140 1426 1144
rect 1446 1138 1450 1142
rect 1502 1138 1506 1142
rect 1526 1138 1530 1142
rect 1550 1138 1554 1142
rect 1574 1138 1578 1142
rect 1622 1138 1626 1142
rect 1662 1138 1666 1142
rect 6 1128 10 1132
rect 70 1128 74 1132
rect 174 1128 178 1132
rect 206 1128 210 1132
rect 246 1128 250 1132
rect 310 1128 314 1132
rect 326 1128 330 1132
rect 422 1128 426 1132
rect 486 1128 490 1132
rect 550 1128 554 1132
rect 1142 1128 1146 1132
rect 1262 1128 1266 1132
rect 1318 1128 1322 1132
rect 1654 1128 1658 1132
rect 30 1118 34 1122
rect 54 1118 58 1122
rect 118 1118 122 1122
rect 198 1118 202 1122
rect 230 1118 234 1122
rect 294 1118 298 1122
rect 350 1118 354 1122
rect 470 1118 474 1122
rect 574 1118 578 1122
rect 590 1118 594 1122
rect 646 1118 650 1122
rect 670 1118 674 1122
rect 702 1118 706 1122
rect 1006 1118 1010 1122
rect 1254 1118 1258 1122
rect 1294 1118 1298 1122
rect 1358 1118 1362 1122
rect 1510 1118 1514 1122
rect 1718 1118 1722 1122
rect 1114 1103 1118 1107
rect 1121 1103 1125 1107
rect 318 1088 322 1092
rect 726 1088 730 1092
rect 1022 1088 1026 1092
rect 1030 1088 1034 1092
rect 1110 1088 1114 1092
rect 1206 1088 1210 1092
rect 1342 1088 1346 1092
rect 1406 1088 1410 1092
rect 1518 1088 1522 1092
rect 1526 1088 1530 1092
rect 6 1078 10 1082
rect 134 1078 138 1082
rect 158 1078 162 1082
rect 198 1078 202 1082
rect 342 1078 346 1082
rect 414 1078 418 1082
rect 454 1078 458 1082
rect 518 1078 522 1082
rect 1310 1078 1314 1082
rect 1414 1078 1418 1082
rect 1422 1078 1426 1082
rect 70 1068 74 1072
rect 126 1068 130 1072
rect 206 1068 210 1072
rect 222 1068 226 1072
rect 270 1068 274 1072
rect 310 1068 314 1072
rect 414 1068 418 1072
rect 478 1068 482 1072
rect 526 1068 530 1072
rect 582 1068 586 1072
rect 718 1068 722 1072
rect 734 1068 738 1072
rect 766 1068 770 1072
rect 1046 1066 1050 1070
rect 1062 1068 1066 1072
rect 1142 1068 1146 1072
rect 1190 1068 1194 1072
rect 1230 1068 1234 1072
rect 1238 1068 1242 1072
rect 1302 1068 1306 1072
rect 1334 1068 1338 1072
rect 1358 1068 1362 1072
rect 1382 1068 1386 1072
rect 1390 1068 1394 1072
rect 1462 1068 1466 1072
rect 1630 1068 1634 1072
rect 1654 1068 1658 1072
rect 30 1058 34 1062
rect 94 1058 98 1062
rect 110 1058 114 1062
rect 158 1058 162 1062
rect 190 1058 194 1062
rect 246 1058 250 1062
rect 286 1058 290 1062
rect 366 1058 370 1062
rect 398 1058 402 1062
rect 438 1058 442 1062
rect 502 1058 506 1062
rect 542 1058 546 1062
rect 558 1058 562 1062
rect 582 1058 586 1062
rect 638 1058 642 1062
rect 670 1058 674 1062
rect 702 1058 706 1062
rect 734 1058 738 1062
rect 790 1058 794 1062
rect 822 1058 826 1062
rect 846 1058 850 1062
rect 878 1058 882 1062
rect 894 1058 898 1062
rect 918 1058 922 1062
rect 966 1058 970 1062
rect 990 1058 994 1062
rect 1070 1058 1074 1062
rect 1094 1058 1098 1062
rect 1166 1058 1170 1062
rect 1222 1058 1226 1062
rect 1246 1058 1250 1062
rect 1278 1058 1282 1062
rect 1294 1058 1298 1062
rect 1454 1059 1458 1063
rect 1558 1058 1562 1062
rect 1590 1059 1594 1063
rect 1646 1059 1650 1063
rect 6 1048 10 1052
rect 30 1048 34 1052
rect 54 1048 58 1052
rect 70 1048 74 1052
rect 102 1048 106 1052
rect 166 1048 170 1052
rect 254 1048 258 1052
rect 278 1048 282 1052
rect 310 1048 314 1052
rect 374 1048 378 1052
rect 406 1048 410 1052
rect 478 1048 482 1052
rect 510 1048 514 1052
rect 558 1048 562 1052
rect 582 1048 586 1052
rect 598 1048 602 1052
rect 646 1048 650 1052
rect 678 1048 682 1052
rect 710 1048 714 1052
rect 758 1048 762 1052
rect 798 1048 802 1052
rect 830 1048 834 1052
rect 838 1048 842 1052
rect 870 1048 874 1052
rect 926 1048 930 1052
rect 1366 1048 1370 1052
rect 38 1038 42 1042
rect 86 1038 90 1042
rect 150 1038 154 1042
rect 158 1038 162 1042
rect 238 1038 242 1042
rect 294 1038 298 1042
rect 358 1038 362 1042
rect 390 1038 394 1042
rect 494 1038 498 1042
rect 502 1038 506 1042
rect 566 1038 570 1042
rect 630 1038 634 1042
rect 662 1038 666 1042
rect 670 1038 674 1042
rect 694 1038 698 1042
rect 782 1038 786 1042
rect 814 1038 818 1042
rect 854 1038 858 1042
rect 886 1038 890 1042
rect 910 1038 914 1042
rect 94 1028 98 1032
rect 638 1028 642 1032
rect 30 1018 34 1022
rect 246 1018 250 1022
rect 262 1018 266 1022
rect 366 1018 370 1022
rect 398 1018 402 1022
rect 702 1018 706 1022
rect 750 1018 754 1022
rect 790 1018 794 1022
rect 822 1018 826 1022
rect 862 1018 866 1022
rect 918 1018 922 1022
rect 1286 1018 1290 1022
rect 1710 1018 1714 1022
rect 602 1003 606 1007
rect 609 1003 613 1007
rect 22 988 26 992
rect 222 988 226 992
rect 478 988 482 992
rect 598 988 602 992
rect 838 988 842 992
rect 878 988 882 992
rect 910 988 914 992
rect 1086 988 1090 992
rect 1262 988 1266 992
rect 1270 988 1274 992
rect 1374 988 1378 992
rect 1390 988 1394 992
rect 1430 988 1434 992
rect 302 978 306 982
rect 718 978 722 982
rect 1686 978 1690 982
rect 54 968 58 972
rect 110 968 114 972
rect 166 968 170 972
rect 214 968 218 972
rect 278 968 282 972
rect 310 968 314 972
rect 366 968 370 972
rect 470 968 474 972
rect 582 968 586 972
rect 598 968 602 972
rect 662 968 666 972
rect 710 968 714 972
rect 742 968 746 972
rect 830 968 834 972
rect 854 968 858 972
rect 886 968 890 972
rect 910 968 914 972
rect 974 968 978 972
rect 126 958 130 962
rect 230 958 234 962
rect 262 958 266 962
rect 294 958 298 962
rect 382 958 386 962
rect 422 958 426 962
rect 486 958 490 962
rect 526 958 530 962
rect 566 958 570 962
rect 726 958 730 962
rect 750 958 754 962
rect 798 958 802 962
rect 814 958 818 962
rect 846 958 850 962
rect 870 958 874 962
rect 902 958 906 962
rect 990 958 994 962
rect 1366 958 1370 962
rect 6 948 10 952
rect 118 948 122 952
rect 222 948 226 952
rect 238 948 242 952
rect 270 948 274 952
rect 286 948 290 952
rect 302 948 306 952
rect 326 948 330 952
rect 374 948 378 952
rect 454 948 458 952
rect 478 948 482 952
rect 558 948 562 952
rect 574 948 578 952
rect 718 948 722 952
rect 750 948 754 952
rect 822 948 826 952
rect 878 948 882 952
rect 918 948 922 952
rect 958 948 962 952
rect 982 948 986 952
rect 998 948 1002 952
rect 1054 948 1058 952
rect 1062 948 1066 952
rect 1094 948 1098 952
rect 1142 948 1146 952
rect 1198 947 1202 951
rect 1302 948 1306 952
rect 1326 948 1330 952
rect 1406 948 1410 952
rect 1462 948 1466 952
rect 1486 948 1490 952
rect 1646 948 1650 952
rect 1710 948 1714 952
rect 78 938 82 942
rect 94 938 98 942
rect 142 938 146 942
rect 158 938 162 942
rect 166 938 170 942
rect 342 938 346 942
rect 430 938 434 942
rect 438 938 442 942
rect 526 938 530 942
rect 542 938 546 942
rect 662 938 666 942
rect 678 938 682 942
rect 694 938 698 942
rect 774 938 778 942
rect 798 938 802 942
rect 862 938 866 942
rect 942 938 946 942
rect 1006 938 1010 942
rect 1022 938 1026 942
rect 1046 938 1050 942
rect 1070 938 1074 942
rect 1102 938 1106 942
rect 1150 938 1154 942
rect 1166 938 1170 942
rect 1182 938 1186 942
rect 1350 938 1354 942
rect 1382 938 1386 942
rect 1510 938 1514 942
rect 1526 938 1530 942
rect 1590 938 1594 942
rect 1606 938 1610 942
rect 1718 938 1722 942
rect 30 928 34 932
rect 70 928 74 932
rect 134 928 138 932
rect 190 928 194 932
rect 254 928 258 932
rect 350 928 354 932
rect 374 928 378 932
rect 390 928 394 932
rect 430 928 434 932
rect 494 928 498 932
rect 622 928 626 932
rect 630 928 634 932
rect 766 928 770 932
rect 798 928 802 932
rect 934 928 938 932
rect 1022 928 1026 932
rect 1086 928 1090 932
rect 1134 928 1138 932
rect 1166 928 1170 932
rect 1398 928 1402 932
rect 1422 928 1426 932
rect 22 918 26 922
rect 118 918 122 922
rect 750 918 754 922
rect 982 918 986 922
rect 1038 918 1042 922
rect 1110 918 1114 922
rect 1694 918 1698 922
rect 1114 903 1118 907
rect 1121 903 1125 907
rect 326 888 330 892
rect 686 888 690 892
rect 862 888 866 892
rect 886 888 890 892
rect 902 888 906 892
rect 1126 888 1130 892
rect 1166 888 1170 892
rect 1198 888 1202 892
rect 1318 888 1322 892
rect 1414 888 1418 892
rect 1430 888 1434 892
rect 1510 888 1514 892
rect 1526 888 1530 892
rect 1646 888 1650 892
rect 1654 888 1658 892
rect 1718 888 1722 892
rect 6 878 10 882
rect 54 878 58 882
rect 62 878 66 882
rect 158 878 162 882
rect 198 878 202 882
rect 374 878 378 882
rect 470 878 474 882
rect 510 878 514 882
rect 574 878 578 882
rect 622 878 626 882
rect 726 878 730 882
rect 838 878 842 882
rect 1422 878 1426 882
rect 22 868 26 872
rect 62 868 66 872
rect 86 868 90 872
rect 174 868 178 872
rect 190 868 194 872
rect 206 868 210 872
rect 246 868 250 872
rect 310 868 314 872
rect 342 868 346 872
rect 366 868 370 872
rect 382 868 386 872
rect 486 868 490 872
rect 518 868 522 872
rect 574 868 578 872
rect 662 868 666 872
rect 702 868 706 872
rect 750 868 754 872
rect 830 868 834 872
rect 838 868 842 872
rect 870 868 874 872
rect 910 868 914 872
rect 1038 868 1042 872
rect 1142 868 1146 872
rect 1182 866 1186 870
rect 1190 868 1194 872
rect 1278 868 1282 872
rect 1294 868 1298 872
rect 1334 868 1338 872
rect 1438 868 1442 872
rect 1454 868 1458 872
rect 1590 868 1594 872
rect 1606 868 1610 872
rect 1622 868 1626 872
rect 1678 868 1682 872
rect 1726 868 1730 872
rect 110 858 114 862
rect 142 858 146 862
rect 174 858 178 862
rect 222 858 226 862
rect 238 858 242 862
rect 270 858 274 862
rect 310 858 314 862
rect 414 858 418 862
rect 446 858 450 862
rect 486 858 490 862
rect 534 858 538 862
rect 558 858 562 862
rect 614 858 618 862
rect 638 858 642 862
rect 726 858 730 862
rect 758 858 762 862
rect 790 858 794 862
rect 814 858 818 862
rect 934 858 938 862
rect 966 858 970 862
rect 998 858 1002 862
rect 1046 858 1050 862
rect 1110 858 1114 862
rect 1158 858 1162 862
rect 1254 858 1258 862
rect 1302 858 1306 862
rect 1350 859 1354 863
rect 1446 858 1450 862
rect 1574 858 1578 862
rect 1630 858 1634 862
rect 1670 858 1674 862
rect 1686 858 1690 862
rect 110 848 114 852
rect 150 848 154 852
rect 190 848 194 852
rect 230 848 234 852
rect 262 848 266 852
rect 318 848 322 852
rect 326 848 330 852
rect 342 848 346 852
rect 398 848 402 852
rect 406 848 410 852
rect 438 848 442 852
rect 502 848 506 852
rect 566 848 570 852
rect 678 848 682 852
rect 686 848 690 852
rect 734 848 738 852
rect 766 848 770 852
rect 798 848 802 852
rect 886 848 890 852
rect 894 848 898 852
rect 942 848 946 852
rect 974 848 978 852
rect 1006 848 1010 852
rect 1710 848 1714 852
rect 6 838 10 842
rect 30 838 34 842
rect 102 838 106 842
rect 134 838 138 842
rect 246 838 250 842
rect 278 838 282 842
rect 302 838 306 842
rect 422 838 426 842
rect 486 838 490 842
rect 550 838 554 842
rect 622 838 626 842
rect 718 838 722 842
rect 750 838 754 842
rect 782 838 786 842
rect 814 838 818 842
rect 926 838 930 842
rect 958 838 962 842
rect 990 838 994 842
rect 1702 838 1706 842
rect 270 828 274 832
rect 670 828 674 832
rect 110 818 114 822
rect 142 818 146 822
rect 390 818 394 822
rect 462 818 466 822
rect 558 818 562 822
rect 790 818 794 822
rect 934 818 938 822
rect 966 818 970 822
rect 998 818 1002 822
rect 1110 818 1114 822
rect 602 803 606 807
rect 609 803 613 807
rect 334 788 338 792
rect 374 788 378 792
rect 398 788 402 792
rect 502 788 506 792
rect 590 788 594 792
rect 638 788 642 792
rect 694 788 698 792
rect 726 788 730 792
rect 814 788 818 792
rect 846 788 850 792
rect 862 788 866 792
rect 870 788 874 792
rect 926 788 930 792
rect 1038 788 1042 792
rect 1262 788 1266 792
rect 1358 788 1362 792
rect 1622 788 1626 792
rect 494 768 498 772
rect 582 768 586 772
rect 630 768 634 772
rect 686 768 690 772
rect 718 768 722 772
rect 822 768 826 772
rect 942 768 946 772
rect 950 768 954 772
rect 6 758 10 762
rect 390 758 394 762
rect 446 758 450 762
rect 510 758 514 762
rect 542 758 546 762
rect 606 758 610 762
rect 646 758 650 762
rect 702 758 706 762
rect 734 758 738 762
rect 806 758 810 762
rect 958 758 962 762
rect 1238 758 1242 762
rect 1462 758 1466 762
rect 62 748 66 752
rect 86 748 90 752
rect 278 748 282 752
rect 358 748 362 752
rect 374 748 378 752
rect 478 748 482 752
rect 502 748 506 752
rect 566 748 570 752
rect 590 748 594 752
rect 638 748 642 752
rect 654 748 658 752
rect 694 748 698 752
rect 726 748 730 752
rect 742 748 746 752
rect 798 748 802 752
rect 814 748 818 752
rect 910 748 914 752
rect 950 748 954 752
rect 966 748 970 752
rect 990 748 994 752
rect 998 748 1002 752
rect 1118 748 1122 752
rect 1166 747 1170 751
rect 1246 748 1250 752
rect 1294 747 1298 751
rect 1366 748 1370 752
rect 1398 748 1402 752
rect 1438 748 1442 752
rect 1470 748 1474 752
rect 1526 748 1530 752
rect 1558 747 1562 751
rect 1590 748 1594 752
rect 1662 748 1666 752
rect 22 738 26 742
rect 46 738 50 742
rect 102 738 106 742
rect 142 738 146 742
rect 158 738 162 742
rect 182 738 186 742
rect 214 738 218 742
rect 222 738 226 742
rect 294 738 298 742
rect 318 738 322 742
rect 406 738 410 742
rect 462 738 466 742
rect 526 738 530 742
rect 758 738 762 742
rect 774 738 778 742
rect 886 740 890 744
rect 894 738 898 742
rect 974 738 978 742
rect 1006 738 1010 742
rect 1094 738 1098 742
rect 1182 738 1186 742
rect 1238 738 1242 742
rect 1278 738 1282 742
rect 1374 738 1378 742
rect 1422 738 1426 742
rect 1438 738 1442 742
rect 1478 738 1482 742
rect 1518 738 1522 742
rect 1638 738 1642 742
rect 54 728 58 732
rect 118 728 122 732
rect 254 728 258 732
rect 262 728 266 732
rect 326 728 330 732
rect 342 728 346 732
rect 358 728 362 732
rect 414 728 418 732
rect 454 728 458 732
rect 518 728 522 732
rect 550 728 554 732
rect 766 728 770 732
rect 838 728 842 732
rect 854 728 858 732
rect 990 728 994 732
rect 1022 728 1026 732
rect 1390 728 1394 732
rect 1430 728 1434 732
rect 1462 728 1466 732
rect 1494 728 1498 732
rect 14 718 18 722
rect 30 718 34 722
rect 78 718 82 722
rect 126 718 130 722
rect 174 718 178 722
rect 190 718 194 722
rect 238 718 242 722
rect 302 718 306 722
rect 670 718 674 722
rect 1014 718 1018 722
rect 1102 718 1106 722
rect 1382 718 1386 722
rect 1486 718 1490 722
rect 1510 718 1514 722
rect 1718 718 1722 722
rect 1114 703 1118 707
rect 1121 703 1125 707
rect 46 688 50 692
rect 390 688 394 692
rect 462 688 466 692
rect 574 688 578 692
rect 590 688 594 692
rect 646 688 650 692
rect 678 688 682 692
rect 702 688 706 692
rect 758 688 762 692
rect 798 688 802 692
rect 830 688 834 692
rect 1110 688 1114 692
rect 1182 688 1186 692
rect 1294 688 1298 692
rect 1446 688 1450 692
rect 1574 688 1578 692
rect 1670 688 1674 692
rect 1694 688 1698 692
rect 54 678 58 682
rect 270 678 274 682
rect 366 678 370 682
rect 422 678 426 682
rect 494 678 498 682
rect 542 678 546 682
rect 622 678 626 682
rect 694 678 698 682
rect 726 678 730 682
rect 734 678 738 682
rect 910 678 914 682
rect 958 678 962 682
rect 1726 678 1730 682
rect 38 668 42 672
rect 62 668 66 672
rect 78 668 82 672
rect 214 668 218 672
rect 230 668 234 672
rect 278 668 282 672
rect 334 668 338 672
rect 374 668 378 672
rect 414 668 418 672
rect 486 668 490 672
rect 494 668 498 672
rect 534 668 538 672
rect 558 668 562 672
rect 606 668 610 672
rect 662 668 666 672
rect 718 668 722 672
rect 766 668 770 672
rect 774 668 778 672
rect 806 668 810 672
rect 942 668 946 672
rect 966 668 970 672
rect 974 668 978 672
rect 982 668 986 672
rect 1022 668 1026 672
rect 1110 668 1114 672
rect 1206 668 1210 672
rect 1318 668 1322 672
rect 1334 668 1338 672
rect 1422 668 1426 672
rect 1470 668 1474 672
rect 1534 668 1538 672
rect 1550 668 1554 672
rect 1590 668 1594 672
rect 1638 668 1642 672
rect 22 658 26 662
rect 94 658 98 662
rect 118 658 122 662
rect 30 648 34 652
rect 86 648 90 652
rect 14 638 18 642
rect 102 638 106 642
rect 166 658 170 662
rect 198 658 202 662
rect 254 658 258 662
rect 294 658 298 662
rect 310 658 314 662
rect 446 658 450 662
rect 526 658 530 662
rect 782 658 786 662
rect 814 658 818 662
rect 862 659 866 663
rect 886 658 890 662
rect 934 658 938 662
rect 990 658 994 662
rect 1006 658 1010 662
rect 1038 659 1042 663
rect 1222 659 1226 663
rect 1286 658 1290 662
rect 1310 658 1314 662
rect 1358 658 1362 662
rect 1430 658 1434 662
rect 1510 658 1514 662
rect 1558 658 1562 662
rect 1606 659 1610 663
rect 1678 658 1682 662
rect 1702 658 1706 662
rect 174 648 178 652
rect 182 648 186 652
rect 246 648 250 652
rect 254 648 258 652
rect 302 648 306 652
rect 342 648 346 652
rect 390 648 394 652
rect 462 648 466 652
rect 470 648 474 652
rect 486 648 490 652
rect 510 648 514 652
rect 526 648 530 652
rect 574 648 578 652
rect 582 648 586 652
rect 958 648 962 652
rect 1422 648 1426 652
rect 134 638 138 642
rect 158 638 162 642
rect 190 638 194 642
rect 214 638 218 642
rect 310 638 314 642
rect 318 638 322 642
rect 414 638 418 642
rect 542 638 546 642
rect 22 618 26 622
rect 46 618 50 622
rect 142 618 146 622
rect 166 618 170 622
rect 190 618 194 622
rect 238 618 242 622
rect 602 603 606 607
rect 609 603 613 607
rect 238 588 242 592
rect 270 588 274 592
rect 446 588 450 592
rect 558 588 562 592
rect 582 588 586 592
rect 702 588 706 592
rect 726 588 730 592
rect 758 588 762 592
rect 798 588 802 592
rect 894 588 898 592
rect 990 588 994 592
rect 998 588 1002 592
rect 1022 588 1026 592
rect 1102 588 1106 592
rect 1166 588 1170 592
rect 1334 588 1338 592
rect 1374 588 1378 592
rect 1654 588 1658 592
rect 1734 588 1738 592
rect 54 578 58 582
rect 78 578 82 582
rect 150 578 154 582
rect 1486 578 1490 582
rect 14 568 18 572
rect 46 568 50 572
rect 142 568 146 572
rect 190 568 194 572
rect 214 568 218 572
rect 246 568 250 572
rect 278 568 282 572
rect 574 568 578 572
rect 718 568 722 572
rect 750 568 754 572
rect 790 568 794 572
rect 1094 568 1098 572
rect 1174 568 1178 572
rect 1366 568 1370 572
rect 1422 568 1426 572
rect 1430 568 1434 572
rect 1454 568 1458 572
rect 1462 568 1466 572
rect 30 558 34 562
rect 62 558 66 562
rect 126 558 130 562
rect 158 558 162 562
rect 198 558 202 562
rect 230 558 234 562
rect 262 558 266 562
rect 350 558 354 562
rect 382 558 386 562
rect 414 558 418 562
rect 590 558 594 562
rect 734 558 738 562
rect 766 558 770 562
rect 1102 558 1106 562
rect 1158 558 1162 562
rect 1350 558 1354 562
rect 1422 558 1426 562
rect 1446 558 1450 562
rect 1542 558 1546 562
rect 1606 558 1610 562
rect 1622 558 1626 562
rect 22 548 26 552
rect 54 548 58 552
rect 110 548 114 552
rect 150 548 154 552
rect 182 548 186 552
rect 190 548 194 552
rect 206 548 210 552
rect 238 548 242 552
rect 270 548 274 552
rect 294 548 298 552
rect 326 548 330 552
rect 358 548 362 552
rect 390 548 394 552
rect 422 548 426 552
rect 494 547 498 551
rect 526 548 530 552
rect 582 548 586 552
rect 638 547 642 551
rect 670 548 674 552
rect 726 548 730 552
rect 758 548 762 552
rect 782 548 786 552
rect 830 547 834 551
rect 862 548 866 552
rect 950 548 954 552
rect 958 548 962 552
rect 1094 548 1098 552
rect 1150 548 1154 552
rect 1166 548 1170 552
rect 1230 548 1234 552
rect 1358 548 1362 552
rect 1406 548 1410 552
rect 1422 548 1426 552
rect 1454 548 1458 552
rect 1598 548 1602 552
rect 1638 548 1642 552
rect 1702 548 1706 552
rect 70 538 74 542
rect 166 538 170 542
rect 310 538 314 542
rect 334 538 338 542
rect 366 538 370 542
rect 398 538 402 542
rect 414 538 418 542
rect 430 538 434 542
rect 462 538 466 542
rect 1006 538 1010 542
rect 1078 538 1082 542
rect 1126 538 1130 542
rect 1222 538 1226 542
rect 1246 538 1250 542
rect 1294 538 1298 542
rect 1342 538 1346 542
rect 1382 538 1386 542
rect 1478 538 1482 542
rect 1518 538 1522 542
rect 1542 538 1546 542
rect 1630 538 1634 542
rect 1694 538 1698 542
rect 22 528 26 532
rect 94 528 98 532
rect 222 528 226 532
rect 318 528 322 532
rect 350 528 354 532
rect 382 528 386 532
rect 446 528 450 532
rect 1190 528 1194 532
rect 1286 528 1290 532
rect 1326 528 1330 532
rect 1382 528 1386 532
rect 1510 528 1514 532
rect 1566 528 1570 532
rect 1582 528 1586 532
rect 1662 528 1666 532
rect 126 518 130 522
rect 1206 518 1210 522
rect 1270 518 1274 522
rect 1310 518 1314 522
rect 1526 518 1530 522
rect 1558 518 1562 522
rect 1678 518 1682 522
rect 1114 503 1118 507
rect 1121 503 1125 507
rect 14 488 18 492
rect 118 488 122 492
rect 166 488 170 492
rect 262 488 266 492
rect 702 488 706 492
rect 1014 488 1018 492
rect 1230 488 1234 492
rect 1422 488 1426 492
rect 1486 488 1490 492
rect 1614 488 1618 492
rect 62 478 66 482
rect 78 478 82 482
rect 134 478 138 482
rect 230 478 234 482
rect 278 478 282 482
rect 382 478 386 482
rect 486 478 490 482
rect 494 478 498 482
rect 534 478 538 482
rect 614 478 618 482
rect 54 468 58 472
rect 102 468 106 472
rect 110 468 114 472
rect 150 468 154 472
rect 222 468 226 472
rect 270 468 274 472
rect 374 468 378 472
rect 382 468 386 472
rect 414 468 418 472
rect 438 468 442 472
rect 470 468 474 472
rect 534 468 538 472
rect 622 468 626 472
rect 638 468 642 472
rect 742 468 746 472
rect 758 468 762 472
rect 782 478 786 482
rect 798 478 802 482
rect 894 478 898 482
rect 934 478 938 482
rect 950 478 954 482
rect 1110 478 1114 482
rect 1214 478 1218 482
rect 1350 478 1354 482
rect 1382 478 1386 482
rect 1534 478 1538 482
rect 1582 478 1586 482
rect 1710 478 1714 482
rect 774 468 778 472
rect 830 468 834 472
rect 886 468 890 472
rect 894 468 898 472
rect 1038 468 1042 472
rect 1046 468 1050 472
rect 1134 468 1138 472
rect 1206 468 1210 472
rect 1334 468 1338 472
rect 1358 468 1362 472
rect 1390 468 1394 472
rect 1406 468 1410 472
rect 1462 468 1466 472
rect 1534 468 1538 472
rect 1598 468 1602 472
rect 1702 468 1706 472
rect 14 458 18 462
rect 38 458 42 462
rect 78 458 82 462
rect 182 458 186 462
rect 206 458 210 462
rect 246 458 250 462
rect 302 458 306 462
rect 342 458 346 462
rect 358 458 362 462
rect 454 458 458 462
rect 470 458 474 462
rect 582 458 586 462
rect 662 458 666 462
rect 686 458 690 462
rect 718 458 722 462
rect 854 458 858 462
rect 870 458 874 462
rect 918 458 922 462
rect 934 458 938 462
rect 974 458 978 462
rect 998 458 1002 462
rect 1022 458 1026 462
rect 1086 458 1090 462
rect 1166 458 1170 462
rect 1190 458 1194 462
rect 1230 458 1234 462
rect 1262 458 1266 462
rect 1294 458 1298 462
rect 1374 458 1378 462
rect 1422 458 1426 462
rect 1478 458 1482 462
rect 1510 458 1514 462
rect 1558 458 1562 462
rect 1582 458 1586 462
rect 1630 458 1634 462
rect 1670 458 1674 462
rect 6 448 10 452
rect 126 448 130 452
rect 166 448 170 452
rect 174 448 178 452
rect 238 448 242 452
rect 286 448 290 452
rect 294 448 298 452
rect 334 448 338 452
rect 406 448 410 452
rect 438 448 442 452
rect 454 448 458 452
rect 558 448 562 452
rect 590 448 594 452
rect 670 448 674 452
rect 686 448 690 452
rect 710 448 714 452
rect 814 448 818 452
rect 830 448 834 452
rect 902 448 906 452
rect 918 448 922 452
rect 982 448 986 452
rect 990 448 994 452
rect 1022 448 1026 452
rect 1062 448 1066 452
rect 1158 448 1162 452
rect 1230 448 1234 452
rect 1254 448 1258 452
rect 1286 448 1290 452
rect 1318 448 1322 452
rect 1414 448 1418 452
rect 1446 448 1450 452
rect 1470 448 1474 452
rect 1502 448 1506 452
rect 1590 448 1594 452
rect 1614 448 1618 452
rect 1622 448 1626 452
rect 1654 448 1658 452
rect 1678 448 1682 452
rect 1686 448 1690 452
rect 22 438 26 442
rect 150 438 154 442
rect 190 438 194 442
rect 254 438 258 442
rect 310 438 314 442
rect 342 438 346 442
rect 438 438 442 442
rect 574 438 578 442
rect 606 438 610 442
rect 654 438 658 442
rect 694 438 698 442
rect 726 438 730 442
rect 854 438 858 442
rect 966 438 970 442
rect 1086 438 1090 442
rect 1174 438 1178 442
rect 1238 438 1242 442
rect 1270 438 1274 442
rect 1302 438 1306 442
rect 1430 438 1434 442
rect 1454 438 1458 442
rect 1486 438 1490 442
rect 1502 438 1506 442
rect 1518 438 1522 442
rect 1574 438 1578 442
rect 1638 438 1642 442
rect 1662 438 1666 442
rect 334 428 338 432
rect 518 428 522 432
rect 846 428 850 432
rect 1262 428 1266 432
rect 182 418 186 422
rect 302 418 306 422
rect 398 418 402 422
rect 422 418 426 422
rect 662 418 666 422
rect 718 418 722 422
rect 822 418 826 422
rect 1142 418 1146 422
rect 1166 418 1170 422
rect 1294 418 1298 422
rect 1630 418 1634 422
rect 602 403 606 407
rect 609 403 613 407
rect 94 388 98 392
rect 118 388 122 392
rect 150 388 154 392
rect 310 388 314 392
rect 526 388 530 392
rect 558 388 562 392
rect 646 388 650 392
rect 678 388 682 392
rect 742 388 746 392
rect 814 388 818 392
rect 894 388 898 392
rect 958 388 962 392
rect 1070 388 1074 392
rect 1094 388 1098 392
rect 1206 388 1210 392
rect 1254 388 1258 392
rect 1286 388 1290 392
rect 1374 388 1378 392
rect 1486 388 1490 392
rect 1566 388 1570 392
rect 1638 388 1642 392
rect 1654 388 1658 392
rect 14 368 18 372
rect 46 368 50 372
rect 86 368 90 372
rect 110 368 114 372
rect 718 378 722 382
rect 854 378 858 382
rect 1238 378 1242 382
rect 182 368 186 372
rect 198 368 202 372
rect 230 368 234 372
rect 238 368 242 372
rect 302 368 306 372
rect 478 368 482 372
rect 550 368 554 372
rect 638 368 642 372
rect 670 368 674 372
rect 710 368 714 372
rect 734 368 738 372
rect 886 368 890 372
rect 950 368 954 372
rect 982 368 986 372
rect 1062 368 1066 372
rect 1102 368 1106 372
rect 1174 368 1178 372
rect 1214 368 1218 372
rect 1262 368 1266 372
rect 1326 368 1330 372
rect 1382 368 1386 372
rect 1430 368 1434 372
rect 1462 368 1466 372
rect 1470 368 1474 372
rect 1478 368 1482 372
rect 1494 368 1498 372
rect 1550 368 1554 372
rect 1558 368 1562 372
rect 1630 368 1634 372
rect 1662 368 1666 372
rect 30 358 34 362
rect 62 358 66 362
rect 70 358 74 362
rect 126 358 130 362
rect 158 358 162 362
rect 214 358 218 362
rect 222 358 226 362
rect 294 358 298 362
rect 390 358 394 362
rect 494 358 498 362
rect 566 358 570 362
rect 574 358 578 362
rect 622 358 626 362
rect 654 358 658 362
rect 686 358 690 362
rect 694 358 698 362
rect 750 358 754 362
rect 758 358 762 362
rect 902 358 906 362
rect 966 358 970 362
rect 998 358 1002 362
rect 1078 358 1082 362
rect 1094 358 1098 362
rect 1190 358 1194 362
rect 1198 358 1202 362
rect 1342 358 1346 362
rect 1366 358 1370 362
rect 1398 358 1402 362
rect 1414 358 1418 362
rect 1446 358 1450 362
rect 1454 358 1458 362
rect 1510 358 1514 362
rect 1614 358 1618 362
rect 1646 358 1650 362
rect 1710 358 1714 362
rect 22 348 26 352
rect 54 348 58 352
rect 78 348 82 352
rect 118 348 122 352
rect 150 348 154 352
rect 166 348 170 352
rect 174 348 178 352
rect 230 348 234 352
rect 254 348 258 352
rect 294 348 298 352
rect 318 348 322 352
rect 390 348 394 352
rect 406 348 410 352
rect 462 348 466 352
rect 486 348 490 352
rect 558 348 562 352
rect 646 348 650 352
rect 678 348 682 352
rect 702 348 706 352
rect 742 348 746 352
rect 758 348 762 352
rect 774 348 778 352
rect 934 348 938 352
rect 958 348 962 352
rect 990 348 994 352
rect 1006 348 1010 352
rect 1038 348 1042 352
rect 1070 348 1074 352
rect 1094 348 1098 352
rect 1182 348 1186 352
rect 1206 348 1210 352
rect 1254 348 1258 352
rect 1326 348 1330 352
rect 1374 348 1378 352
rect 1430 348 1434 352
rect 1462 348 1466 352
rect 1502 348 1506 352
rect 1518 348 1522 352
rect 1542 348 1546 352
rect 1582 348 1586 352
rect 1606 348 1610 352
rect 1622 348 1626 352
rect 1654 348 1658 352
rect 14 338 18 342
rect 46 338 50 342
rect 198 338 202 342
rect 278 338 282 342
rect 334 338 338 342
rect 382 338 386 342
rect 446 338 450 342
rect 534 338 538 342
rect 598 338 602 342
rect 614 338 618 342
rect 830 338 834 342
rect 862 338 866 342
rect 886 338 890 342
rect 918 338 922 342
rect 982 338 986 342
rect 1022 338 1026 342
rect 1134 338 1138 342
rect 1158 338 1162 342
rect 1230 338 1234 342
rect 1278 338 1282 342
rect 1302 338 1306 342
rect 1358 338 1362 342
rect 1414 338 1418 342
rect 1526 338 1530 342
rect 1710 338 1714 342
rect 278 328 282 332
rect 342 328 346 332
rect 358 328 362 332
rect 430 328 434 332
rect 438 328 442 332
rect 486 328 490 332
rect 502 328 506 332
rect 574 328 578 332
rect 798 328 802 332
rect 830 328 834 332
rect 870 328 874 332
rect 910 328 914 332
rect 1030 328 1034 332
rect 1038 328 1042 332
rect 1126 328 1130 332
rect 1182 328 1186 332
rect 1294 328 1298 332
rect 1326 328 1330 332
rect 1678 328 1682 332
rect 814 318 818 322
rect 1350 318 1354 322
rect 1590 318 1594 322
rect 1114 303 1118 307
rect 1121 303 1125 307
rect 22 288 26 292
rect 46 288 50 292
rect 86 288 90 292
rect 150 288 154 292
rect 182 288 186 292
rect 214 288 218 292
rect 470 288 474 292
rect 566 288 570 292
rect 590 288 594 292
rect 638 288 642 292
rect 662 288 666 292
rect 750 288 754 292
rect 766 288 770 292
rect 790 288 794 292
rect 822 288 826 292
rect 982 288 986 292
rect 1014 288 1018 292
rect 1054 288 1058 292
rect 1078 288 1082 292
rect 1174 288 1178 292
rect 1262 288 1266 292
rect 1366 288 1370 292
rect 1382 288 1386 292
rect 1438 288 1442 292
rect 1470 288 1474 292
rect 1494 288 1498 292
rect 1518 288 1522 292
rect 1550 288 1554 292
rect 1678 288 1682 292
rect 1718 288 1722 292
rect 6 278 10 282
rect 70 278 74 282
rect 110 278 114 282
rect 278 278 282 282
rect 302 278 306 282
rect 390 278 394 282
rect 398 278 402 282
rect 406 278 410 282
rect 414 278 418 282
rect 454 278 458 282
rect 494 278 498 282
rect 678 278 682 282
rect 702 278 706 282
rect 846 278 850 282
rect 878 278 882 282
rect 926 278 930 282
rect 950 278 954 282
rect 1030 278 1034 282
rect 1190 278 1194 282
rect 1278 278 1282 282
rect 1398 278 1402 282
rect 1566 278 1570 282
rect 1686 278 1690 282
rect 38 268 42 272
rect 62 268 66 272
rect 270 268 274 272
rect 390 268 394 272
rect 446 268 450 272
rect 502 268 506 272
rect 646 268 650 272
rect 670 268 674 272
rect 710 268 714 272
rect 782 268 786 272
rect 854 268 858 272
rect 894 268 898 272
rect 1062 268 1066 272
rect 1102 268 1106 272
rect 1158 268 1162 272
rect 1182 268 1186 272
rect 1198 268 1202 272
rect 1254 268 1258 272
rect 1286 268 1290 272
rect 1374 268 1378 272
rect 1406 268 1410 272
rect 1542 268 1546 272
rect 1614 268 1618 272
rect 1694 268 1698 272
rect 94 258 98 262
rect 126 258 130 262
rect 142 258 146 262
rect 174 258 178 262
rect 198 258 202 262
rect 238 258 242 262
rect 254 258 258 262
rect 286 258 290 262
rect 342 258 346 262
rect 366 258 370 262
rect 518 258 522 262
rect 542 258 546 262
rect 574 258 578 262
rect 622 258 626 262
rect 694 258 698 262
rect 742 258 746 262
rect 806 258 810 262
rect 822 258 826 262
rect 886 258 890 262
rect 950 258 954 262
rect 982 258 986 262
rect 1006 258 1010 262
rect 1086 258 1090 262
rect 1126 258 1130 262
rect 1158 258 1162 262
rect 1214 258 1218 262
rect 1238 258 1242 262
rect 1302 258 1306 262
rect 1326 258 1330 262
rect 1350 258 1354 262
rect 1422 258 1426 262
rect 1446 258 1450 262
rect 1486 258 1490 262
rect 1518 258 1522 262
rect 1582 258 1586 262
rect 1622 258 1626 262
rect 102 248 106 252
rect 134 248 138 252
rect 166 248 170 252
rect 222 248 226 252
rect 310 248 314 252
rect 326 248 330 252
rect 334 248 338 252
rect 446 248 450 252
rect 550 248 554 252
rect 582 248 586 252
rect 614 248 618 252
rect 654 248 658 252
rect 734 248 738 252
rect 766 248 770 252
rect 814 248 818 252
rect 870 248 874 252
rect 958 248 962 252
rect 998 248 1002 252
rect 1078 248 1082 252
rect 1142 248 1146 252
rect 1166 248 1170 252
rect 1246 248 1250 252
rect 1270 248 1274 252
rect 1334 248 1338 252
rect 1342 248 1346 252
rect 1390 248 1394 252
rect 1502 248 1506 252
rect 1510 248 1514 252
rect 1558 248 1562 252
rect 86 238 90 242
rect 150 238 154 242
rect 182 238 186 242
rect 230 238 234 242
rect 342 238 346 242
rect 350 238 354 242
rect 534 238 538 242
rect 542 238 546 242
rect 566 238 570 242
rect 742 238 746 242
rect 750 238 754 242
rect 830 238 834 242
rect 942 238 946 242
rect 998 238 1002 242
rect 1014 238 1018 242
rect 1086 238 1090 242
rect 1230 238 1234 242
rect 1318 238 1322 242
rect 1358 238 1362 242
rect 1446 238 1450 242
rect 1526 238 1530 242
rect 230 228 234 232
rect 1238 228 1242 232
rect 1326 228 1330 232
rect 902 218 906 222
rect 1470 218 1474 222
rect 602 203 606 207
rect 609 203 613 207
rect 14 188 18 192
rect 110 188 114 192
rect 150 188 154 192
rect 198 188 202 192
rect 238 188 242 192
rect 270 188 274 192
rect 326 188 330 192
rect 494 188 498 192
rect 574 188 578 192
rect 670 188 674 192
rect 750 188 754 192
rect 822 188 826 192
rect 854 188 858 192
rect 918 188 922 192
rect 1014 188 1018 192
rect 1078 188 1082 192
rect 1118 188 1122 192
rect 1222 188 1226 192
rect 1254 188 1258 192
rect 1406 188 1410 192
rect 1470 188 1474 192
rect 1590 188 1594 192
rect 1622 188 1626 192
rect 1310 178 1314 182
rect 38 168 42 172
rect 102 168 106 172
rect 158 168 162 172
rect 190 168 194 172
rect 214 168 218 172
rect 246 168 250 172
rect 278 168 282 172
rect 334 168 338 172
rect 454 168 458 172
rect 502 168 506 172
rect 678 168 682 172
rect 726 168 730 172
rect 830 168 834 172
rect 862 168 866 172
rect 926 168 930 172
rect 1022 168 1026 172
rect 1086 168 1090 172
rect 1134 168 1138 172
rect 1230 168 1234 172
rect 1262 168 1266 172
rect 1438 168 1442 172
rect 1478 168 1482 172
rect 1598 168 1602 172
rect 1630 168 1634 172
rect 54 158 58 162
rect 126 158 130 162
rect 142 158 146 162
rect 182 158 186 162
rect 222 158 226 162
rect 230 158 234 162
rect 262 158 266 162
rect 318 158 322 162
rect 470 158 474 162
rect 510 158 514 162
rect 558 158 562 162
rect 662 158 666 162
rect 694 158 698 162
rect 734 158 738 162
rect 806 158 810 162
rect 814 158 818 162
rect 846 158 850 162
rect 878 158 882 162
rect 910 158 914 162
rect 974 158 978 162
rect 1038 158 1042 162
rect 1110 158 1114 162
rect 1150 158 1154 162
rect 1190 158 1194 162
rect 1246 158 1250 162
rect 1278 158 1282 162
rect 1390 158 1394 162
rect 1422 158 1426 162
rect 1494 158 1498 162
rect 1534 158 1538 162
rect 1582 158 1586 162
rect 1614 158 1618 162
rect 1646 158 1650 162
rect 46 148 50 152
rect 62 148 66 152
rect 110 148 114 152
rect 150 148 154 152
rect 182 148 186 152
rect 238 148 242 152
rect 270 148 274 152
rect 294 148 298 152
rect 326 148 330 152
rect 350 148 354 152
rect 382 148 386 152
rect 414 148 418 152
rect 454 148 458 152
rect 510 148 514 152
rect 526 148 530 152
rect 582 148 586 152
rect 638 148 642 152
rect 654 148 658 152
rect 686 148 690 152
rect 758 148 762 152
rect 822 148 826 152
rect 854 148 858 152
rect 918 148 922 152
rect 942 148 946 152
rect 1030 148 1034 152
rect 1070 148 1074 152
rect 1094 148 1098 152
rect 1142 148 1146 152
rect 1158 148 1162 152
rect 1238 148 1242 152
rect 1270 148 1274 152
rect 1286 148 1290 152
rect 1342 148 1346 152
rect 1422 148 1426 152
rect 1438 148 1442 152
rect 1486 148 1490 152
rect 1502 148 1506 152
rect 1534 148 1538 152
rect 1550 148 1554 152
rect 1590 148 1594 152
rect 1622 148 1626 152
rect 1654 148 1658 152
rect 1662 148 1666 152
rect 1710 148 1714 152
rect 1734 148 1738 152
rect 22 138 26 142
rect 78 138 82 142
rect 134 138 138 142
rect 206 138 210 142
rect 374 138 378 142
rect 406 138 410 142
rect 438 138 442 142
rect 446 138 450 142
rect 478 138 482 142
rect 486 138 490 142
rect 542 138 546 142
rect 710 138 714 142
rect 790 138 794 142
rect 894 138 898 142
rect 958 138 962 142
rect 1054 138 1058 142
rect 1174 138 1178 142
rect 1206 138 1210 142
rect 1326 138 1330 142
rect 1358 138 1362 142
rect 1374 138 1378 142
rect 1414 138 1418 142
rect 1518 138 1522 142
rect 1694 138 1698 142
rect 46 128 50 132
rect 86 128 90 132
rect 310 128 314 132
rect 374 128 378 132
rect 406 128 410 132
rect 438 128 442 132
rect 550 128 554 132
rect 598 128 602 132
rect 622 128 626 132
rect 702 128 706 132
rect 774 128 778 132
rect 782 128 786 132
rect 902 128 906 132
rect 966 128 970 132
rect 1006 128 1010 132
rect 1046 128 1050 132
rect 1182 128 1186 132
rect 1214 128 1218 132
rect 1334 128 1338 132
rect 1366 128 1370 132
rect 1374 128 1378 132
rect 1462 128 1466 132
rect 1526 128 1530 132
rect 1566 128 1570 132
rect 1686 128 1690 132
rect 1302 118 1306 122
rect 1114 103 1118 107
rect 1121 103 1125 107
rect 14 88 18 92
rect 70 88 74 92
rect 150 88 154 92
rect 174 88 178 92
rect 230 88 234 92
rect 270 88 274 92
rect 302 88 306 92
rect 342 88 346 92
rect 358 88 362 92
rect 470 88 474 92
rect 518 88 522 92
rect 558 88 562 92
rect 574 88 578 92
rect 646 88 650 92
rect 670 88 674 92
rect 694 88 698 92
rect 726 88 730 92
rect 758 88 762 92
rect 838 88 842 92
rect 878 88 882 92
rect 910 88 914 92
rect 1006 88 1010 92
rect 1038 88 1042 92
rect 1094 88 1098 92
rect 1150 88 1154 92
rect 1198 88 1202 92
rect 1238 88 1242 92
rect 1262 88 1266 92
rect 1318 88 1322 92
rect 1366 88 1370 92
rect 1390 88 1394 92
rect 1414 88 1418 92
rect 1446 88 1450 92
rect 1478 88 1482 92
rect 1502 88 1506 92
rect 1542 88 1546 92
rect 1574 88 1578 92
rect 1606 88 1610 92
rect 1670 88 1674 92
rect 1718 88 1722 92
rect 118 78 122 82
rect 126 78 130 82
rect 166 78 170 82
rect 254 78 258 82
rect 318 78 322 82
rect 438 78 442 82
rect 454 78 458 82
rect 494 78 498 82
rect 510 78 514 82
rect 614 78 618 82
rect 654 78 658 82
rect 678 78 682 82
rect 742 78 746 82
rect 782 78 786 82
rect 806 78 810 82
rect 814 78 818 82
rect 854 78 858 82
rect 926 78 930 82
rect 958 78 962 82
rect 1062 78 1066 82
rect 1070 78 1074 82
rect 1190 78 1194 82
rect 1278 78 1282 82
rect 1286 78 1290 82
rect 1302 78 1306 82
rect 1342 78 1346 82
rect 1430 78 1434 82
rect 1518 78 1522 82
rect 1550 78 1554 82
rect 1582 78 1586 82
rect 6 68 10 72
rect 30 68 34 72
rect 46 68 50 72
rect 134 68 138 72
rect 190 68 194 72
rect 262 68 266 72
rect 286 68 290 72
rect 326 68 330 72
rect 350 68 354 72
rect 366 68 370 72
rect 430 68 434 72
rect 462 68 466 72
rect 542 68 546 72
rect 582 68 586 72
rect 710 68 714 72
rect 750 68 754 72
rect 846 68 850 72
rect 886 68 890 72
rect 934 68 938 72
rect 958 68 962 72
rect 998 68 1002 72
rect 1022 68 1026 72
rect 1030 68 1034 72
rect 1102 68 1106 72
rect 1126 68 1130 72
rect 1222 68 1226 72
rect 1246 68 1250 72
rect 1334 68 1338 72
rect 1358 68 1362 72
rect 1382 68 1386 72
rect 1398 68 1402 72
rect 1422 68 1426 72
rect 1462 68 1466 72
rect 1486 68 1490 72
rect 1526 68 1530 72
rect 1558 68 1562 72
rect 1590 68 1594 72
rect 1662 68 1666 72
rect 1694 68 1698 72
rect 1702 66 1706 70
rect 94 58 98 62
rect 166 58 170 62
rect 198 58 202 62
rect 222 58 226 62
rect 414 58 418 62
rect 422 58 426 62
rect 478 58 482 62
rect 590 58 594 62
rect 790 58 794 62
rect 958 58 962 62
rect 974 58 978 62
rect 990 58 994 62
rect 1166 58 1170 62
rect 1222 58 1226 62
rect 1286 58 1290 62
rect 1686 58 1690 62
rect 22 48 26 52
rect 30 48 34 52
rect 46 48 50 52
rect 78 48 82 52
rect 174 48 178 52
rect 278 48 282 52
rect 342 48 346 52
rect 374 48 378 52
rect 390 48 394 52
rect 478 48 482 52
rect 558 48 562 52
rect 566 48 570 52
rect 686 48 690 52
rect 950 48 954 52
rect 974 48 978 52
rect 1006 48 1010 52
rect 1142 48 1146 52
rect 1238 48 1242 52
rect 1358 48 1362 52
rect 1406 48 1410 52
rect 1470 48 1474 52
rect 1494 48 1498 52
rect 414 38 418 42
rect 1374 38 1378 42
rect 446 18 450 22
rect 602 3 606 7
rect 609 3 613 7
<< metal2 >>
rect 62 1638 66 1642
rect 198 1638 202 1642
rect 294 1638 298 1642
rect 414 1638 418 1642
rect 446 1638 450 1642
rect 550 1641 554 1642
rect 542 1638 554 1641
rect 566 1638 570 1642
rect 630 1638 634 1642
rect 646 1638 650 1642
rect 670 1638 674 1642
rect 694 1638 698 1642
rect 710 1638 714 1642
rect 726 1638 730 1642
rect 750 1638 754 1642
rect 766 1638 770 1642
rect 1230 1638 1234 1642
rect 62 1592 65 1638
rect 62 1562 65 1588
rect 118 1562 121 1588
rect 158 1552 161 1558
rect 186 1548 190 1551
rect 198 1551 201 1638
rect 294 1631 297 1638
rect 294 1628 305 1631
rect 278 1572 281 1608
rect 206 1562 209 1568
rect 194 1548 201 1551
rect 94 1542 97 1548
rect 130 1538 134 1541
rect 162 1538 166 1541
rect 186 1538 190 1541
rect 218 1538 222 1541
rect 6 1522 9 1528
rect 6 1462 9 1518
rect 22 1471 25 1518
rect 14 1468 25 1471
rect 6 1352 9 1448
rect 14 1442 17 1468
rect 38 1462 41 1468
rect 46 1462 49 1538
rect 82 1528 86 1531
rect 62 1492 65 1518
rect 110 1482 113 1528
rect 118 1482 121 1538
rect 54 1472 57 1478
rect 26 1458 30 1461
rect 22 1402 25 1418
rect 30 1412 33 1448
rect 54 1432 57 1468
rect 62 1462 65 1478
rect 70 1462 73 1468
rect 134 1462 137 1468
rect 142 1462 145 1538
rect 246 1532 249 1568
rect 258 1538 265 1541
rect 282 1538 286 1541
rect 82 1458 86 1461
rect 22 1382 25 1388
rect 6 1261 9 1348
rect 22 1338 30 1341
rect 22 1322 25 1338
rect 38 1331 41 1398
rect 62 1381 65 1458
rect 118 1452 121 1458
rect 150 1451 153 1518
rect 182 1482 185 1518
rect 198 1482 201 1488
rect 170 1468 174 1471
rect 158 1462 161 1468
rect 182 1462 185 1468
rect 146 1448 153 1451
rect 70 1442 73 1448
rect 58 1378 65 1381
rect 46 1362 49 1368
rect 54 1352 57 1378
rect 86 1362 89 1408
rect 106 1368 110 1371
rect 118 1362 121 1368
rect 46 1342 49 1348
rect 54 1332 57 1348
rect 78 1332 81 1338
rect 38 1328 49 1331
rect 14 1292 17 1298
rect 22 1272 25 1318
rect 6 1258 14 1261
rect 6 1232 9 1248
rect 14 1212 17 1218
rect 22 1202 25 1268
rect 38 1242 41 1318
rect 46 1262 49 1328
rect 86 1302 89 1358
rect 94 1342 97 1348
rect 118 1342 121 1348
rect 78 1262 81 1268
rect 94 1262 97 1318
rect 6 1142 9 1148
rect 38 1132 41 1138
rect 10 1128 14 1131
rect 6 1082 9 1098
rect 14 1062 17 1088
rect 10 1048 14 1051
rect 22 992 25 1128
rect 30 1062 33 1118
rect 30 1032 33 1048
rect 38 1042 41 1058
rect 6 952 9 978
rect 30 941 33 1018
rect 30 938 41 941
rect 30 922 33 928
rect 6 882 9 898
rect 22 882 25 918
rect 22 872 25 878
rect 6 762 9 838
rect 22 742 25 868
rect 38 862 41 938
rect 30 842 33 848
rect 22 732 25 738
rect 6 632 9 648
rect 14 642 17 718
rect 30 661 33 718
rect 26 658 33 661
rect 38 672 41 798
rect 46 772 49 1218
rect 54 1192 57 1248
rect 70 1162 73 1218
rect 70 1132 73 1138
rect 54 1062 57 1118
rect 78 1102 81 1258
rect 86 1242 89 1248
rect 102 1242 105 1278
rect 126 1262 129 1368
rect 134 1362 137 1378
rect 158 1362 161 1418
rect 146 1358 150 1361
rect 174 1361 177 1418
rect 170 1358 177 1361
rect 190 1362 193 1478
rect 206 1452 209 1518
rect 214 1462 217 1468
rect 198 1412 201 1448
rect 222 1442 225 1518
rect 246 1482 249 1528
rect 262 1482 265 1538
rect 302 1532 305 1628
rect 358 1562 361 1588
rect 374 1562 377 1568
rect 362 1558 366 1561
rect 322 1538 326 1541
rect 310 1532 313 1538
rect 334 1532 337 1548
rect 398 1542 401 1548
rect 354 1538 358 1541
rect 378 1538 382 1541
rect 282 1528 286 1531
rect 242 1468 246 1471
rect 254 1442 257 1468
rect 262 1462 265 1478
rect 270 1452 273 1518
rect 294 1472 297 1518
rect 302 1512 305 1528
rect 306 1478 310 1481
rect 318 1472 321 1518
rect 358 1482 361 1488
rect 354 1468 358 1471
rect 282 1458 286 1461
rect 378 1458 382 1461
rect 314 1448 318 1451
rect 214 1372 217 1418
rect 230 1362 233 1388
rect 182 1342 185 1348
rect 158 1322 161 1338
rect 206 1332 209 1338
rect 114 1248 118 1251
rect 142 1241 145 1318
rect 166 1271 169 1318
rect 138 1238 145 1241
rect 158 1268 169 1271
rect 158 1242 161 1268
rect 170 1258 174 1261
rect 166 1232 169 1238
rect 174 1222 177 1248
rect 110 1182 113 1218
rect 122 1168 126 1171
rect 110 1162 113 1168
rect 134 1162 137 1218
rect 142 1162 145 1218
rect 130 1158 134 1161
rect 182 1152 185 1308
rect 190 1242 193 1318
rect 206 1272 209 1328
rect 214 1322 217 1338
rect 222 1282 225 1318
rect 230 1312 233 1348
rect 254 1331 257 1438
rect 334 1432 337 1458
rect 390 1452 393 1518
rect 398 1492 401 1538
rect 406 1532 409 1538
rect 398 1462 401 1488
rect 414 1462 417 1638
rect 446 1612 449 1638
rect 446 1562 449 1608
rect 534 1562 537 1578
rect 542 1562 545 1638
rect 422 1552 425 1558
rect 494 1542 497 1558
rect 542 1552 545 1558
rect 518 1542 521 1548
rect 426 1538 430 1541
rect 450 1538 454 1541
rect 422 1482 425 1508
rect 418 1458 425 1461
rect 286 1392 289 1418
rect 262 1372 265 1378
rect 282 1358 286 1361
rect 294 1352 297 1428
rect 302 1362 305 1418
rect 334 1362 337 1418
rect 374 1402 377 1418
rect 322 1358 326 1361
rect 378 1358 382 1361
rect 398 1352 401 1458
rect 406 1362 409 1368
rect 294 1342 297 1348
rect 330 1338 334 1341
rect 302 1332 305 1338
rect 358 1332 361 1338
rect 254 1328 265 1331
rect 230 1272 233 1288
rect 254 1281 257 1318
rect 250 1278 257 1281
rect 214 1262 217 1268
rect 198 1242 201 1258
rect 210 1248 214 1251
rect 206 1232 209 1248
rect 198 1192 201 1218
rect 138 1148 150 1151
rect 166 1142 169 1148
rect 110 1122 113 1138
rect 174 1122 177 1128
rect 54 1042 57 1048
rect 62 1022 65 1098
rect 74 1068 81 1071
rect 70 1042 73 1048
rect 54 962 57 968
rect 62 951 65 1018
rect 54 948 65 951
rect 78 952 81 1068
rect 94 1062 97 1068
rect 102 1052 105 1098
rect 110 1062 113 1068
rect 118 1062 121 1118
rect 134 1082 137 1118
rect 158 1072 161 1078
rect 86 1042 89 1048
rect 94 1032 97 1038
rect 126 1002 129 1068
rect 154 1058 158 1061
rect 166 1042 169 1048
rect 146 1038 150 1041
rect 106 968 110 971
rect 130 958 134 961
rect 158 952 161 1038
rect 182 1031 185 1148
rect 210 1128 214 1131
rect 198 1082 201 1118
rect 206 1092 209 1128
rect 238 1122 241 1138
rect 246 1132 249 1278
rect 262 1271 265 1328
rect 386 1328 390 1331
rect 270 1282 273 1328
rect 258 1268 265 1271
rect 270 1262 273 1268
rect 222 1072 225 1078
rect 210 1068 214 1071
rect 190 1032 193 1058
rect 182 1028 190 1031
rect 222 992 225 1058
rect 230 1041 233 1118
rect 254 1112 257 1138
rect 246 1062 249 1068
rect 262 1051 265 1218
rect 278 1162 281 1328
rect 326 1322 329 1328
rect 406 1322 409 1348
rect 286 1272 289 1318
rect 294 1272 297 1278
rect 290 1258 294 1261
rect 290 1238 294 1241
rect 302 1222 305 1248
rect 318 1242 321 1318
rect 326 1262 329 1268
rect 350 1262 353 1318
rect 318 1192 321 1208
rect 298 1168 302 1171
rect 270 1072 273 1108
rect 278 1092 281 1158
rect 286 1152 289 1168
rect 310 1132 313 1138
rect 282 1058 286 1061
rect 258 1048 265 1051
rect 230 1038 238 1041
rect 170 968 174 971
rect 210 968 214 971
rect 230 962 233 968
rect 238 952 241 1028
rect 246 952 249 1018
rect 254 962 257 1048
rect 278 1042 281 1048
rect 294 1042 297 1118
rect 310 1072 313 1118
rect 318 1092 321 1168
rect 326 1152 329 1218
rect 334 1192 337 1248
rect 342 1222 345 1248
rect 358 1232 361 1238
rect 338 1168 342 1171
rect 326 1132 329 1138
rect 342 1112 345 1158
rect 350 1152 353 1218
rect 366 1171 369 1318
rect 390 1272 393 1318
rect 406 1282 409 1308
rect 402 1278 406 1281
rect 390 1252 393 1258
rect 378 1248 382 1251
rect 386 1238 390 1241
rect 414 1212 417 1248
rect 422 1222 425 1458
rect 438 1452 441 1518
rect 446 1482 449 1538
rect 510 1532 513 1538
rect 466 1518 470 1521
rect 446 1462 449 1478
rect 446 1422 449 1428
rect 446 1362 449 1368
rect 430 1322 433 1338
rect 438 1282 441 1348
rect 454 1332 457 1508
rect 486 1492 489 1528
rect 530 1518 534 1521
rect 502 1512 505 1518
rect 502 1482 505 1488
rect 466 1478 470 1481
rect 462 1452 465 1458
rect 478 1392 481 1468
rect 502 1462 505 1468
rect 518 1441 521 1518
rect 534 1472 537 1478
rect 530 1458 534 1461
rect 518 1438 526 1441
rect 510 1401 513 1418
rect 510 1398 521 1401
rect 502 1362 505 1368
rect 474 1348 478 1351
rect 494 1342 497 1358
rect 502 1282 505 1348
rect 510 1292 513 1388
rect 518 1362 521 1398
rect 542 1352 545 1548
rect 558 1542 561 1548
rect 566 1532 569 1638
rect 630 1612 633 1638
rect 600 1603 602 1607
rect 606 1603 609 1607
rect 613 1603 616 1607
rect 646 1582 649 1638
rect 670 1582 673 1638
rect 694 1612 697 1638
rect 710 1592 713 1638
rect 630 1562 633 1578
rect 586 1548 590 1551
rect 566 1502 569 1528
rect 550 1482 553 1498
rect 554 1448 558 1451
rect 574 1442 577 1508
rect 606 1482 609 1548
rect 614 1542 617 1558
rect 622 1552 625 1558
rect 646 1542 649 1548
rect 642 1468 646 1471
rect 582 1462 585 1468
rect 590 1452 593 1458
rect 622 1442 625 1468
rect 654 1462 657 1468
rect 646 1442 649 1448
rect 662 1442 665 1518
rect 670 1472 673 1478
rect 678 1462 681 1588
rect 726 1572 729 1638
rect 686 1532 689 1568
rect 698 1558 702 1561
rect 718 1542 721 1548
rect 750 1542 753 1638
rect 758 1552 761 1558
rect 706 1538 710 1541
rect 686 1482 689 1528
rect 686 1462 689 1468
rect 678 1452 681 1458
rect 682 1448 686 1451
rect 694 1442 697 1518
rect 706 1478 710 1481
rect 718 1431 721 1538
rect 766 1532 769 1638
rect 1230 1612 1233 1638
rect 1402 1568 1406 1571
rect 1462 1568 1470 1571
rect 1506 1568 1510 1571
rect 786 1558 790 1561
rect 806 1552 809 1568
rect 902 1562 905 1568
rect 1158 1562 1161 1568
rect 978 1558 982 1561
rect 1074 1558 1078 1561
rect 1170 1558 1174 1561
rect 1298 1558 1302 1561
rect 998 1552 1001 1558
rect 774 1532 777 1548
rect 930 1548 934 1551
rect 746 1528 750 1531
rect 734 1492 737 1518
rect 758 1491 761 1528
rect 750 1488 761 1491
rect 750 1482 753 1488
rect 726 1462 729 1478
rect 758 1472 761 1478
rect 738 1468 742 1471
rect 750 1462 753 1468
rect 718 1428 729 1431
rect 550 1362 553 1368
rect 558 1352 561 1418
rect 566 1372 569 1378
rect 574 1361 577 1398
rect 582 1382 585 1418
rect 600 1403 602 1407
rect 606 1403 609 1407
rect 613 1403 616 1407
rect 678 1362 681 1368
rect 574 1358 582 1361
rect 618 1358 622 1361
rect 702 1352 705 1418
rect 718 1362 721 1418
rect 566 1342 569 1348
rect 574 1342 577 1348
rect 654 1342 657 1348
rect 522 1338 526 1341
rect 546 1338 550 1341
rect 602 1338 606 1341
rect 642 1338 646 1341
rect 566 1332 569 1338
rect 642 1328 646 1331
rect 510 1272 513 1288
rect 430 1242 433 1248
rect 362 1168 369 1171
rect 374 1162 377 1168
rect 390 1162 393 1168
rect 446 1162 449 1268
rect 462 1262 465 1268
rect 526 1262 529 1268
rect 482 1258 486 1261
rect 498 1248 502 1251
rect 474 1238 478 1241
rect 534 1241 537 1318
rect 566 1292 569 1328
rect 546 1258 550 1261
rect 562 1248 566 1251
rect 534 1238 542 1241
rect 550 1232 553 1238
rect 582 1222 585 1258
rect 590 1242 593 1318
rect 630 1262 633 1318
rect 638 1282 641 1328
rect 646 1272 649 1278
rect 662 1272 665 1278
rect 678 1262 681 1338
rect 686 1282 689 1318
rect 610 1238 614 1241
rect 622 1232 625 1258
rect 486 1172 489 1218
rect 600 1203 602 1207
rect 606 1203 609 1207
rect 613 1203 616 1207
rect 526 1182 529 1188
rect 458 1168 462 1171
rect 558 1162 561 1188
rect 574 1172 577 1178
rect 482 1158 486 1161
rect 402 1148 406 1151
rect 338 1078 342 1081
rect 310 1052 313 1058
rect 262 1022 265 1038
rect 262 962 265 1018
rect 282 968 286 971
rect 294 962 297 978
rect 302 972 305 978
rect 350 972 353 1118
rect 362 1058 366 1061
rect 358 1042 361 1048
rect 366 992 369 1018
rect 314 968 321 971
rect 362 968 366 971
rect 162 948 169 951
rect 54 882 57 948
rect 78 942 81 948
rect 118 942 121 948
rect 94 932 97 938
rect 134 932 137 948
rect 166 942 169 948
rect 62 882 65 888
rect 58 868 62 871
rect 70 812 73 928
rect 118 892 121 918
rect 142 912 145 938
rect 158 932 161 938
rect 174 882 177 948
rect 222 942 225 948
rect 254 932 257 938
rect 190 922 193 928
rect 190 902 193 918
rect 154 878 158 881
rect 194 878 198 881
rect 86 872 89 878
rect 110 862 113 868
rect 110 842 113 848
rect 98 838 102 841
rect 118 832 121 878
rect 138 858 142 861
rect 106 818 110 821
rect 70 802 73 808
rect 46 742 49 758
rect 58 748 62 751
rect 82 748 86 751
rect 102 732 105 738
rect 110 732 113 778
rect 118 732 121 828
rect 134 822 137 838
rect 142 752 145 818
rect 138 738 142 741
rect 50 728 54 731
rect 46 692 49 718
rect 54 682 57 708
rect 62 672 65 698
rect 78 682 81 718
rect 102 712 105 728
rect 150 722 153 848
rect 158 842 161 878
rect 174 872 177 878
rect 194 868 198 871
rect 174 852 177 858
rect 186 848 190 851
rect 206 822 209 868
rect 222 862 225 868
rect 230 852 233 878
rect 238 862 241 888
rect 262 882 265 958
rect 270 952 273 958
rect 306 948 310 951
rect 286 942 289 948
rect 318 941 321 968
rect 374 961 377 1048
rect 382 1041 385 1148
rect 430 1142 433 1158
rect 470 1142 473 1148
rect 498 1138 502 1141
rect 390 1122 393 1138
rect 446 1132 449 1138
rect 510 1132 513 1138
rect 518 1132 521 1138
rect 414 1082 417 1118
rect 394 1058 398 1061
rect 402 1048 406 1051
rect 382 1038 390 1041
rect 398 1012 401 1018
rect 414 1002 417 1068
rect 414 982 417 998
rect 422 981 425 1128
rect 486 1122 489 1128
rect 518 1122 521 1128
rect 550 1122 553 1128
rect 478 1118 486 1121
rect 470 1102 473 1118
rect 438 1062 441 1068
rect 454 1022 457 1078
rect 478 1072 481 1118
rect 498 1058 502 1061
rect 510 1052 513 1088
rect 518 1082 521 1118
rect 558 1092 561 1158
rect 610 1148 614 1151
rect 566 1142 569 1148
rect 590 1122 593 1128
rect 574 1072 577 1118
rect 590 1071 593 1118
rect 622 1082 625 1218
rect 630 1162 633 1248
rect 662 1172 665 1258
rect 674 1248 678 1251
rect 686 1242 689 1258
rect 694 1251 697 1338
rect 702 1332 705 1338
rect 726 1332 729 1428
rect 750 1362 753 1418
rect 734 1342 737 1358
rect 750 1332 753 1338
rect 702 1282 705 1328
rect 710 1262 713 1268
rect 694 1248 705 1251
rect 678 1171 681 1218
rect 702 1182 705 1248
rect 710 1242 713 1248
rect 718 1242 721 1318
rect 734 1272 737 1278
rect 758 1271 761 1448
rect 766 1372 769 1488
rect 774 1462 777 1488
rect 790 1482 793 1518
rect 786 1468 790 1471
rect 798 1452 801 1488
rect 782 1362 785 1438
rect 790 1362 793 1418
rect 774 1342 777 1348
rect 766 1282 769 1308
rect 758 1268 769 1271
rect 734 1252 737 1258
rect 766 1252 769 1268
rect 774 1261 777 1318
rect 782 1312 785 1358
rect 806 1342 809 1538
rect 838 1482 841 1528
rect 814 1431 817 1458
rect 822 1442 825 1478
rect 854 1472 857 1538
rect 870 1532 873 1547
rect 942 1542 945 1548
rect 966 1542 969 1548
rect 862 1472 865 1478
rect 842 1458 846 1461
rect 814 1428 825 1431
rect 814 1362 817 1368
rect 822 1341 825 1428
rect 830 1352 833 1418
rect 854 1362 857 1468
rect 870 1462 873 1508
rect 878 1472 881 1498
rect 866 1458 870 1461
rect 886 1412 889 1538
rect 910 1532 913 1538
rect 910 1502 913 1528
rect 938 1518 942 1521
rect 910 1482 913 1488
rect 950 1482 953 1538
rect 958 1512 961 1538
rect 982 1522 985 1548
rect 998 1532 1001 1538
rect 1006 1522 1009 1558
rect 1094 1552 1097 1558
rect 1162 1548 1166 1551
rect 1174 1542 1177 1558
rect 1242 1548 1246 1551
rect 1298 1548 1302 1551
rect 1314 1548 1318 1551
rect 1182 1542 1185 1548
rect 1138 1538 1142 1541
rect 1154 1538 1158 1541
rect 990 1492 993 1508
rect 894 1472 897 1478
rect 958 1472 961 1478
rect 922 1468 926 1471
rect 894 1452 897 1468
rect 902 1462 905 1468
rect 938 1458 942 1461
rect 894 1362 897 1418
rect 910 1392 913 1418
rect 926 1372 929 1458
rect 950 1452 953 1458
rect 946 1448 950 1451
rect 934 1372 937 1438
rect 942 1432 945 1438
rect 938 1368 942 1371
rect 838 1342 841 1348
rect 822 1338 833 1341
rect 774 1258 782 1261
rect 670 1168 681 1171
rect 694 1172 697 1178
rect 710 1171 713 1218
rect 718 1192 721 1228
rect 702 1168 713 1171
rect 670 1152 673 1168
rect 682 1158 686 1161
rect 702 1152 705 1168
rect 710 1152 713 1158
rect 646 1102 649 1118
rect 670 1112 673 1118
rect 702 1092 705 1118
rect 586 1068 593 1071
rect 526 1052 529 1068
rect 542 1062 545 1068
rect 554 1058 558 1061
rect 578 1058 582 1061
rect 590 1048 598 1051
rect 478 1042 481 1048
rect 490 1038 494 1041
rect 502 1032 505 1038
rect 478 992 481 998
rect 422 978 433 981
rect 422 962 425 968
rect 374 958 382 961
rect 326 952 329 958
rect 370 948 374 951
rect 318 938 329 941
rect 338 938 342 941
rect 326 892 329 938
rect 374 932 377 938
rect 346 928 350 931
rect 342 882 345 928
rect 382 882 385 958
rect 370 878 374 881
rect 310 872 313 878
rect 342 872 345 878
rect 246 861 249 868
rect 246 858 254 861
rect 262 852 265 868
rect 274 858 278 861
rect 314 858 318 861
rect 302 842 305 858
rect 342 852 345 858
rect 314 848 318 851
rect 330 848 337 851
rect 250 838 257 841
rect 254 831 257 838
rect 254 828 270 831
rect 158 762 161 818
rect 206 782 209 818
rect 158 742 161 758
rect 82 668 86 671
rect 38 662 41 668
rect 94 662 97 668
rect 34 648 38 651
rect 90 648 94 651
rect 102 642 105 668
rect 42 618 46 621
rect 14 492 17 568
rect 22 552 25 618
rect 30 562 33 618
rect 82 578 86 581
rect 54 572 57 578
rect 42 568 46 571
rect 62 562 65 578
rect 30 552 33 558
rect 110 552 113 678
rect 126 672 129 718
rect 122 658 126 661
rect 134 651 137 678
rect 166 662 169 748
rect 178 738 182 741
rect 226 738 230 741
rect 214 732 217 738
rect 174 662 177 718
rect 126 648 137 651
rect 102 548 110 551
rect 54 542 57 548
rect 22 532 25 538
rect 54 472 57 508
rect 70 502 73 538
rect 90 528 94 531
rect 78 482 81 488
rect 66 478 70 481
rect 38 462 41 468
rect 18 458 22 461
rect 6 452 9 458
rect 78 442 81 458
rect 26 438 30 441
rect 46 372 49 418
rect 94 392 97 498
rect 102 482 105 548
rect 118 492 121 608
rect 126 562 129 648
rect 158 642 161 658
rect 134 612 137 638
rect 134 522 137 598
rect 142 572 145 618
rect 150 572 153 578
rect 158 562 161 578
rect 166 572 169 618
rect 174 582 177 648
rect 182 562 185 648
rect 190 642 193 718
rect 230 682 233 738
rect 254 732 257 768
rect 278 752 281 838
rect 326 762 329 798
rect 334 792 337 848
rect 294 742 297 748
rect 318 732 321 738
rect 326 732 329 758
rect 358 752 361 878
rect 378 868 382 871
rect 366 832 369 868
rect 390 852 393 928
rect 406 852 409 958
rect 430 942 433 978
rect 466 968 470 971
rect 526 962 529 968
rect 558 962 561 1048
rect 582 1042 585 1048
rect 570 1038 574 1041
rect 590 991 593 1048
rect 622 1041 625 1068
rect 670 1062 673 1088
rect 718 1072 721 1178
rect 726 1092 729 1248
rect 734 1072 737 1158
rect 766 1072 769 1248
rect 790 1242 793 1318
rect 806 1272 809 1338
rect 814 1322 817 1328
rect 814 1292 817 1308
rect 830 1292 833 1338
rect 846 1332 849 1338
rect 846 1272 849 1328
rect 854 1292 857 1358
rect 890 1348 894 1351
rect 782 1142 785 1147
rect 798 1122 801 1218
rect 806 1192 809 1268
rect 862 1252 865 1348
rect 878 1332 881 1348
rect 902 1342 905 1348
rect 918 1342 921 1358
rect 926 1352 929 1368
rect 946 1358 950 1361
rect 958 1352 961 1378
rect 966 1372 969 1478
rect 998 1472 1001 1478
rect 986 1468 993 1471
rect 990 1462 993 1468
rect 978 1458 982 1461
rect 978 1448 985 1451
rect 974 1352 977 1358
rect 942 1342 945 1348
rect 834 1248 838 1251
rect 806 1172 809 1188
rect 886 1172 889 1258
rect 902 1192 905 1338
rect 974 1292 977 1338
rect 982 1322 985 1448
rect 998 1402 1001 1468
rect 1006 1422 1009 1518
rect 1014 1512 1017 1528
rect 1046 1522 1049 1528
rect 1062 1522 1065 1538
rect 1094 1532 1097 1538
rect 1118 1532 1121 1538
rect 1022 1482 1025 1488
rect 1030 1482 1033 1518
rect 1112 1503 1114 1507
rect 1118 1503 1121 1507
rect 1125 1503 1128 1507
rect 1102 1472 1105 1478
rect 1090 1468 1094 1471
rect 1122 1468 1126 1471
rect 1018 1458 1022 1461
rect 1038 1451 1041 1468
rect 1134 1462 1137 1528
rect 1142 1472 1145 1538
rect 1158 1462 1161 1468
rect 1058 1458 1062 1461
rect 1074 1458 1078 1461
rect 1034 1448 1041 1451
rect 1066 1448 1070 1451
rect 1014 1432 1017 1438
rect 994 1388 998 1391
rect 990 1362 993 1368
rect 998 1352 1001 1378
rect 1006 1362 1009 1418
rect 954 1278 958 1281
rect 914 1259 918 1262
rect 950 1192 953 1278
rect 982 1252 985 1318
rect 990 1292 993 1328
rect 1014 1292 1017 1398
rect 1030 1392 1033 1418
rect 1022 1372 1025 1388
rect 1038 1362 1041 1448
rect 1094 1442 1097 1448
rect 1078 1432 1081 1438
rect 1070 1428 1078 1431
rect 1022 1342 1025 1348
rect 1030 1292 1033 1338
rect 1038 1302 1041 1358
rect 1006 1272 1009 1278
rect 1014 1272 1017 1288
rect 1038 1282 1041 1288
rect 1046 1272 1049 1328
rect 990 1252 993 1258
rect 962 1248 966 1251
rect 1026 1248 1030 1251
rect 1046 1232 1049 1268
rect 1054 1242 1057 1408
rect 1062 1392 1065 1428
rect 914 1188 918 1191
rect 870 1152 873 1158
rect 838 1142 841 1147
rect 634 1058 638 1061
rect 646 1052 649 1058
rect 678 1052 681 1058
rect 682 1048 686 1051
rect 622 1038 630 1041
rect 638 1032 641 1048
rect 686 1038 694 1041
rect 662 1032 665 1038
rect 670 1032 673 1038
rect 600 1003 602 1007
rect 606 1003 609 1007
rect 613 1003 616 1007
rect 590 988 598 991
rect 578 968 582 971
rect 602 968 606 971
rect 482 958 486 961
rect 562 958 566 961
rect 454 952 457 958
rect 474 948 478 951
rect 570 948 574 951
rect 438 942 441 948
rect 558 942 561 948
rect 434 938 438 941
rect 522 938 526 941
rect 414 862 417 868
rect 398 822 401 848
rect 374 792 377 818
rect 390 812 393 818
rect 398 792 401 798
rect 414 772 417 848
rect 422 812 425 838
rect 266 728 270 731
rect 346 728 350 731
rect 242 718 249 721
rect 214 672 217 678
rect 230 672 233 678
rect 198 662 201 668
rect 246 652 249 718
rect 254 662 257 708
rect 278 682 281 718
rect 302 712 305 718
rect 266 678 270 681
rect 278 672 281 678
rect 334 672 337 728
rect 358 692 361 728
rect 366 682 369 718
rect 374 672 377 748
rect 390 692 393 758
rect 294 662 297 668
rect 306 658 310 661
rect 258 648 262 651
rect 298 648 302 651
rect 318 642 321 648
rect 214 632 217 638
rect 310 632 313 638
rect 334 632 337 668
rect 342 652 345 658
rect 386 648 390 651
rect 406 642 409 738
rect 414 732 417 768
rect 430 762 433 928
rect 494 902 497 928
rect 470 882 473 898
rect 514 878 518 881
rect 438 852 441 878
rect 446 852 449 858
rect 438 802 441 848
rect 470 842 473 878
rect 486 872 489 878
rect 486 852 489 858
rect 498 848 502 851
rect 490 838 494 841
rect 462 802 465 818
rect 502 792 505 818
rect 490 768 494 771
rect 446 762 449 768
rect 510 762 513 848
rect 518 832 521 868
rect 454 732 457 758
rect 478 752 481 758
rect 498 748 502 751
rect 526 742 529 928
rect 534 862 537 868
rect 542 832 545 938
rect 630 932 633 1018
rect 662 962 665 968
rect 678 942 681 978
rect 622 922 625 928
rect 622 882 625 918
rect 662 882 665 938
rect 686 892 689 1038
rect 702 1031 705 1058
rect 710 1052 713 1068
rect 694 1028 705 1031
rect 694 972 697 1028
rect 706 1018 710 1021
rect 718 991 721 1068
rect 718 988 729 991
rect 718 972 721 978
rect 710 962 713 968
rect 726 962 729 988
rect 718 942 721 948
rect 698 938 702 941
rect 578 878 582 881
rect 662 872 665 878
rect 702 872 705 928
rect 578 868 582 871
rect 554 858 558 861
rect 618 858 622 861
rect 570 848 574 851
rect 554 838 558 841
rect 626 838 630 841
rect 638 832 641 858
rect 678 842 681 848
rect 558 772 561 818
rect 600 803 602 807
rect 606 803 609 807
rect 613 803 616 807
rect 594 788 598 791
rect 642 788 646 791
rect 546 758 550 761
rect 570 748 574 751
rect 462 732 465 738
rect 522 728 526 731
rect 462 692 465 708
rect 422 682 425 688
rect 486 672 489 728
rect 494 682 497 688
rect 418 668 422 671
rect 498 668 502 671
rect 446 662 449 668
rect 526 662 529 728
rect 542 682 545 748
rect 582 741 585 768
rect 610 758 614 761
rect 590 752 593 758
rect 574 738 585 741
rect 550 722 553 728
rect 554 718 561 721
rect 558 672 561 718
rect 574 692 577 738
rect 590 692 593 728
rect 606 672 609 758
rect 630 732 633 768
rect 638 752 641 768
rect 646 762 649 768
rect 654 752 657 828
rect 670 822 673 828
rect 686 822 689 848
rect 694 792 697 818
rect 658 748 662 751
rect 646 692 649 728
rect 622 682 625 688
rect 670 682 673 718
rect 678 692 681 768
rect 686 732 689 768
rect 702 762 705 788
rect 698 748 705 751
rect 694 682 697 738
rect 702 692 705 748
rect 670 671 673 678
rect 666 668 673 671
rect 710 672 713 918
rect 726 912 729 958
rect 726 872 729 878
rect 722 858 726 861
rect 734 852 737 1058
rect 758 1052 761 1058
rect 778 1038 782 1041
rect 790 1032 793 1058
rect 802 1048 806 1051
rect 814 1042 817 1098
rect 822 1062 825 1068
rect 894 1062 897 1068
rect 838 1052 841 1058
rect 826 1048 830 1051
rect 846 1042 849 1058
rect 870 1052 873 1058
rect 878 1041 881 1058
rect 870 1038 881 1041
rect 854 1032 857 1038
rect 742 972 745 978
rect 750 962 753 1018
rect 790 1002 793 1018
rect 822 1012 825 1018
rect 842 988 846 991
rect 854 972 857 978
rect 834 968 838 971
rect 814 962 817 968
rect 802 958 806 961
rect 842 958 846 961
rect 862 952 865 1018
rect 870 992 873 1038
rect 878 992 881 1028
rect 886 1002 889 1038
rect 874 958 878 961
rect 746 948 750 951
rect 818 948 822 951
rect 798 942 801 948
rect 762 928 766 931
rect 774 922 777 938
rect 862 932 865 938
rect 866 928 873 931
rect 750 882 753 918
rect 798 902 801 928
rect 750 861 753 868
rect 746 858 753 861
rect 758 862 761 868
rect 766 852 769 858
rect 718 832 721 838
rect 726 792 729 838
rect 734 792 737 848
rect 750 802 753 838
rect 722 768 726 771
rect 738 758 742 761
rect 730 748 734 751
rect 746 748 750 751
rect 758 742 761 778
rect 774 742 777 888
rect 786 858 790 861
rect 794 848 798 851
rect 782 832 785 838
rect 790 752 793 818
rect 806 762 809 908
rect 838 882 841 928
rect 862 892 865 918
rect 870 872 873 928
rect 878 922 881 948
rect 886 892 889 968
rect 902 962 905 1168
rect 926 1152 929 1168
rect 1070 1151 1073 1428
rect 1086 1342 1089 1348
rect 1094 1342 1097 1348
rect 1110 1342 1113 1458
rect 1134 1452 1137 1458
rect 1134 1441 1137 1448
rect 1150 1442 1153 1458
rect 1166 1452 1169 1478
rect 1174 1472 1177 1498
rect 1198 1492 1201 1498
rect 1206 1481 1209 1518
rect 1198 1478 1209 1481
rect 1214 1482 1217 1538
rect 1222 1532 1225 1548
rect 1230 1532 1233 1538
rect 1182 1452 1185 1458
rect 1198 1452 1201 1478
rect 1206 1462 1209 1468
rect 1222 1462 1225 1518
rect 1230 1472 1233 1528
rect 1238 1522 1241 1538
rect 1250 1528 1254 1531
rect 1310 1531 1313 1538
rect 1306 1528 1313 1531
rect 1318 1532 1321 1548
rect 1326 1542 1329 1548
rect 1330 1528 1334 1531
rect 1134 1438 1145 1441
rect 1126 1392 1129 1438
rect 1134 1392 1137 1398
rect 1078 1332 1081 1338
rect 1110 1332 1113 1338
rect 1112 1303 1114 1307
rect 1118 1303 1121 1307
rect 1125 1303 1128 1307
rect 1118 1272 1121 1278
rect 1102 1263 1105 1268
rect 1142 1222 1145 1438
rect 1158 1432 1161 1448
rect 1206 1442 1209 1448
rect 1206 1352 1209 1438
rect 1222 1422 1225 1458
rect 1238 1452 1241 1488
rect 1270 1482 1273 1508
rect 1286 1482 1289 1528
rect 1342 1522 1345 1528
rect 1254 1462 1257 1468
rect 1246 1362 1249 1458
rect 1270 1452 1273 1458
rect 1254 1371 1257 1438
rect 1286 1412 1289 1418
rect 1286 1392 1289 1408
rect 1274 1388 1278 1391
rect 1294 1382 1297 1468
rect 1326 1462 1329 1468
rect 1302 1402 1305 1448
rect 1318 1442 1321 1458
rect 1326 1392 1329 1418
rect 1350 1392 1353 1538
rect 1366 1492 1369 1558
rect 1430 1552 1433 1558
rect 1374 1512 1377 1518
rect 1374 1492 1377 1508
rect 1358 1392 1361 1448
rect 1366 1402 1369 1458
rect 1382 1412 1385 1548
rect 1390 1422 1393 1538
rect 1414 1532 1417 1548
rect 1422 1532 1425 1538
rect 1438 1532 1441 1538
rect 1446 1522 1449 1548
rect 1454 1511 1457 1558
rect 1446 1508 1457 1511
rect 1446 1492 1449 1508
rect 1462 1502 1465 1568
rect 1478 1562 1481 1568
rect 1470 1552 1473 1558
rect 1518 1552 1521 1568
rect 1590 1562 1593 1568
rect 1554 1558 1558 1561
rect 1482 1548 1486 1551
rect 1470 1532 1473 1538
rect 1486 1512 1489 1548
rect 1494 1501 1497 1548
rect 1514 1538 1518 1541
rect 1526 1532 1529 1548
rect 1534 1522 1537 1558
rect 1594 1548 1598 1551
rect 1546 1538 1550 1541
rect 1486 1498 1497 1501
rect 1462 1472 1465 1498
rect 1486 1492 1489 1498
rect 1426 1468 1430 1471
rect 1450 1468 1454 1471
rect 1398 1462 1401 1468
rect 1406 1442 1409 1458
rect 1430 1452 1433 1458
rect 1422 1432 1425 1448
rect 1438 1412 1441 1468
rect 1462 1392 1465 1458
rect 1494 1422 1497 1468
rect 1390 1382 1393 1388
rect 1254 1368 1262 1371
rect 1266 1368 1270 1371
rect 1374 1362 1377 1368
rect 1306 1358 1310 1361
rect 1410 1358 1414 1361
rect 1162 1348 1166 1351
rect 1150 1342 1153 1348
rect 1182 1332 1185 1338
rect 1162 1328 1166 1331
rect 1218 1328 1222 1331
rect 1158 1292 1161 1298
rect 1150 1242 1153 1268
rect 1166 1252 1169 1318
rect 1174 1282 1177 1328
rect 1198 1322 1201 1328
rect 1238 1302 1241 1358
rect 1250 1348 1254 1351
rect 1330 1348 1334 1351
rect 1362 1348 1390 1351
rect 1442 1348 1449 1351
rect 1246 1292 1249 1308
rect 1182 1282 1185 1288
rect 1162 1148 1166 1151
rect 974 1112 977 1147
rect 990 1062 993 1138
rect 914 1058 918 1061
rect 926 1042 929 1048
rect 910 1032 913 1038
rect 966 1032 969 1058
rect 990 1052 993 1058
rect 1006 1052 1009 1118
rect 1030 1092 1033 1108
rect 1112 1103 1114 1107
rect 1118 1103 1121 1107
rect 1125 1103 1128 1107
rect 1114 1088 1118 1091
rect 1022 1082 1025 1088
rect 1046 1070 1049 1088
rect 1142 1072 1145 1128
rect 1174 1092 1177 1278
rect 1270 1272 1273 1318
rect 1278 1302 1281 1338
rect 1278 1262 1281 1278
rect 1194 1258 1198 1261
rect 1210 1258 1214 1261
rect 1234 1258 1238 1261
rect 1242 1248 1246 1251
rect 1214 1242 1217 1248
rect 1206 1192 1209 1238
rect 1214 1162 1217 1238
rect 1262 1232 1265 1258
rect 1286 1222 1289 1348
rect 1302 1311 1305 1338
rect 1314 1328 1321 1331
rect 1302 1308 1310 1311
rect 1294 1301 1297 1308
rect 1294 1298 1305 1301
rect 1294 1282 1297 1288
rect 1302 1282 1305 1298
rect 1310 1282 1313 1308
rect 1318 1282 1321 1328
rect 1326 1272 1329 1348
rect 1334 1332 1337 1338
rect 1342 1322 1345 1348
rect 1370 1338 1374 1341
rect 1402 1338 1406 1341
rect 1422 1322 1425 1348
rect 1430 1302 1433 1338
rect 1438 1332 1441 1338
rect 1362 1278 1366 1281
rect 1310 1262 1313 1268
rect 1358 1262 1361 1268
rect 1346 1258 1350 1261
rect 1222 1152 1225 1218
rect 1238 1152 1241 1158
rect 1246 1152 1249 1218
rect 1278 1152 1281 1158
rect 1302 1152 1305 1158
rect 1330 1148 1334 1151
rect 1206 1092 1209 1148
rect 1238 1122 1241 1138
rect 1066 1068 1070 1071
rect 1098 1058 1102 1061
rect 1070 1052 1073 1058
rect 1166 1052 1169 1058
rect 1190 1052 1193 1068
rect 910 992 913 998
rect 918 972 921 1018
rect 974 972 977 1018
rect 910 951 913 968
rect 990 962 993 1038
rect 1086 992 1089 1028
rect 902 948 913 951
rect 922 948 958 951
rect 978 948 982 951
rect 902 892 905 948
rect 930 928 934 931
rect 910 872 913 928
rect 942 892 945 938
rect 990 922 993 958
rect 998 952 1001 958
rect 1062 952 1065 968
rect 1094 952 1097 988
rect 1142 952 1145 1008
rect 1222 1002 1225 1058
rect 1022 942 1025 948
rect 1054 942 1057 948
rect 1202 947 1206 950
rect 1098 938 1102 941
rect 1162 938 1166 941
rect 826 868 830 871
rect 814 852 817 858
rect 814 792 817 838
rect 802 748 814 751
rect 774 732 777 738
rect 734 682 737 708
rect 758 692 761 718
rect 766 682 769 728
rect 798 692 801 728
rect 822 722 825 768
rect 830 692 833 858
rect 838 782 841 868
rect 934 862 937 878
rect 962 858 966 861
rect 946 848 950 851
rect 846 792 849 838
rect 862 792 865 828
rect 870 792 873 848
rect 886 842 889 848
rect 894 832 897 848
rect 926 842 929 848
rect 954 838 958 841
rect 926 792 929 828
rect 934 802 937 818
rect 950 772 953 778
rect 938 768 942 771
rect 958 762 961 768
rect 966 762 969 818
rect 974 772 977 848
rect 982 792 985 918
rect 990 842 993 878
rect 1006 872 1009 938
rect 1046 932 1049 938
rect 998 862 1001 868
rect 998 812 1001 818
rect 998 752 1001 788
rect 1006 772 1009 848
rect 946 748 950 751
rect 962 748 966 751
rect 986 748 990 751
rect 838 732 841 738
rect 854 712 857 728
rect 722 678 726 681
rect 714 668 718 671
rect 534 662 537 668
rect 470 652 473 658
rect 582 652 585 658
rect 490 648 494 651
rect 506 648 510 651
rect 462 642 465 648
rect 526 642 529 648
rect 418 638 422 641
rect 546 638 550 641
rect 190 572 193 618
rect 238 612 241 618
rect 234 588 238 591
rect 274 588 278 591
rect 198 562 201 578
rect 206 552 209 588
rect 214 572 217 578
rect 246 572 249 588
rect 274 568 278 571
rect 258 558 262 561
rect 230 552 233 558
rect 294 552 297 558
rect 194 548 198 551
rect 242 548 246 551
rect 274 548 278 551
rect 150 542 153 548
rect 182 542 185 548
rect 310 542 313 618
rect 170 538 174 541
rect 218 528 222 531
rect 102 472 105 478
rect 110 472 113 478
rect 102 462 105 468
rect 126 452 129 518
rect 134 482 137 518
rect 150 472 153 518
rect 262 492 265 538
rect 318 532 321 628
rect 406 602 409 638
rect 558 592 561 648
rect 574 642 577 648
rect 582 592 585 638
rect 590 602 593 618
rect 600 603 602 607
rect 606 603 609 607
rect 613 603 616 607
rect 450 588 454 591
rect 350 562 353 568
rect 358 552 361 578
rect 382 562 385 568
rect 414 562 417 568
rect 386 548 390 551
rect 418 548 422 551
rect 326 532 329 548
rect 462 542 465 588
rect 526 552 529 578
rect 566 568 574 571
rect 494 542 497 547
rect 394 538 398 541
rect 318 522 321 528
rect 334 512 337 538
rect 354 528 358 531
rect 162 488 166 491
rect 282 478 286 481
rect 150 462 153 468
rect 186 458 190 461
rect 162 448 166 451
rect 178 448 182 451
rect 150 442 153 448
rect 198 441 201 478
rect 230 472 233 478
rect 222 462 225 468
rect 210 458 214 461
rect 194 438 201 441
rect 118 392 121 438
rect 182 422 185 428
rect 18 368 22 371
rect 70 362 73 388
rect 58 358 62 361
rect 10 338 14 341
rect 6 282 9 298
rect 14 192 17 328
rect 22 322 25 348
rect 30 332 33 358
rect 74 348 78 351
rect 46 342 49 348
rect 54 342 57 348
rect 22 292 25 308
rect 46 292 49 318
rect 86 292 89 368
rect 110 352 113 368
rect 126 362 129 388
rect 122 348 126 351
rect 70 282 73 288
rect 110 282 113 288
rect 38 272 41 278
rect 62 272 65 278
rect 14 92 17 168
rect 22 162 25 178
rect 34 168 38 171
rect 54 162 57 188
rect 62 172 65 268
rect 122 258 126 261
rect 82 238 86 241
rect 22 142 25 158
rect 62 152 65 158
rect 50 148 54 151
rect 22 82 25 138
rect 46 132 49 138
rect 70 92 73 238
rect 94 232 97 258
rect 102 242 105 248
rect 78 142 81 198
rect 110 192 113 258
rect 134 252 137 408
rect 150 392 153 398
rect 158 362 161 388
rect 166 352 169 358
rect 174 352 177 378
rect 182 362 185 368
rect 198 362 201 368
rect 150 292 153 348
rect 182 292 185 348
rect 206 341 209 448
rect 238 392 241 448
rect 246 422 249 458
rect 254 432 257 438
rect 230 372 233 378
rect 242 368 249 371
rect 226 358 230 361
rect 214 352 217 358
rect 202 338 209 341
rect 194 258 198 261
rect 134 242 137 248
rect 142 242 145 258
rect 162 248 166 251
rect 86 132 89 168
rect 102 132 105 168
rect 126 152 129 158
rect 110 142 113 148
rect 134 142 137 238
rect 150 192 153 238
rect 174 222 177 258
rect 182 212 185 238
rect 198 192 201 238
rect 206 182 209 338
rect 222 332 225 358
rect 234 348 238 351
rect 246 332 249 368
rect 254 342 257 348
rect 214 292 217 318
rect 222 252 225 328
rect 270 322 273 468
rect 346 458 358 461
rect 286 452 289 458
rect 294 412 297 448
rect 302 431 305 458
rect 330 448 334 451
rect 314 438 318 441
rect 346 438 350 441
rect 334 432 337 438
rect 302 428 313 431
rect 302 412 305 418
rect 310 392 313 428
rect 366 402 369 538
rect 414 532 417 538
rect 386 528 390 531
rect 374 472 377 518
rect 430 502 433 538
rect 442 528 446 531
rect 486 482 489 508
rect 498 478 502 481
rect 538 478 545 481
rect 382 472 385 478
rect 414 472 417 478
rect 438 472 441 478
rect 470 472 473 478
rect 406 452 409 468
rect 454 462 457 468
rect 438 452 441 458
rect 470 452 473 458
rect 458 448 462 451
rect 442 438 446 441
rect 518 432 521 438
rect 278 342 281 388
rect 398 382 401 418
rect 302 372 305 378
rect 422 362 425 418
rect 290 358 294 361
rect 394 358 398 361
rect 318 352 321 358
rect 290 348 294 351
rect 390 342 393 348
rect 278 282 281 328
rect 334 322 337 338
rect 382 332 385 338
rect 362 328 366 331
rect 342 292 345 328
rect 406 292 409 348
rect 430 332 433 418
rect 526 392 529 428
rect 470 368 478 371
rect 438 332 441 358
rect 462 342 465 348
rect 302 282 305 288
rect 390 282 393 288
rect 282 278 286 281
rect 274 268 278 271
rect 230 242 233 268
rect 242 258 254 261
rect 282 258 286 261
rect 234 228 238 231
rect 238 192 241 208
rect 142 162 145 178
rect 194 168 198 171
rect 86 82 89 128
rect 118 82 121 98
rect 126 82 129 88
rect 46 72 49 78
rect 86 72 89 78
rect 10 68 14 71
rect 34 68 38 71
rect 86 61 89 68
rect 86 58 94 61
rect 22 52 25 58
rect 34 48 38 51
rect 74 48 78 51
rect 46 12 49 48
rect 134 12 137 68
rect 46 -18 49 8
rect 46 -22 50 -18
rect 134 -19 138 -18
rect 142 -19 145 98
rect 150 92 153 148
rect 158 142 161 168
rect 206 162 209 178
rect 214 172 217 178
rect 222 162 225 168
rect 178 158 182 161
rect 234 158 238 161
rect 186 148 190 151
rect 206 142 209 158
rect 238 142 241 148
rect 246 142 249 168
rect 174 92 177 128
rect 166 82 169 88
rect 206 72 209 138
rect 230 92 233 138
rect 254 82 257 208
rect 262 162 265 248
rect 270 192 273 218
rect 282 168 286 171
rect 294 152 297 258
rect 326 252 329 278
rect 398 272 401 278
rect 406 272 409 278
rect 366 262 369 268
rect 346 258 350 261
rect 338 248 342 251
rect 310 242 313 248
rect 274 148 278 151
rect 270 92 273 138
rect 194 68 198 71
rect 258 68 262 71
rect 282 68 286 71
rect 222 62 225 68
rect 294 62 297 148
rect 302 92 305 168
rect 318 162 321 248
rect 354 238 361 241
rect 342 232 345 238
rect 326 182 329 188
rect 338 168 345 171
rect 330 148 334 151
rect 310 132 313 138
rect 342 92 345 168
rect 350 152 353 158
rect 358 92 361 238
rect 374 142 377 178
rect 390 162 393 268
rect 414 212 417 278
rect 438 271 441 328
rect 446 322 449 338
rect 454 282 457 328
rect 470 292 473 368
rect 494 362 497 378
rect 482 348 486 351
rect 486 332 489 338
rect 502 322 505 328
rect 498 278 502 281
rect 438 268 446 271
rect 502 262 505 268
rect 450 248 454 251
rect 414 192 417 208
rect 494 192 497 218
rect 458 168 462 171
rect 382 152 385 158
rect 414 142 417 148
rect 446 142 449 148
rect 402 138 406 141
rect 434 138 438 141
rect 454 132 457 148
rect 370 128 374 131
rect 402 128 406 131
rect 434 128 438 131
rect 458 128 465 131
rect 322 78 326 81
rect 322 68 326 71
rect 346 68 350 71
rect 362 68 366 71
rect 162 58 166 61
rect 202 58 206 61
rect 174 42 177 48
rect 278 22 281 48
rect 134 -22 145 -19
rect 158 -18 161 8
rect 294 -18 297 58
rect 374 52 377 68
rect 414 62 417 128
rect 426 68 430 71
rect 390 52 393 58
rect 422 52 425 58
rect 346 48 350 51
rect 414 42 417 48
rect 438 32 441 78
rect 454 52 457 78
rect 462 72 465 128
rect 470 92 473 158
rect 478 142 481 148
rect 502 142 505 168
rect 510 162 513 378
rect 534 362 537 468
rect 542 372 545 478
rect 558 442 561 448
rect 566 431 569 568
rect 590 562 593 598
rect 702 592 705 638
rect 726 592 729 668
rect 734 632 737 678
rect 766 672 769 678
rect 774 672 777 678
rect 806 672 809 678
rect 886 671 889 740
rect 894 682 897 738
rect 910 682 913 748
rect 1022 742 1025 928
rect 1038 891 1041 918
rect 1038 888 1049 891
rect 1038 872 1041 878
rect 1038 792 1041 868
rect 1046 862 1049 888
rect 974 712 977 738
rect 990 732 993 738
rect 886 668 897 671
rect 938 668 942 671
rect 670 552 673 578
rect 714 568 718 571
rect 734 562 737 618
rect 758 592 761 628
rect 774 592 777 668
rect 782 652 785 658
rect 814 642 817 658
rect 798 592 801 618
rect 862 602 865 659
rect 886 572 889 658
rect 894 592 897 668
rect 930 658 934 661
rect 746 568 750 571
rect 762 558 766 561
rect 578 548 582 551
rect 638 542 641 547
rect 614 472 617 478
rect 638 472 641 478
rect 582 452 585 458
rect 590 442 593 448
rect 606 442 609 448
rect 558 428 569 431
rect 574 432 577 438
rect 558 392 561 428
rect 590 382 593 438
rect 600 403 602 407
rect 606 403 609 407
rect 613 403 616 407
rect 622 392 625 468
rect 646 392 649 498
rect 702 492 705 538
rect 726 532 729 548
rect 758 542 761 548
rect 782 542 785 548
rect 662 462 665 468
rect 718 462 721 468
rect 678 458 686 461
rect 678 452 681 458
rect 714 448 718 451
rect 670 442 673 448
rect 654 432 657 438
rect 534 342 537 358
rect 534 322 537 338
rect 550 332 553 368
rect 562 358 566 361
rect 626 358 630 361
rect 558 342 561 348
rect 566 292 569 348
rect 574 342 577 358
rect 614 342 617 348
rect 578 328 582 331
rect 590 292 593 318
rect 598 272 601 338
rect 522 258 526 261
rect 538 258 542 261
rect 550 252 553 268
rect 614 262 617 338
rect 638 292 641 368
rect 654 362 657 378
rect 662 362 665 418
rect 670 412 673 438
rect 678 392 681 428
rect 686 382 689 448
rect 726 442 729 478
rect 758 472 761 518
rect 790 502 793 568
rect 830 551 833 558
rect 862 552 865 568
rect 950 552 953 688
rect 958 672 961 678
rect 966 672 969 678
rect 982 672 985 678
rect 990 672 993 728
rect 1006 722 1009 738
rect 1026 728 1030 731
rect 1014 692 1017 718
rect 974 662 977 668
rect 1002 658 1006 661
rect 958 652 961 658
rect 990 592 993 658
rect 998 592 1001 638
rect 958 552 961 568
rect 798 482 801 508
rect 950 482 953 528
rect 1006 502 1009 538
rect 786 478 790 481
rect 938 478 942 481
rect 894 472 897 478
rect 746 468 750 471
rect 826 468 830 471
rect 698 438 702 441
rect 718 391 721 418
rect 710 388 721 391
rect 742 392 745 428
rect 650 358 654 361
rect 670 351 673 368
rect 686 362 689 378
rect 710 372 713 388
rect 722 378 726 381
rect 694 352 697 358
rect 702 352 705 358
rect 662 348 673 351
rect 646 342 649 348
rect 662 292 665 348
rect 678 332 681 348
rect 734 342 737 368
rect 762 358 766 361
rect 750 352 753 358
rect 774 352 777 468
rect 886 462 889 468
rect 918 462 921 468
rect 858 458 870 461
rect 814 452 817 458
rect 934 452 937 458
rect 922 448 926 451
rect 762 348 766 351
rect 778 348 793 351
rect 742 322 745 348
rect 750 292 753 328
rect 766 292 769 338
rect 678 282 681 288
rect 698 278 702 281
rect 570 258 574 261
rect 626 258 630 261
rect 582 252 585 258
rect 610 248 614 251
rect 534 242 537 248
rect 542 232 545 238
rect 566 232 569 238
rect 574 192 577 248
rect 622 222 625 258
rect 514 148 518 151
rect 526 142 529 148
rect 542 142 545 158
rect 486 132 489 138
rect 494 82 497 118
rect 518 92 521 138
rect 550 82 553 128
rect 558 92 561 158
rect 582 152 585 168
rect 574 92 577 148
rect 478 62 481 68
rect 478 42 481 48
rect 510 32 513 78
rect 542 72 545 78
rect 582 72 585 78
rect 590 62 593 218
rect 600 203 602 207
rect 606 203 609 207
rect 613 203 616 207
rect 638 172 641 278
rect 650 268 654 271
rect 674 268 678 271
rect 690 258 694 261
rect 638 152 641 168
rect 622 132 625 138
rect 618 128 622 131
rect 598 122 601 128
rect 646 92 649 168
rect 654 152 657 248
rect 670 192 673 248
rect 674 168 678 171
rect 662 152 665 158
rect 686 152 689 168
rect 694 162 697 208
rect 710 182 713 268
rect 734 252 737 278
rect 734 212 737 248
rect 742 242 745 258
rect 750 231 753 238
rect 742 228 753 231
rect 734 172 737 208
rect 726 162 729 168
rect 670 92 673 108
rect 694 92 697 148
rect 710 142 713 158
rect 734 152 737 158
rect 742 132 745 228
rect 750 192 753 218
rect 758 152 761 288
rect 782 272 785 338
rect 790 292 793 348
rect 798 332 801 418
rect 814 392 817 408
rect 822 362 825 418
rect 814 282 817 318
rect 822 292 825 348
rect 830 342 833 448
rect 902 442 905 448
rect 966 442 969 468
rect 974 442 977 458
rect 990 452 993 498
rect 1014 492 1017 628
rect 1022 592 1025 668
rect 1042 659 1046 662
rect 1022 572 1025 588
rect 1034 468 1038 471
rect 1022 462 1025 468
rect 1046 462 1049 468
rect 1002 458 1006 461
rect 858 438 862 441
rect 846 432 849 438
rect 894 392 897 408
rect 858 378 862 381
rect 886 362 889 368
rect 898 358 902 361
rect 910 342 913 398
rect 950 372 953 408
rect 958 392 961 438
rect 982 382 985 448
rect 974 371 977 378
rect 974 368 982 371
rect 970 358 974 361
rect 934 352 937 358
rect 954 348 958 351
rect 990 342 993 348
rect 866 338 870 341
rect 890 338 894 341
rect 978 338 982 341
rect 910 332 913 338
rect 834 328 838 331
rect 866 328 870 331
rect 918 322 921 338
rect 910 301 913 318
rect 918 312 921 318
rect 910 298 921 301
rect 850 278 854 281
rect 858 268 865 271
rect 802 258 806 261
rect 766 222 769 248
rect 782 132 785 148
rect 790 132 793 138
rect 654 82 657 88
rect 702 82 705 128
rect 726 92 729 118
rect 758 92 761 128
rect 774 102 777 128
rect 610 78 614 81
rect 678 62 681 78
rect 710 72 713 78
rect 742 72 745 78
rect 750 72 753 78
rect 782 62 785 78
rect 798 61 801 258
rect 810 248 814 251
rect 822 192 825 258
rect 830 222 833 238
rect 814 162 817 168
rect 806 152 809 158
rect 814 152 817 158
rect 822 152 825 158
rect 830 122 833 168
rect 838 92 841 168
rect 846 162 849 268
rect 854 192 857 218
rect 862 202 865 268
rect 870 252 873 258
rect 878 192 881 278
rect 894 272 897 278
rect 886 262 889 268
rect 858 168 862 171
rect 878 162 881 168
rect 846 121 849 158
rect 854 152 857 158
rect 894 151 897 268
rect 906 218 910 221
rect 918 192 921 298
rect 926 282 929 298
rect 982 292 985 308
rect 998 292 1001 358
rect 1006 352 1009 358
rect 1014 292 1017 458
rect 1022 442 1025 448
rect 1046 402 1049 458
rect 1058 448 1062 451
rect 1022 342 1025 358
rect 1030 332 1033 368
rect 1046 362 1049 398
rect 1062 372 1065 408
rect 1070 392 1073 938
rect 1090 928 1094 931
rect 1114 918 1118 921
rect 1112 903 1114 907
rect 1118 903 1121 907
rect 1125 903 1128 907
rect 1134 891 1137 928
rect 1130 888 1137 891
rect 1138 868 1142 871
rect 1114 858 1118 861
rect 1094 742 1097 838
rect 1094 642 1097 738
rect 1110 732 1113 818
rect 1118 772 1121 848
rect 1118 752 1121 768
rect 1102 682 1105 718
rect 1112 703 1114 707
rect 1118 703 1121 707
rect 1125 703 1128 707
rect 1114 688 1118 691
rect 1150 672 1153 938
rect 1162 928 1166 931
rect 1182 921 1185 938
rect 1174 918 1185 921
rect 1166 892 1169 908
rect 1174 882 1177 918
rect 1194 888 1198 891
rect 1182 870 1185 888
rect 1230 872 1233 1068
rect 1238 1022 1241 1068
rect 1246 1062 1249 1148
rect 1254 1062 1257 1118
rect 1246 1012 1249 1058
rect 1262 1022 1265 1128
rect 1270 1122 1273 1138
rect 1294 1122 1297 1148
rect 1318 1122 1321 1128
rect 1278 1062 1281 1078
rect 1294 1071 1297 1118
rect 1306 1078 1310 1081
rect 1294 1068 1302 1071
rect 1326 1062 1329 1138
rect 1342 1092 1345 1228
rect 1374 1222 1377 1278
rect 1382 1272 1385 1288
rect 1414 1272 1417 1288
rect 1446 1282 1449 1348
rect 1470 1341 1473 1368
rect 1478 1352 1481 1398
rect 1502 1372 1505 1458
rect 1510 1442 1513 1478
rect 1542 1462 1545 1508
rect 1550 1472 1553 1528
rect 1566 1472 1569 1538
rect 1574 1492 1577 1548
rect 1598 1512 1601 1538
rect 1614 1532 1617 1558
rect 1646 1542 1649 1547
rect 1606 1492 1609 1518
rect 1614 1482 1617 1518
rect 1510 1392 1513 1438
rect 1526 1402 1529 1458
rect 1550 1442 1553 1468
rect 1558 1442 1561 1448
rect 1574 1432 1577 1458
rect 1586 1448 1590 1451
rect 1550 1392 1553 1398
rect 1534 1382 1537 1388
rect 1574 1382 1577 1418
rect 1590 1392 1593 1408
rect 1598 1372 1601 1478
rect 1654 1472 1657 1538
rect 1658 1468 1662 1471
rect 1658 1458 1662 1461
rect 1614 1442 1617 1458
rect 1614 1422 1617 1438
rect 1670 1392 1673 1438
rect 1678 1432 1681 1528
rect 1578 1368 1582 1371
rect 1630 1362 1633 1368
rect 1514 1358 1518 1361
rect 1682 1358 1686 1361
rect 1470 1338 1481 1341
rect 1458 1328 1462 1331
rect 1426 1278 1430 1281
rect 1398 1232 1401 1248
rect 1350 1162 1353 1218
rect 1390 1162 1393 1218
rect 1438 1192 1441 1268
rect 1446 1232 1449 1248
rect 1454 1192 1457 1298
rect 1470 1282 1473 1308
rect 1478 1292 1481 1338
rect 1494 1302 1497 1358
rect 1486 1272 1489 1278
rect 1510 1271 1513 1338
rect 1534 1281 1537 1348
rect 1562 1340 1566 1343
rect 1582 1342 1585 1358
rect 1590 1352 1593 1358
rect 1666 1348 1670 1351
rect 1646 1342 1649 1348
rect 1654 1342 1657 1348
rect 1694 1342 1697 1478
rect 1626 1338 1630 1341
rect 1666 1338 1670 1341
rect 1542 1302 1545 1338
rect 1546 1288 1550 1291
rect 1534 1278 1545 1281
rect 1506 1268 1513 1271
rect 1362 1158 1369 1161
rect 1354 1148 1358 1151
rect 1358 1072 1361 1118
rect 1366 1072 1369 1158
rect 1406 1152 1409 1158
rect 1410 1148 1417 1151
rect 1274 1058 1278 1061
rect 1298 1058 1302 1061
rect 1262 992 1265 998
rect 1270 992 1273 998
rect 1286 902 1289 1018
rect 1302 952 1305 1048
rect 1194 868 1198 871
rect 1158 852 1161 858
rect 1166 742 1169 747
rect 1230 741 1233 868
rect 1254 862 1257 898
rect 1318 892 1321 1038
rect 1334 1032 1337 1068
rect 1374 1052 1377 1148
rect 1414 1142 1417 1148
rect 1438 1148 1446 1151
rect 1462 1151 1465 1268
rect 1494 1172 1497 1258
rect 1470 1162 1473 1168
rect 1478 1152 1481 1158
rect 1494 1152 1497 1168
rect 1510 1162 1513 1268
rect 1534 1262 1537 1268
rect 1518 1172 1521 1248
rect 1526 1162 1529 1168
rect 1514 1158 1518 1161
rect 1542 1152 1545 1278
rect 1550 1272 1553 1278
rect 1558 1192 1561 1258
rect 1566 1252 1569 1318
rect 1574 1302 1577 1338
rect 1582 1272 1585 1288
rect 1590 1252 1593 1298
rect 1598 1292 1601 1338
rect 1614 1322 1617 1328
rect 1630 1312 1633 1328
rect 1614 1272 1617 1278
rect 1662 1272 1665 1318
rect 1622 1268 1630 1271
rect 1606 1262 1609 1268
rect 1622 1262 1625 1268
rect 1610 1248 1614 1251
rect 1566 1242 1569 1248
rect 1582 1162 1585 1168
rect 1462 1148 1470 1151
rect 1402 1138 1406 1141
rect 1382 1122 1385 1138
rect 1422 1132 1425 1140
rect 1406 1092 1409 1128
rect 1414 1082 1417 1088
rect 1422 1082 1425 1118
rect 1382 1072 1385 1078
rect 1394 1068 1398 1071
rect 1370 1048 1374 1051
rect 1366 962 1369 1008
rect 1374 992 1377 1028
rect 1382 992 1385 1018
rect 1390 992 1393 1048
rect 1426 988 1430 991
rect 1326 942 1329 948
rect 1350 942 1353 948
rect 1366 892 1369 958
rect 1382 942 1385 988
rect 1438 981 1441 1148
rect 1446 1132 1449 1138
rect 1454 1042 1457 1059
rect 1430 978 1441 981
rect 1402 948 1406 951
rect 1294 872 1297 878
rect 1262 792 1265 848
rect 1278 832 1281 868
rect 1298 858 1302 861
rect 1334 832 1337 868
rect 1350 852 1353 859
rect 1238 751 1241 758
rect 1238 748 1246 751
rect 1278 742 1281 828
rect 1398 792 1401 928
rect 1422 922 1425 928
rect 1410 888 1414 891
rect 1422 882 1425 898
rect 1430 892 1433 978
rect 1438 872 1441 878
rect 1446 862 1449 958
rect 1462 952 1465 1068
rect 1454 872 1457 908
rect 1478 872 1481 1148
rect 1542 1142 1545 1148
rect 1566 1142 1569 1158
rect 1606 1152 1609 1158
rect 1614 1152 1617 1238
rect 1598 1142 1601 1148
rect 1622 1142 1625 1258
rect 1662 1142 1665 1268
rect 1670 1262 1673 1268
rect 1674 1148 1678 1151
rect 1522 1138 1526 1141
rect 1618 1138 1622 1141
rect 1502 1132 1505 1138
rect 1510 962 1513 1118
rect 1518 1092 1521 1138
rect 1550 1132 1553 1138
rect 1574 1132 1577 1138
rect 1526 1092 1529 1128
rect 1654 1072 1657 1128
rect 1710 1112 1713 1418
rect 1718 1352 1721 1358
rect 1718 1152 1721 1318
rect 1558 952 1561 1058
rect 1590 1042 1593 1059
rect 1362 788 1366 791
rect 1366 752 1369 758
rect 1398 752 1401 768
rect 1438 752 1441 798
rect 1230 738 1238 741
rect 1094 582 1097 638
rect 1102 592 1105 668
rect 1110 642 1113 668
rect 1166 592 1169 718
rect 1182 692 1185 738
rect 1182 672 1185 688
rect 1278 682 1281 738
rect 1294 692 1297 747
rect 1206 672 1209 678
rect 1334 672 1337 678
rect 1286 662 1289 668
rect 1318 662 1321 668
rect 1222 652 1225 659
rect 1306 658 1310 661
rect 1362 658 1366 661
rect 1374 592 1377 738
rect 1394 728 1398 731
rect 1382 662 1385 718
rect 1422 692 1425 738
rect 1430 732 1433 738
rect 1422 672 1425 688
rect 1422 658 1430 661
rect 1422 652 1425 658
rect 1338 588 1342 591
rect 1078 542 1081 578
rect 1090 568 1094 571
rect 1178 568 1182 571
rect 1154 558 1158 561
rect 1078 362 1081 498
rect 1086 462 1089 538
rect 1086 442 1089 448
rect 1094 392 1097 548
rect 1102 502 1105 558
rect 1154 548 1158 551
rect 1122 538 1126 541
rect 1166 512 1169 548
rect 1190 532 1193 568
rect 1342 558 1350 561
rect 1226 548 1230 551
rect 1342 542 1345 558
rect 1358 552 1361 578
rect 1422 572 1425 578
rect 1430 572 1433 578
rect 1366 562 1369 568
rect 1426 558 1430 561
rect 1406 552 1409 558
rect 1226 538 1230 541
rect 1250 538 1254 541
rect 1290 538 1294 541
rect 1374 538 1382 541
rect 1112 503 1114 507
rect 1118 503 1121 507
rect 1125 503 1128 507
rect 1206 502 1209 518
rect 1110 432 1113 478
rect 1110 422 1113 428
rect 1094 362 1097 378
rect 1102 372 1105 398
rect 1082 358 1086 361
rect 1042 348 1046 351
rect 1074 348 1081 351
rect 1038 302 1041 328
rect 950 272 953 278
rect 950 252 953 258
rect 958 252 961 288
rect 982 262 985 268
rect 1006 262 1009 268
rect 1002 248 1006 251
rect 942 222 945 238
rect 930 168 934 171
rect 886 148 897 151
rect 910 152 913 158
rect 942 152 945 158
rect 922 148 926 151
rect 846 118 854 121
rect 806 82 809 88
rect 846 82 849 108
rect 878 92 881 118
rect 854 82 857 88
rect 858 78 865 81
rect 814 72 817 78
rect 846 72 849 78
rect 794 58 801 61
rect 558 52 561 58
rect 566 42 569 48
rect 686 22 689 48
rect 450 18 454 21
rect 798 12 801 58
rect 600 3 602 7
rect 606 3 609 7
rect 613 3 616 7
rect 158 -22 162 -18
rect 294 -22 298 -18
rect 790 -19 793 8
rect 814 -18 817 8
rect 838 -18 841 68
rect 862 -18 865 78
rect 886 72 889 148
rect 958 142 961 198
rect 974 162 977 168
rect 894 132 897 138
rect 902 112 905 128
rect 910 92 913 128
rect 966 112 969 128
rect 998 121 1001 238
rect 1014 192 1017 238
rect 1030 212 1033 278
rect 1038 182 1041 298
rect 1054 292 1057 298
rect 1078 292 1081 348
rect 1094 342 1097 348
rect 1126 332 1129 458
rect 1134 452 1137 468
rect 1170 458 1174 461
rect 1154 448 1158 451
rect 1142 362 1145 418
rect 1066 268 1070 271
rect 1086 271 1089 328
rect 1112 303 1114 307
rect 1118 303 1121 307
rect 1125 303 1128 307
rect 1078 268 1089 271
rect 1102 272 1105 278
rect 1078 252 1081 268
rect 1090 258 1097 261
rect 1006 132 1009 178
rect 1018 168 1022 171
rect 1042 158 1046 161
rect 1010 128 1017 131
rect 998 118 1009 121
rect 1006 92 1009 118
rect 918 78 926 81
rect 962 78 966 81
rect 918 32 921 78
rect 930 68 934 71
rect 962 68 966 71
rect 990 62 993 88
rect 998 72 1001 78
rect 978 58 982 61
rect 958 51 961 58
rect 1006 52 1009 58
rect 958 48 974 51
rect 918 12 921 28
rect 950 22 953 48
rect 918 -18 921 8
rect 982 -18 985 8
rect 798 -19 802 -18
rect 790 -22 802 -19
rect 814 -22 818 -18
rect 838 -22 842 -18
rect 862 -22 866 -18
rect 918 -22 922 -18
rect 982 -22 986 -18
rect 1014 -19 1017 128
rect 1022 72 1025 158
rect 1034 148 1038 151
rect 1054 142 1057 238
rect 1086 222 1089 238
rect 1078 192 1081 218
rect 1094 192 1097 258
rect 1110 212 1113 288
rect 1126 262 1129 268
rect 1134 232 1137 338
rect 1142 292 1145 358
rect 1150 272 1153 448
rect 1182 441 1185 498
rect 1214 482 1217 538
rect 1282 528 1286 531
rect 1270 511 1273 518
rect 1266 508 1273 511
rect 1230 492 1233 508
rect 1286 502 1289 528
rect 1206 472 1209 478
rect 1210 468 1214 471
rect 1190 462 1193 468
rect 1234 458 1238 461
rect 1266 458 1270 461
rect 1298 458 1302 461
rect 1178 438 1185 441
rect 1250 448 1254 451
rect 1278 448 1286 451
rect 1166 402 1169 418
rect 1206 392 1209 408
rect 1162 338 1166 341
rect 1174 312 1177 368
rect 1198 362 1201 378
rect 1186 358 1190 361
rect 1182 342 1185 348
rect 1206 342 1209 348
rect 1190 331 1193 338
rect 1186 328 1193 331
rect 1214 302 1217 368
rect 1230 342 1233 448
rect 1270 442 1273 448
rect 1242 438 1246 441
rect 1262 432 1265 438
rect 1254 392 1257 418
rect 1242 378 1246 381
rect 1254 342 1257 348
rect 1230 332 1233 338
rect 1174 292 1177 298
rect 1262 292 1265 368
rect 1278 362 1281 448
rect 1310 441 1313 518
rect 1326 492 1329 528
rect 1334 472 1337 518
rect 1306 438 1313 441
rect 1318 442 1321 448
rect 1342 442 1345 538
rect 1350 482 1353 538
rect 1374 472 1377 538
rect 1386 528 1393 531
rect 1390 482 1393 528
rect 1422 492 1425 548
rect 1438 532 1441 738
rect 1446 692 1449 848
rect 1454 842 1457 868
rect 1486 852 1489 948
rect 1510 942 1513 948
rect 1526 942 1529 948
rect 1510 892 1513 918
rect 1590 912 1593 938
rect 1526 892 1529 898
rect 1606 872 1609 938
rect 1630 922 1633 1068
rect 1646 1052 1649 1059
rect 1646 892 1649 948
rect 1654 892 1657 1038
rect 1682 978 1686 981
rect 1694 971 1697 1108
rect 1686 968 1697 971
rect 1702 1018 1710 1021
rect 1626 868 1630 871
rect 1674 868 1678 871
rect 1462 762 1465 768
rect 1470 752 1473 808
rect 1522 748 1526 751
rect 1558 751 1561 758
rect 1522 738 1526 741
rect 1478 732 1481 738
rect 1494 732 1497 738
rect 1458 728 1462 731
rect 1470 662 1473 668
rect 1486 652 1489 718
rect 1510 662 1513 718
rect 1574 692 1577 858
rect 1590 752 1593 868
rect 1686 862 1689 968
rect 1622 858 1630 861
rect 1622 792 1625 858
rect 1534 672 1537 678
rect 1550 672 1553 688
rect 1590 672 1593 748
rect 1638 672 1641 738
rect 1590 662 1593 668
rect 1554 658 1558 661
rect 1606 652 1609 659
rect 1654 592 1657 848
rect 1662 752 1665 788
rect 1670 692 1673 858
rect 1678 662 1681 858
rect 1694 792 1697 918
rect 1702 862 1705 1018
rect 1718 951 1721 1118
rect 1714 948 1721 951
rect 1714 938 1718 941
rect 1710 852 1713 898
rect 1718 892 1721 918
rect 1726 892 1729 1218
rect 1726 872 1729 878
rect 1702 842 1705 848
rect 1714 718 1718 721
rect 1694 692 1697 698
rect 1702 662 1705 718
rect 1730 678 1734 681
rect 1486 582 1489 588
rect 1454 572 1457 578
rect 1462 572 1465 578
rect 1510 572 1513 578
rect 1446 542 1449 558
rect 1458 548 1462 551
rect 1298 418 1302 421
rect 1286 392 1289 408
rect 1358 392 1361 468
rect 1370 458 1374 461
rect 1374 392 1377 448
rect 1382 382 1385 478
rect 1390 472 1393 478
rect 1462 472 1465 478
rect 1478 472 1481 538
rect 1486 492 1489 528
rect 1466 468 1470 471
rect 1330 368 1334 371
rect 1370 358 1374 361
rect 1342 352 1345 358
rect 1326 342 1329 348
rect 1278 332 1281 338
rect 1294 302 1297 328
rect 1194 278 1198 281
rect 1158 272 1161 278
rect 1178 268 1182 271
rect 1158 252 1161 258
rect 1146 248 1150 251
rect 1166 222 1169 248
rect 1038 92 1041 118
rect 1046 92 1049 128
rect 1062 122 1065 178
rect 1074 148 1078 151
rect 1086 132 1089 168
rect 1110 162 1113 208
rect 1118 192 1121 218
rect 1174 182 1177 268
rect 1198 242 1201 268
rect 1218 258 1222 261
rect 1234 258 1238 261
rect 1246 252 1249 288
rect 1278 282 1281 298
rect 1302 291 1305 338
rect 1322 328 1326 331
rect 1294 288 1305 291
rect 1258 268 1262 271
rect 1230 242 1233 248
rect 1238 232 1241 238
rect 1226 188 1230 191
rect 1134 172 1137 178
rect 1098 148 1102 151
rect 1126 132 1129 168
rect 1150 162 1153 178
rect 1226 168 1230 171
rect 1158 152 1161 158
rect 1146 148 1153 151
rect 1150 141 1153 148
rect 1166 141 1169 158
rect 1190 152 1193 158
rect 1238 152 1241 178
rect 1246 162 1249 208
rect 1254 192 1257 248
rect 1270 172 1273 248
rect 1286 222 1289 268
rect 1294 232 1297 288
rect 1302 262 1305 268
rect 1322 258 1326 261
rect 1342 252 1345 328
rect 1350 271 1353 318
rect 1358 302 1361 338
rect 1366 332 1369 358
rect 1374 332 1377 348
rect 1366 292 1369 318
rect 1382 292 1385 368
rect 1390 352 1393 468
rect 1406 462 1409 468
rect 1422 462 1425 468
rect 1442 448 1446 451
rect 1414 422 1417 448
rect 1470 442 1473 448
rect 1434 438 1454 441
rect 1426 368 1430 371
rect 1398 362 1401 368
rect 1414 362 1417 368
rect 1446 362 1449 418
rect 1478 402 1481 458
rect 1494 452 1497 558
rect 1510 532 1513 568
rect 1546 558 1550 561
rect 1518 532 1521 538
rect 1510 452 1513 458
rect 1498 448 1502 451
rect 1526 441 1529 518
rect 1542 481 1545 538
rect 1566 532 1569 588
rect 1602 558 1606 561
rect 1614 558 1622 561
rect 1598 532 1601 548
rect 1578 528 1582 531
rect 1538 478 1545 481
rect 1558 481 1561 518
rect 1566 492 1569 528
rect 1558 478 1569 481
rect 1542 472 1545 478
rect 1522 438 1529 441
rect 1534 462 1537 468
rect 1486 422 1489 438
rect 1502 422 1505 438
rect 1486 392 1489 408
rect 1510 402 1513 438
rect 1482 368 1486 371
rect 1490 368 1494 371
rect 1414 342 1417 348
rect 1430 342 1433 348
rect 1398 282 1401 298
rect 1438 292 1441 338
rect 1446 322 1449 358
rect 1454 352 1457 358
rect 1462 352 1465 368
rect 1470 361 1473 368
rect 1510 362 1513 398
rect 1534 392 1537 458
rect 1542 422 1545 468
rect 1558 462 1561 468
rect 1566 441 1569 478
rect 1582 472 1585 478
rect 1598 472 1601 528
rect 1614 492 1617 558
rect 1642 548 1646 551
rect 1630 542 1633 548
rect 1662 532 1665 608
rect 1734 592 1737 628
rect 1702 542 1705 548
rect 1694 532 1697 538
rect 1662 502 1665 528
rect 1578 458 1582 461
rect 1566 438 1574 441
rect 1590 432 1593 448
rect 1566 392 1569 418
rect 1562 368 1566 371
rect 1470 358 1481 361
rect 1374 272 1377 278
rect 1350 268 1361 271
rect 1402 268 1406 271
rect 1350 252 1353 258
rect 1358 252 1361 268
rect 1422 262 1425 268
rect 1442 258 1446 261
rect 1310 182 1313 188
rect 1150 138 1169 141
rect 1174 142 1177 148
rect 1094 92 1097 128
rect 1112 103 1114 107
rect 1118 103 1121 107
rect 1125 103 1128 107
rect 1150 92 1153 128
rect 1030 72 1033 88
rect 1058 78 1062 81
rect 1074 78 1078 81
rect 1102 72 1105 88
rect 1122 68 1126 71
rect 1022 22 1025 68
rect 1038 -18 1041 18
rect 1062 -18 1065 8
rect 1078 -18 1081 18
rect 1102 -18 1105 18
rect 1134 -18 1137 78
rect 1166 62 1169 68
rect 1146 58 1153 61
rect 1142 52 1145 58
rect 1150 -18 1153 58
rect 1174 12 1177 138
rect 1206 132 1209 138
rect 1182 112 1185 128
rect 1190 82 1193 118
rect 1214 112 1217 128
rect 1198 92 1201 108
rect 1238 92 1241 108
rect 1166 -18 1169 8
rect 1022 -19 1026 -18
rect 1014 -22 1026 -19
rect 1038 -22 1042 -18
rect 1062 -22 1066 -18
rect 1078 -22 1082 -18
rect 1102 -22 1106 -18
rect 1134 -22 1138 -18
rect 1150 -22 1154 -18
rect 1166 -22 1170 -18
rect 1190 -19 1193 78
rect 1246 72 1249 118
rect 1262 92 1265 168
rect 1274 158 1278 161
rect 1282 148 1286 151
rect 1270 141 1273 148
rect 1294 141 1297 148
rect 1270 138 1297 141
rect 1302 122 1305 128
rect 1318 92 1321 238
rect 1326 232 1329 248
rect 1334 212 1337 248
rect 1390 242 1393 248
rect 1354 238 1358 241
rect 1406 192 1409 238
rect 1438 172 1441 178
rect 1418 158 1422 161
rect 1342 152 1345 158
rect 1354 138 1358 141
rect 1378 138 1382 141
rect 1326 132 1329 138
rect 1286 82 1289 88
rect 1326 82 1329 128
rect 1334 122 1337 128
rect 1366 122 1369 128
rect 1366 92 1369 108
rect 1374 102 1377 128
rect 1382 92 1385 98
rect 1390 92 1393 158
rect 1410 138 1414 141
rect 1226 68 1230 71
rect 1222 12 1225 58
rect 1278 52 1281 78
rect 1290 58 1294 61
rect 1238 42 1241 48
rect 1198 -19 1202 -18
rect 1190 -22 1202 -19
rect 1214 -19 1217 8
rect 1238 -18 1241 8
rect 1262 -18 1265 38
rect 1278 -18 1281 48
rect 1302 32 1305 78
rect 1334 72 1337 88
rect 1342 72 1345 78
rect 1382 72 1385 88
rect 1398 72 1401 98
rect 1414 92 1417 108
rect 1422 102 1425 148
rect 1438 122 1441 148
rect 1422 72 1425 98
rect 1446 92 1449 238
rect 1462 201 1465 328
rect 1478 322 1481 358
rect 1514 348 1518 351
rect 1502 322 1505 348
rect 1526 342 1529 358
rect 1542 342 1545 348
rect 1470 292 1473 318
rect 1494 292 1497 318
rect 1518 292 1521 318
rect 1486 262 1489 268
rect 1526 262 1529 338
rect 1550 292 1553 368
rect 1586 348 1590 351
rect 1566 282 1569 288
rect 1538 268 1542 271
rect 1510 252 1513 258
rect 1518 252 1521 258
rect 1470 212 1473 218
rect 1462 198 1473 201
rect 1470 192 1473 198
rect 1478 172 1481 248
rect 1502 242 1505 248
rect 1530 238 1534 241
rect 1494 162 1497 208
rect 1502 152 1505 158
rect 1490 148 1494 151
rect 1510 141 1513 168
rect 1502 138 1513 141
rect 1518 142 1521 188
rect 1542 162 1545 268
rect 1582 262 1585 348
rect 1590 302 1593 318
rect 1598 282 1601 468
rect 1630 462 1633 468
rect 1678 462 1681 518
rect 1694 482 1697 528
rect 1702 472 1705 518
rect 1710 482 1713 488
rect 1610 448 1614 451
rect 1614 402 1617 418
rect 1614 362 1617 398
rect 1622 372 1625 448
rect 1638 442 1641 448
rect 1654 442 1657 448
rect 1662 442 1665 458
rect 1670 452 1673 458
rect 1686 452 1689 458
rect 1678 442 1681 448
rect 1630 392 1633 418
rect 1638 392 1641 408
rect 1622 362 1625 368
rect 1630 362 1633 368
rect 1646 362 1649 428
rect 1654 392 1657 398
rect 1678 382 1681 438
rect 1702 372 1705 448
rect 1662 362 1665 368
rect 1706 358 1710 361
rect 1610 348 1614 351
rect 1626 348 1630 351
rect 1614 272 1617 338
rect 1558 202 1561 248
rect 1582 192 1585 258
rect 1590 192 1593 238
rect 1614 221 1617 268
rect 1626 258 1630 261
rect 1606 218 1617 221
rect 1594 168 1598 171
rect 1530 158 1534 161
rect 1578 158 1582 161
rect 1538 148 1542 151
rect 1586 148 1590 151
rect 1458 128 1462 131
rect 1478 92 1481 138
rect 1502 92 1505 138
rect 1526 102 1529 128
rect 1542 92 1545 108
rect 1550 102 1553 148
rect 1566 122 1569 128
rect 1574 92 1577 148
rect 1598 142 1601 158
rect 1354 68 1358 71
rect 1358 52 1361 58
rect 1406 52 1409 58
rect 1430 52 1433 78
rect 1462 72 1465 88
rect 1486 72 1489 88
rect 1518 82 1521 88
rect 1550 82 1553 88
rect 1578 78 1582 81
rect 1526 72 1529 78
rect 1590 72 1593 118
rect 1606 92 1609 218
rect 1614 162 1617 208
rect 1622 192 1625 248
rect 1646 212 1649 358
rect 1658 348 1662 351
rect 1678 332 1681 338
rect 1682 288 1686 291
rect 1682 278 1686 281
rect 1694 272 1697 308
rect 1710 282 1713 338
rect 1718 292 1721 348
rect 1630 152 1633 168
rect 1642 158 1646 161
rect 1654 152 1657 198
rect 1710 152 1713 188
rect 1622 112 1625 148
rect 1662 142 1665 148
rect 1662 92 1665 138
rect 1686 132 1689 148
rect 1694 132 1697 138
rect 1682 128 1686 131
rect 1670 92 1673 98
rect 1718 92 1721 258
rect 1662 72 1665 78
rect 1690 68 1694 71
rect 1494 52 1497 68
rect 1470 42 1473 48
rect 1374 32 1377 38
rect 1326 -18 1329 8
rect 1526 -18 1529 68
rect 1558 22 1561 68
rect 1706 66 1710 69
rect 1734 62 1737 148
rect 1690 58 1694 61
rect 1558 -18 1561 18
rect 1222 -19 1226 -18
rect 1214 -22 1226 -19
rect 1238 -22 1242 -18
rect 1262 -22 1266 -18
rect 1278 -22 1282 -18
rect 1326 -22 1330 -18
rect 1526 -22 1530 -18
rect 1558 -22 1562 -18
<< m3contact >>
rect 62 1588 66 1592
rect 118 1588 122 1592
rect 158 1558 162 1562
rect 190 1548 194 1552
rect 278 1608 282 1612
rect 206 1568 210 1572
rect 246 1568 250 1572
rect 94 1538 98 1542
rect 126 1538 130 1542
rect 166 1538 170 1542
rect 182 1538 186 1542
rect 222 1538 226 1542
rect 6 1518 10 1522
rect 38 1468 42 1472
rect 6 1458 10 1462
rect 6 1448 10 1452
rect 86 1528 90 1532
rect 110 1528 114 1532
rect 62 1488 66 1492
rect 54 1478 58 1482
rect 118 1478 122 1482
rect 30 1458 34 1462
rect 46 1458 50 1462
rect 70 1468 74 1472
rect 254 1538 258 1542
rect 286 1538 290 1542
rect 182 1518 186 1522
rect 62 1458 66 1462
rect 78 1458 82 1462
rect 134 1458 138 1462
rect 142 1458 146 1462
rect 54 1428 58 1432
rect 30 1408 34 1412
rect 22 1398 26 1402
rect 38 1398 42 1402
rect 22 1388 26 1392
rect 54 1378 58 1382
rect 118 1448 122 1452
rect 198 1488 202 1492
rect 190 1478 194 1482
rect 158 1468 162 1472
rect 174 1468 178 1472
rect 182 1468 186 1472
rect 70 1438 74 1442
rect 86 1408 90 1412
rect 46 1368 50 1372
rect 134 1378 138 1382
rect 110 1368 114 1372
rect 118 1368 122 1372
rect 126 1368 130 1372
rect 46 1348 50 1352
rect 54 1348 58 1352
rect 78 1328 82 1332
rect 22 1318 26 1322
rect 14 1298 18 1302
rect 14 1258 18 1262
rect 6 1248 10 1252
rect 6 1228 10 1232
rect 14 1208 18 1212
rect 118 1348 122 1352
rect 94 1338 98 1342
rect 86 1298 90 1302
rect 78 1268 82 1272
rect 102 1278 106 1282
rect 54 1248 58 1252
rect 22 1198 26 1202
rect 6 1148 10 1152
rect 14 1128 18 1132
rect 22 1128 26 1132
rect 38 1128 42 1132
rect 6 1098 10 1102
rect 14 1088 18 1092
rect 14 1058 18 1062
rect 14 1048 18 1052
rect 38 1058 42 1062
rect 30 1028 34 1032
rect 6 978 10 982
rect 6 948 10 952
rect 30 918 34 922
rect 6 898 10 902
rect 22 878 26 882
rect 38 858 42 862
rect 30 848 34 852
rect 38 798 42 802
rect 22 728 26 732
rect 6 648 10 652
rect 54 1188 58 1192
rect 70 1158 74 1162
rect 70 1138 74 1142
rect 150 1358 154 1362
rect 158 1358 162 1362
rect 214 1468 218 1472
rect 206 1448 210 1452
rect 358 1588 362 1592
rect 366 1558 370 1562
rect 374 1558 378 1562
rect 398 1548 402 1552
rect 318 1538 322 1542
rect 350 1538 354 1542
rect 382 1538 386 1542
rect 286 1528 290 1532
rect 310 1528 314 1532
rect 334 1528 338 1532
rect 246 1478 250 1482
rect 246 1468 250 1472
rect 262 1458 266 1462
rect 302 1508 306 1512
rect 302 1478 306 1482
rect 358 1488 362 1492
rect 318 1468 322 1472
rect 350 1468 354 1472
rect 278 1458 282 1462
rect 382 1458 386 1462
rect 310 1448 314 1452
rect 254 1438 258 1442
rect 198 1408 202 1412
rect 230 1388 234 1392
rect 214 1368 218 1372
rect 182 1348 186 1352
rect 206 1328 210 1332
rect 158 1318 162 1322
rect 110 1248 114 1252
rect 86 1238 90 1242
rect 182 1308 186 1312
rect 174 1258 178 1262
rect 166 1238 170 1242
rect 134 1218 138 1222
rect 174 1218 178 1222
rect 110 1178 114 1182
rect 110 1168 114 1172
rect 118 1168 122 1172
rect 126 1158 130 1162
rect 142 1158 146 1162
rect 214 1318 218 1322
rect 406 1528 410 1532
rect 446 1608 450 1612
rect 534 1578 538 1582
rect 422 1558 426 1562
rect 542 1558 546 1562
rect 518 1548 522 1552
rect 558 1548 562 1552
rect 422 1538 426 1542
rect 446 1538 450 1542
rect 494 1538 498 1542
rect 422 1508 426 1512
rect 398 1458 402 1462
rect 294 1428 298 1432
rect 334 1428 338 1432
rect 286 1388 290 1392
rect 262 1368 266 1372
rect 286 1358 290 1362
rect 374 1398 378 1402
rect 302 1358 306 1362
rect 326 1358 330 1362
rect 334 1358 338 1362
rect 382 1358 386 1362
rect 406 1368 410 1372
rect 294 1348 298 1352
rect 398 1348 402 1352
rect 326 1338 330 1342
rect 254 1318 258 1322
rect 230 1308 234 1312
rect 230 1288 234 1292
rect 222 1278 226 1282
rect 206 1268 210 1272
rect 214 1268 218 1272
rect 214 1248 218 1252
rect 198 1238 202 1242
rect 206 1228 210 1232
rect 198 1188 202 1192
rect 166 1148 170 1152
rect 110 1118 114 1122
rect 134 1118 138 1122
rect 174 1118 178 1122
rect 62 1098 66 1102
rect 78 1098 82 1102
rect 102 1098 106 1102
rect 54 1058 58 1062
rect 54 1038 58 1042
rect 70 1038 74 1042
rect 62 1018 66 1022
rect 54 958 58 962
rect 94 1068 98 1072
rect 110 1068 114 1072
rect 158 1068 162 1072
rect 118 1058 122 1062
rect 86 1048 90 1052
rect 94 1038 98 1042
rect 150 1058 154 1062
rect 142 1038 146 1042
rect 166 1038 170 1042
rect 126 998 130 1002
rect 102 968 106 972
rect 134 958 138 962
rect 214 1128 218 1132
rect 198 1118 202 1122
rect 278 1328 282 1332
rect 302 1328 306 1332
rect 358 1328 362 1332
rect 390 1328 394 1332
rect 270 1278 274 1282
rect 270 1268 274 1272
rect 262 1218 266 1222
rect 238 1118 242 1122
rect 206 1088 210 1092
rect 222 1078 226 1082
rect 214 1068 218 1072
rect 222 1058 226 1062
rect 190 1028 194 1032
rect 254 1108 258 1112
rect 246 1068 250 1072
rect 326 1318 330 1322
rect 390 1318 394 1322
rect 406 1318 410 1322
rect 286 1268 290 1272
rect 294 1268 298 1272
rect 286 1258 290 1262
rect 294 1238 298 1242
rect 326 1268 330 1272
rect 334 1248 338 1252
rect 302 1218 306 1222
rect 318 1208 322 1212
rect 302 1168 306 1172
rect 318 1168 322 1172
rect 270 1108 274 1112
rect 310 1138 314 1142
rect 310 1118 314 1122
rect 278 1088 282 1092
rect 278 1058 282 1062
rect 238 1028 242 1032
rect 174 968 178 972
rect 206 968 210 972
rect 230 968 234 972
rect 358 1228 362 1232
rect 342 1218 346 1222
rect 334 1188 338 1192
rect 334 1168 338 1172
rect 326 1148 330 1152
rect 326 1138 330 1142
rect 406 1308 410 1312
rect 398 1278 402 1282
rect 382 1248 386 1252
rect 390 1248 394 1252
rect 382 1238 386 1242
rect 510 1528 514 1532
rect 462 1518 466 1522
rect 454 1508 458 1512
rect 446 1478 450 1482
rect 438 1448 442 1452
rect 446 1428 450 1432
rect 446 1368 450 1372
rect 438 1348 442 1352
rect 430 1318 434 1322
rect 518 1518 522 1522
rect 526 1518 530 1522
rect 502 1508 506 1512
rect 486 1488 490 1492
rect 502 1488 506 1492
rect 462 1478 466 1482
rect 462 1458 466 1462
rect 502 1458 506 1462
rect 534 1468 538 1472
rect 526 1458 530 1462
rect 478 1388 482 1392
rect 510 1388 514 1392
rect 502 1368 506 1372
rect 494 1358 498 1362
rect 470 1348 474 1352
rect 502 1348 506 1352
rect 454 1328 458 1332
rect 630 1608 634 1612
rect 602 1603 606 1607
rect 609 1603 613 1607
rect 694 1608 698 1612
rect 678 1588 682 1592
rect 710 1588 714 1592
rect 630 1578 634 1582
rect 646 1578 650 1582
rect 670 1578 674 1582
rect 622 1558 626 1562
rect 582 1548 586 1552
rect 606 1548 610 1552
rect 574 1508 578 1512
rect 550 1498 554 1502
rect 566 1498 570 1502
rect 558 1448 562 1452
rect 646 1548 650 1552
rect 582 1468 586 1472
rect 646 1468 650 1472
rect 654 1468 658 1472
rect 590 1458 594 1462
rect 646 1448 650 1452
rect 670 1478 674 1482
rect 686 1568 690 1572
rect 726 1568 730 1572
rect 702 1558 706 1562
rect 718 1548 722 1552
rect 758 1558 762 1562
rect 702 1538 706 1542
rect 750 1538 754 1542
rect 686 1478 690 1482
rect 686 1468 690 1472
rect 678 1458 682 1462
rect 686 1448 690 1452
rect 702 1478 706 1482
rect 622 1438 626 1442
rect 646 1438 650 1442
rect 1230 1608 1234 1612
rect 902 1568 906 1572
rect 1398 1568 1402 1572
rect 1478 1568 1482 1572
rect 1510 1568 1514 1572
rect 1590 1568 1594 1572
rect 790 1558 794 1562
rect 974 1558 978 1562
rect 998 1558 1002 1562
rect 1006 1558 1010 1562
rect 1070 1558 1074 1562
rect 1158 1558 1162 1562
rect 1166 1558 1170 1562
rect 1294 1558 1298 1562
rect 1430 1558 1434 1562
rect 774 1548 778 1552
rect 806 1548 810 1552
rect 934 1548 938 1552
rect 806 1538 810 1542
rect 854 1538 858 1542
rect 742 1528 746 1532
rect 766 1528 770 1532
rect 734 1488 738 1492
rect 766 1488 770 1492
rect 774 1488 778 1492
rect 726 1478 730 1482
rect 742 1468 746 1472
rect 758 1468 762 1472
rect 750 1458 754 1462
rect 758 1448 762 1452
rect 550 1368 554 1372
rect 574 1398 578 1402
rect 566 1378 570 1382
rect 602 1403 606 1407
rect 609 1403 613 1407
rect 582 1378 586 1382
rect 678 1368 682 1372
rect 614 1358 618 1362
rect 542 1348 546 1352
rect 558 1348 562 1352
rect 574 1348 578 1352
rect 654 1348 658 1352
rect 702 1348 706 1352
rect 526 1338 530 1342
rect 550 1338 554 1342
rect 566 1338 570 1342
rect 606 1338 610 1342
rect 646 1338 650 1342
rect 694 1338 698 1342
rect 566 1328 570 1332
rect 638 1328 642 1332
rect 510 1288 514 1292
rect 462 1268 466 1272
rect 526 1268 530 1272
rect 430 1238 434 1242
rect 422 1218 426 1222
rect 414 1208 418 1212
rect 374 1168 378 1172
rect 390 1168 394 1172
rect 478 1258 482 1262
rect 502 1248 506 1252
rect 470 1238 474 1242
rect 542 1258 546 1262
rect 566 1248 570 1252
rect 550 1228 554 1232
rect 646 1278 650 1282
rect 662 1278 666 1282
rect 686 1278 690 1282
rect 630 1258 634 1262
rect 662 1258 666 1262
rect 686 1258 690 1262
rect 590 1238 594 1242
rect 606 1238 610 1242
rect 622 1228 626 1232
rect 582 1218 586 1222
rect 602 1203 606 1207
rect 609 1203 613 1207
rect 526 1188 530 1192
rect 558 1188 562 1192
rect 454 1168 458 1172
rect 486 1168 490 1172
rect 574 1178 578 1182
rect 430 1158 434 1162
rect 446 1158 450 1162
rect 486 1158 490 1162
rect 382 1148 386 1152
rect 406 1148 410 1152
rect 342 1108 346 1112
rect 334 1078 338 1082
rect 310 1058 314 1062
rect 262 1038 266 1042
rect 278 1038 282 1042
rect 294 978 298 982
rect 286 968 290 972
rect 358 1058 362 1062
rect 358 1048 362 1052
rect 374 1048 378 1052
rect 366 988 370 992
rect 302 968 306 972
rect 350 968 354 972
rect 358 968 362 972
rect 254 958 258 962
rect 270 958 274 962
rect 78 948 82 952
rect 134 948 138 952
rect 158 948 162 952
rect 118 938 122 942
rect 174 948 178 952
rect 246 948 250 952
rect 94 928 98 932
rect 62 888 66 892
rect 54 868 58 872
rect 158 928 162 932
rect 142 908 146 912
rect 118 888 122 892
rect 222 938 226 942
rect 254 938 258 942
rect 190 918 194 922
rect 190 898 194 902
rect 238 888 242 892
rect 86 878 90 882
rect 118 878 122 882
rect 150 878 154 882
rect 174 878 178 882
rect 190 878 194 882
rect 230 878 234 882
rect 110 868 114 872
rect 94 838 98 842
rect 110 838 114 842
rect 134 858 138 862
rect 118 828 122 832
rect 102 818 106 822
rect 70 808 74 812
rect 70 798 74 802
rect 110 778 114 782
rect 46 768 50 772
rect 46 758 50 762
rect 54 748 58 752
rect 78 748 82 752
rect 134 818 138 822
rect 142 748 146 752
rect 134 738 138 742
rect 46 728 50 732
rect 102 728 106 732
rect 110 728 114 732
rect 46 718 50 722
rect 54 708 58 712
rect 62 698 66 702
rect 198 868 202 872
rect 222 868 226 872
rect 174 848 178 852
rect 182 848 186 852
rect 158 838 162 842
rect 310 948 314 952
rect 286 938 290 942
rect 326 958 330 962
rect 470 1138 474 1142
rect 502 1138 506 1142
rect 446 1128 450 1132
rect 510 1128 514 1132
rect 518 1128 522 1132
rect 390 1118 394 1122
rect 414 1118 418 1122
rect 390 1058 394 1062
rect 398 1048 402 1052
rect 398 1008 402 1012
rect 414 998 418 1002
rect 414 978 418 982
rect 486 1118 490 1122
rect 518 1118 522 1122
rect 550 1118 554 1122
rect 470 1098 474 1102
rect 438 1068 442 1072
rect 510 1088 514 1092
rect 494 1058 498 1062
rect 614 1148 618 1152
rect 566 1138 570 1142
rect 590 1128 594 1132
rect 558 1088 562 1092
rect 542 1068 546 1072
rect 574 1068 578 1072
rect 678 1248 682 1252
rect 734 1358 738 1362
rect 750 1358 754 1362
rect 702 1328 706 1332
rect 750 1328 754 1332
rect 702 1278 706 1282
rect 710 1268 714 1272
rect 734 1278 738 1282
rect 798 1488 802 1492
rect 790 1478 794 1482
rect 790 1468 794 1472
rect 782 1438 786 1442
rect 790 1418 794 1422
rect 774 1338 778 1342
rect 766 1308 770 1312
rect 734 1258 738 1262
rect 822 1478 826 1482
rect 942 1538 946 1542
rect 966 1538 970 1542
rect 870 1528 874 1532
rect 870 1508 874 1512
rect 862 1478 866 1482
rect 854 1468 858 1472
rect 846 1458 850 1462
rect 814 1368 818 1372
rect 878 1498 882 1502
rect 862 1458 866 1462
rect 910 1528 914 1532
rect 934 1518 938 1522
rect 910 1498 914 1502
rect 910 1488 914 1492
rect 998 1528 1002 1532
rect 1094 1548 1098 1552
rect 1166 1548 1170 1552
rect 1238 1548 1242 1552
rect 1294 1548 1298 1552
rect 1310 1548 1314 1552
rect 1326 1548 1330 1552
rect 1118 1538 1122 1542
rect 1142 1538 1146 1542
rect 1150 1538 1154 1542
rect 1182 1538 1186 1542
rect 982 1518 986 1522
rect 1006 1518 1010 1522
rect 958 1508 962 1512
rect 990 1508 994 1512
rect 894 1478 898 1482
rect 950 1478 954 1482
rect 958 1478 962 1482
rect 966 1478 970 1482
rect 902 1468 906 1472
rect 926 1468 930 1472
rect 926 1458 930 1462
rect 934 1458 938 1462
rect 950 1458 954 1462
rect 894 1448 898 1452
rect 910 1418 914 1422
rect 886 1408 890 1412
rect 942 1448 946 1452
rect 942 1438 946 1442
rect 958 1378 962 1382
rect 926 1368 930 1372
rect 942 1368 946 1372
rect 854 1358 858 1362
rect 838 1348 842 1352
rect 846 1338 850 1342
rect 782 1308 786 1312
rect 726 1248 730 1252
rect 710 1238 714 1242
rect 718 1228 722 1232
rect 694 1178 698 1182
rect 702 1178 706 1182
rect 718 1178 722 1182
rect 630 1158 634 1162
rect 686 1158 690 1162
rect 710 1148 714 1152
rect 670 1108 674 1112
rect 646 1098 650 1102
rect 670 1088 674 1092
rect 702 1088 706 1092
rect 622 1078 626 1082
rect 622 1068 626 1072
rect 550 1058 554 1062
rect 574 1058 578 1062
rect 526 1048 530 1052
rect 478 1038 482 1042
rect 486 1038 490 1042
rect 502 1028 506 1032
rect 454 1018 458 1022
rect 478 998 482 1002
rect 422 968 426 972
rect 406 958 410 962
rect 366 948 370 952
rect 334 938 338 942
rect 374 938 378 942
rect 342 928 346 932
rect 262 878 266 882
rect 310 878 314 882
rect 342 878 346 882
rect 358 878 362 882
rect 366 878 370 882
rect 382 878 386 882
rect 262 868 266 872
rect 254 858 258 862
rect 278 858 282 862
rect 302 858 306 862
rect 318 858 322 862
rect 342 858 346 862
rect 310 848 314 852
rect 158 818 162 822
rect 206 818 210 822
rect 206 778 210 782
rect 254 768 258 772
rect 158 758 162 762
rect 166 748 170 752
rect 150 718 154 722
rect 102 708 106 712
rect 78 678 82 682
rect 110 678 114 682
rect 86 668 90 672
rect 94 668 98 672
rect 102 668 106 672
rect 38 658 42 662
rect 38 648 42 652
rect 94 648 98 652
rect 6 628 10 632
rect 30 618 34 622
rect 38 618 42 622
rect 62 578 66 582
rect 86 578 90 582
rect 38 568 42 572
rect 54 568 58 572
rect 134 678 138 682
rect 126 668 130 672
rect 126 658 130 662
rect 174 738 178 742
rect 230 738 234 742
rect 214 728 218 732
rect 158 658 162 662
rect 174 658 178 662
rect 118 608 122 612
rect 30 548 34 552
rect 22 538 26 542
rect 54 538 58 542
rect 54 508 58 512
rect 86 528 90 532
rect 70 498 74 502
rect 94 498 98 502
rect 78 488 82 492
rect 70 478 74 482
rect 38 468 42 472
rect 6 458 10 462
rect 22 458 26 462
rect 30 438 34 442
rect 78 438 82 442
rect 46 418 50 422
rect 134 608 138 612
rect 134 598 138 602
rect 158 578 162 582
rect 150 568 154 572
rect 174 578 178 582
rect 166 568 170 572
rect 326 798 330 802
rect 326 758 330 762
rect 294 748 298 752
rect 374 868 378 872
rect 462 968 466 972
rect 526 968 530 972
rect 574 1038 578 1042
rect 582 1038 586 1042
rect 734 1158 738 1162
rect 814 1328 818 1332
rect 814 1308 818 1312
rect 886 1348 890 1352
rect 782 1138 786 1142
rect 942 1358 946 1362
rect 998 1468 1002 1472
rect 974 1458 978 1462
rect 990 1458 994 1462
rect 966 1368 970 1372
rect 974 1358 978 1362
rect 902 1338 906 1342
rect 918 1338 922 1342
rect 942 1338 946 1342
rect 974 1338 978 1342
rect 878 1328 882 1332
rect 838 1248 842 1252
rect 862 1248 866 1252
rect 806 1188 810 1192
rect 1094 1528 1098 1532
rect 1046 1518 1050 1522
rect 1062 1518 1066 1522
rect 1014 1508 1018 1512
rect 1022 1488 1026 1492
rect 1114 1503 1118 1507
rect 1121 1503 1125 1507
rect 1030 1478 1034 1482
rect 1102 1478 1106 1482
rect 1094 1468 1098 1472
rect 1126 1468 1130 1472
rect 1014 1458 1018 1462
rect 1174 1498 1178 1502
rect 1198 1498 1202 1502
rect 1166 1478 1170 1482
rect 1142 1468 1146 1472
rect 1158 1468 1162 1472
rect 1062 1458 1066 1462
rect 1070 1458 1074 1462
rect 1110 1458 1114 1462
rect 1150 1458 1154 1462
rect 1070 1448 1074 1452
rect 1014 1428 1018 1432
rect 1006 1418 1010 1422
rect 1030 1418 1034 1422
rect 998 1398 1002 1402
rect 990 1388 994 1392
rect 998 1378 1002 1382
rect 990 1358 994 1362
rect 1014 1398 1018 1402
rect 990 1328 994 1332
rect 982 1318 986 1322
rect 958 1278 962 1282
rect 910 1259 914 1263
rect 1022 1388 1026 1392
rect 1094 1438 1098 1442
rect 1062 1428 1066 1432
rect 1078 1428 1082 1432
rect 1054 1408 1058 1412
rect 1022 1338 1026 1342
rect 1030 1338 1034 1342
rect 1038 1298 1042 1302
rect 1014 1288 1018 1292
rect 1006 1278 1010 1282
rect 1038 1278 1042 1282
rect 1046 1268 1050 1272
rect 990 1258 994 1262
rect 958 1248 962 1252
rect 982 1248 986 1252
rect 1022 1248 1026 1252
rect 1046 1228 1050 1232
rect 918 1188 922 1192
rect 950 1188 954 1192
rect 806 1168 810 1172
rect 902 1168 906 1172
rect 870 1158 874 1162
rect 838 1138 842 1142
rect 798 1118 802 1122
rect 814 1098 818 1102
rect 710 1068 714 1072
rect 766 1068 770 1072
rect 630 1058 634 1062
rect 646 1058 650 1062
rect 678 1058 682 1062
rect 638 1048 642 1052
rect 686 1048 690 1052
rect 662 1028 666 1032
rect 670 1028 674 1032
rect 630 1018 634 1022
rect 602 1003 606 1007
rect 609 1003 613 1007
rect 574 968 578 972
rect 606 968 610 972
rect 454 958 458 962
rect 478 958 482 962
rect 558 958 562 962
rect 438 948 442 952
rect 470 948 474 952
rect 566 948 570 952
rect 518 938 522 942
rect 558 938 562 942
rect 526 928 530 932
rect 414 868 418 872
rect 390 848 394 852
rect 414 848 418 852
rect 366 828 370 832
rect 374 818 378 822
rect 398 818 402 822
rect 390 808 394 812
rect 398 798 402 802
rect 422 808 426 812
rect 414 768 418 772
rect 358 748 362 752
rect 270 728 274 732
rect 318 728 322 732
rect 334 728 338 732
rect 350 728 354 732
rect 214 678 218 682
rect 230 678 234 682
rect 198 668 202 672
rect 278 718 282 722
rect 254 708 258 712
rect 302 708 306 712
rect 262 678 266 682
rect 278 678 282 682
rect 366 718 370 722
rect 358 688 362 692
rect 294 668 298 672
rect 302 658 306 662
rect 262 648 266 652
rect 294 648 298 652
rect 318 648 322 652
rect 342 658 346 662
rect 382 648 386 652
rect 470 898 474 902
rect 494 898 498 902
rect 438 878 442 882
rect 486 878 490 882
rect 518 878 522 882
rect 446 848 450 852
rect 486 848 490 852
rect 494 848 498 852
rect 510 848 514 852
rect 470 838 474 842
rect 494 838 498 842
rect 502 818 506 822
rect 438 798 442 802
rect 462 798 466 802
rect 446 768 450 772
rect 486 768 490 772
rect 518 828 522 832
rect 430 758 434 762
rect 454 758 458 762
rect 478 758 482 762
rect 494 748 498 752
rect 534 868 538 872
rect 678 978 682 982
rect 662 958 666 962
rect 622 918 626 922
rect 710 1018 714 1022
rect 758 1058 762 1062
rect 694 968 698 972
rect 718 968 722 972
rect 710 958 714 962
rect 702 938 706 942
rect 718 938 722 942
rect 702 928 706 932
rect 582 878 586 882
rect 662 878 666 882
rect 710 918 714 922
rect 582 868 586 872
rect 550 858 554 862
rect 622 858 626 862
rect 574 848 578 852
rect 558 838 562 842
rect 630 838 634 842
rect 678 838 682 842
rect 542 828 546 832
rect 638 828 642 832
rect 654 828 658 832
rect 602 803 606 807
rect 609 803 613 807
rect 598 788 602 792
rect 646 788 650 792
rect 558 768 562 772
rect 638 768 642 772
rect 646 768 650 772
rect 550 758 554 762
rect 542 748 546 752
rect 574 748 578 752
rect 462 728 466 732
rect 486 728 490 732
rect 526 728 530 732
rect 462 708 466 712
rect 422 688 426 692
rect 494 688 498 692
rect 422 668 426 672
rect 446 668 450 672
rect 502 668 506 672
rect 590 758 594 762
rect 614 758 618 762
rect 550 718 554 722
rect 590 728 594 732
rect 670 818 674 822
rect 686 818 690 822
rect 694 818 698 822
rect 702 788 706 792
rect 678 768 682 772
rect 662 748 666 752
rect 630 728 634 732
rect 646 728 650 732
rect 622 688 626 692
rect 694 738 698 742
rect 686 728 690 732
rect 670 678 674 682
rect 726 908 730 912
rect 726 868 730 872
rect 718 858 722 862
rect 774 1038 778 1042
rect 806 1048 810 1052
rect 822 1068 826 1072
rect 894 1068 898 1072
rect 838 1058 842 1062
rect 870 1058 874 1062
rect 822 1048 826 1052
rect 846 1038 850 1042
rect 790 1028 794 1032
rect 854 1028 858 1032
rect 742 978 746 982
rect 822 1008 826 1012
rect 790 998 794 1002
rect 846 988 850 992
rect 854 978 858 982
rect 814 968 818 972
rect 838 968 842 972
rect 750 958 754 962
rect 806 958 810 962
rect 838 958 842 962
rect 878 1028 882 1032
rect 886 998 890 1002
rect 870 988 874 992
rect 878 958 882 962
rect 742 948 746 952
rect 798 948 802 952
rect 814 948 818 952
rect 862 948 866 952
rect 758 928 762 932
rect 838 928 842 932
rect 862 928 866 932
rect 774 918 778 922
rect 806 908 810 912
rect 798 898 802 902
rect 774 888 778 892
rect 750 878 754 882
rect 758 868 762 872
rect 742 858 746 862
rect 766 858 770 862
rect 734 848 738 852
rect 726 838 730 842
rect 718 828 722 832
rect 750 798 754 802
rect 734 788 738 792
rect 758 778 762 782
rect 726 768 730 772
rect 742 758 746 762
rect 734 748 738 752
rect 750 748 754 752
rect 782 858 786 862
rect 790 848 794 852
rect 782 828 786 832
rect 862 918 866 922
rect 878 918 882 922
rect 926 1148 930 1152
rect 1094 1348 1098 1352
rect 1134 1448 1138 1452
rect 1126 1438 1130 1442
rect 1230 1538 1234 1542
rect 1222 1528 1226 1532
rect 1222 1518 1226 1522
rect 1214 1478 1218 1482
rect 1206 1468 1210 1472
rect 1254 1528 1258 1532
rect 1302 1528 1306 1532
rect 1318 1528 1322 1532
rect 1326 1528 1330 1532
rect 1238 1518 1242 1522
rect 1270 1508 1274 1512
rect 1238 1488 1242 1492
rect 1158 1448 1162 1452
rect 1182 1448 1186 1452
rect 1134 1398 1138 1402
rect 1086 1338 1090 1342
rect 1110 1338 1114 1342
rect 1078 1328 1082 1332
rect 1114 1303 1118 1307
rect 1121 1303 1125 1307
rect 1118 1278 1122 1282
rect 1102 1268 1106 1272
rect 1206 1438 1210 1442
rect 1342 1518 1346 1522
rect 1286 1478 1290 1482
rect 1254 1468 1258 1472
rect 1254 1458 1258 1462
rect 1270 1458 1274 1462
rect 1222 1418 1226 1422
rect 1286 1418 1290 1422
rect 1286 1408 1290 1412
rect 1278 1388 1282 1392
rect 1326 1458 1330 1462
rect 1318 1438 1322 1442
rect 1326 1418 1330 1422
rect 1302 1398 1306 1402
rect 1382 1548 1386 1552
rect 1414 1548 1418 1552
rect 1374 1518 1378 1522
rect 1374 1508 1378 1512
rect 1366 1488 1370 1492
rect 1358 1448 1362 1452
rect 1390 1538 1394 1542
rect 1422 1538 1426 1542
rect 1438 1528 1442 1532
rect 1446 1518 1450 1522
rect 1550 1558 1554 1562
rect 1470 1548 1474 1552
rect 1478 1548 1482 1552
rect 1494 1548 1498 1552
rect 1518 1548 1522 1552
rect 1470 1528 1474 1532
rect 1486 1508 1490 1512
rect 1462 1498 1466 1502
rect 1510 1538 1514 1542
rect 1526 1528 1530 1532
rect 1598 1548 1602 1552
rect 1550 1538 1554 1542
rect 1550 1528 1554 1532
rect 1534 1518 1538 1522
rect 1542 1508 1546 1512
rect 1422 1468 1426 1472
rect 1446 1468 1450 1472
rect 1462 1468 1466 1472
rect 1398 1458 1402 1462
rect 1430 1448 1434 1452
rect 1406 1438 1410 1442
rect 1422 1428 1426 1432
rect 1390 1418 1394 1422
rect 1382 1408 1386 1412
rect 1438 1408 1442 1412
rect 1366 1398 1370 1402
rect 1494 1418 1498 1422
rect 1478 1398 1482 1402
rect 1350 1388 1354 1392
rect 1390 1388 1394 1392
rect 1294 1378 1298 1382
rect 1270 1368 1274 1372
rect 1374 1368 1378 1372
rect 1310 1358 1314 1362
rect 1414 1358 1418 1362
rect 1150 1348 1154 1352
rect 1166 1348 1170 1352
rect 1206 1348 1210 1352
rect 1158 1328 1162 1332
rect 1174 1328 1178 1332
rect 1182 1328 1186 1332
rect 1222 1328 1226 1332
rect 1166 1318 1170 1322
rect 1158 1298 1162 1302
rect 1198 1318 1202 1322
rect 1246 1348 1250 1352
rect 1334 1348 1338 1352
rect 1438 1348 1442 1352
rect 1270 1318 1274 1322
rect 1246 1308 1250 1312
rect 1238 1298 1242 1302
rect 1182 1288 1186 1292
rect 1150 1238 1154 1242
rect 1142 1218 1146 1222
rect 1166 1148 1170 1152
rect 974 1108 978 1112
rect 910 1058 914 1062
rect 926 1048 930 1052
rect 926 1038 930 1042
rect 1030 1108 1034 1112
rect 1114 1103 1118 1107
rect 1121 1103 1125 1107
rect 1046 1088 1050 1092
rect 1118 1088 1122 1092
rect 1022 1078 1026 1082
rect 1278 1298 1282 1302
rect 1278 1278 1282 1282
rect 1198 1258 1202 1262
rect 1214 1258 1218 1262
rect 1230 1258 1234 1262
rect 1214 1248 1218 1252
rect 1238 1248 1242 1252
rect 1206 1238 1210 1242
rect 1262 1228 1266 1232
rect 1302 1338 1306 1342
rect 1294 1308 1298 1312
rect 1310 1328 1314 1332
rect 1310 1308 1314 1312
rect 1294 1278 1298 1282
rect 1318 1278 1322 1282
rect 1334 1328 1338 1332
rect 1374 1338 1378 1342
rect 1406 1338 1410 1342
rect 1438 1338 1442 1342
rect 1342 1318 1346 1322
rect 1422 1318 1426 1322
rect 1430 1298 1434 1302
rect 1382 1288 1386 1292
rect 1414 1288 1418 1292
rect 1366 1278 1370 1282
rect 1310 1258 1314 1262
rect 1350 1258 1354 1262
rect 1358 1258 1362 1262
rect 1342 1228 1346 1232
rect 1222 1218 1226 1222
rect 1246 1218 1250 1222
rect 1286 1218 1290 1222
rect 1238 1158 1242 1162
rect 1278 1158 1282 1162
rect 1302 1158 1306 1162
rect 1206 1148 1210 1152
rect 1294 1148 1298 1152
rect 1326 1148 1330 1152
rect 1238 1118 1242 1122
rect 1174 1088 1178 1092
rect 1070 1068 1074 1072
rect 1230 1068 1234 1072
rect 1102 1058 1106 1062
rect 990 1048 994 1052
rect 1006 1048 1010 1052
rect 1070 1048 1074 1052
rect 1166 1048 1170 1052
rect 1190 1048 1194 1052
rect 990 1038 994 1042
rect 910 1028 914 1032
rect 966 1028 970 1032
rect 974 1018 978 1022
rect 910 998 914 1002
rect 918 968 922 972
rect 902 958 906 962
rect 1086 1028 1090 1032
rect 1142 1008 1146 1012
rect 1094 988 1098 992
rect 1062 968 1066 972
rect 998 958 1002 962
rect 974 948 978 952
rect 910 928 914 932
rect 926 928 930 932
rect 1222 998 1226 1002
rect 1022 948 1026 952
rect 1206 947 1210 951
rect 1054 938 1058 942
rect 1094 938 1098 942
rect 1158 938 1162 942
rect 990 918 994 922
rect 942 888 946 892
rect 934 878 938 882
rect 822 868 826 872
rect 830 858 834 862
rect 814 848 818 852
rect 806 758 810 762
rect 790 748 794 752
rect 774 728 778 732
rect 798 728 802 732
rect 758 718 762 722
rect 734 708 738 712
rect 822 718 826 722
rect 958 858 962 862
rect 870 848 874 852
rect 926 848 930 852
rect 950 848 954 852
rect 974 848 978 852
rect 846 838 850 842
rect 862 828 866 832
rect 886 838 890 842
rect 950 838 954 842
rect 894 828 898 832
rect 926 828 930 832
rect 934 798 938 802
rect 838 778 842 782
rect 950 778 954 782
rect 934 768 938 772
rect 958 768 962 772
rect 990 878 994 882
rect 1046 928 1050 932
rect 998 868 1002 872
rect 1006 868 1010 872
rect 998 808 1002 812
rect 982 788 986 792
rect 998 788 1002 792
rect 974 768 978 772
rect 966 758 970 762
rect 1006 768 1010 772
rect 942 748 946 752
rect 958 748 962 752
rect 982 748 986 752
rect 838 738 842 742
rect 854 708 858 712
rect 718 678 722 682
rect 766 678 770 682
rect 774 678 778 682
rect 806 678 810 682
rect 710 668 714 672
rect 726 668 730 672
rect 470 658 474 662
rect 534 658 538 662
rect 582 658 586 662
rect 494 648 498 652
rect 502 648 506 652
rect 558 648 562 652
rect 406 638 410 642
rect 422 638 426 642
rect 462 638 466 642
rect 526 638 530 642
rect 550 638 554 642
rect 214 628 218 632
rect 310 628 314 632
rect 318 628 322 632
rect 334 628 338 632
rect 310 618 314 622
rect 238 608 242 612
rect 206 588 210 592
rect 230 588 234 592
rect 246 588 250 592
rect 278 588 282 592
rect 198 578 202 582
rect 182 558 186 562
rect 214 578 218 582
rect 270 568 274 572
rect 254 558 258 562
rect 294 558 298 562
rect 198 548 202 552
rect 230 548 234 552
rect 246 548 250 552
rect 278 548 282 552
rect 150 538 154 542
rect 174 538 178 542
rect 182 538 186 542
rect 262 538 266 542
rect 214 528 218 532
rect 134 518 138 522
rect 150 518 154 522
rect 102 478 106 482
rect 110 478 114 482
rect 102 458 106 462
rect 406 598 410 602
rect 574 638 578 642
rect 582 638 586 642
rect 702 638 706 642
rect 590 618 594 622
rect 602 603 606 607
rect 609 603 613 607
rect 590 598 594 602
rect 454 588 458 592
rect 462 588 466 592
rect 358 578 362 582
rect 350 568 354 572
rect 382 568 386 572
rect 414 568 418 572
rect 382 548 386 552
rect 414 548 418 552
rect 526 578 530 582
rect 390 538 394 542
rect 494 538 498 542
rect 326 528 330 532
rect 318 518 322 522
rect 358 528 362 532
rect 334 508 338 512
rect 158 488 162 492
rect 198 478 202 482
rect 286 478 290 482
rect 150 458 154 462
rect 190 458 194 462
rect 150 448 154 452
rect 158 448 162 452
rect 182 448 186 452
rect 118 438 122 442
rect 230 468 234 472
rect 270 468 274 472
rect 214 458 218 462
rect 222 458 226 462
rect 206 448 210 452
rect 182 428 186 432
rect 134 408 138 412
rect 70 388 74 392
rect 126 388 130 392
rect 22 368 26 372
rect 54 358 58 362
rect 6 338 10 342
rect 14 328 18 332
rect 6 298 10 302
rect 46 348 50 352
rect 70 348 74 352
rect 54 338 58 342
rect 30 328 34 332
rect 22 318 26 322
rect 46 318 50 322
rect 22 308 26 312
rect 110 348 114 352
rect 126 348 130 352
rect 70 288 74 292
rect 110 288 114 292
rect 38 278 42 282
rect 62 278 66 282
rect 14 188 18 192
rect 54 188 58 192
rect 22 178 26 182
rect 14 168 18 172
rect 30 168 34 172
rect 110 258 114 262
rect 118 258 122 262
rect 70 238 74 242
rect 78 238 82 242
rect 62 168 66 172
rect 22 158 26 162
rect 62 158 66 162
rect 54 148 58 152
rect 46 138 50 142
rect 102 248 106 252
rect 102 238 106 242
rect 94 228 98 232
rect 78 198 82 202
rect 150 398 154 402
rect 158 388 162 392
rect 174 378 178 382
rect 166 358 170 362
rect 182 358 186 362
rect 198 358 202 362
rect 182 348 186 352
rect 254 428 258 432
rect 246 418 250 422
rect 238 388 242 392
rect 230 378 234 382
rect 230 358 234 362
rect 214 348 218 352
rect 190 258 194 262
rect 134 248 138 252
rect 158 248 162 252
rect 134 238 138 242
rect 142 238 146 242
rect 86 168 90 172
rect 126 148 130 152
rect 198 238 202 242
rect 174 218 178 222
rect 182 208 186 212
rect 238 348 242 352
rect 254 338 258 342
rect 222 328 226 332
rect 246 328 250 332
rect 214 318 218 322
rect 286 458 290 462
rect 326 448 330 452
rect 318 438 322 442
rect 334 438 338 442
rect 350 438 354 442
rect 294 408 298 412
rect 302 408 306 412
rect 390 528 394 532
rect 414 528 418 532
rect 374 518 378 522
rect 438 528 442 532
rect 486 508 490 512
rect 430 498 434 502
rect 382 478 386 482
rect 414 478 418 482
rect 438 478 442 482
rect 470 478 474 482
rect 502 478 506 482
rect 382 468 386 472
rect 406 468 410 472
rect 454 468 458 472
rect 534 468 538 472
rect 438 458 442 462
rect 462 448 466 452
rect 470 448 474 452
rect 446 438 450 442
rect 518 438 522 442
rect 526 428 530 432
rect 430 418 434 422
rect 366 398 370 402
rect 278 388 282 392
rect 302 378 306 382
rect 398 378 402 382
rect 286 358 290 362
rect 318 358 322 362
rect 398 358 402 362
rect 422 358 426 362
rect 286 348 290 352
rect 390 338 394 342
rect 270 318 274 322
rect 366 328 370 332
rect 382 328 386 332
rect 334 318 338 322
rect 494 378 498 382
rect 510 378 514 382
rect 438 358 442 362
rect 462 338 466 342
rect 302 288 306 292
rect 342 288 346 292
rect 390 288 394 292
rect 406 288 410 292
rect 286 278 290 282
rect 326 278 330 282
rect 230 268 234 272
rect 278 268 282 272
rect 222 248 226 252
rect 278 258 282 262
rect 294 258 298 262
rect 262 248 266 252
rect 238 228 242 232
rect 238 208 242 212
rect 254 208 258 212
rect 142 178 146 182
rect 206 178 210 182
rect 214 178 218 182
rect 198 168 202 172
rect 110 138 114 142
rect 102 128 106 132
rect 118 98 122 102
rect 142 98 146 102
rect 126 88 130 92
rect 22 78 26 82
rect 46 78 50 82
rect 86 78 90 82
rect 14 68 18 72
rect 38 68 42 72
rect 86 68 90 72
rect 22 58 26 62
rect 38 48 42 52
rect 70 48 74 52
rect 46 8 50 12
rect 134 8 138 12
rect 222 168 226 172
rect 174 158 178 162
rect 206 158 210 162
rect 238 158 242 162
rect 190 148 194 152
rect 158 138 162 142
rect 230 138 234 142
rect 238 138 242 142
rect 246 138 250 142
rect 174 128 178 132
rect 166 88 170 92
rect 270 218 274 222
rect 286 168 290 172
rect 366 268 370 272
rect 398 268 402 272
rect 406 268 410 272
rect 350 258 354 262
rect 318 248 322 252
rect 342 248 346 252
rect 310 238 314 242
rect 302 168 306 172
rect 278 148 282 152
rect 270 138 274 142
rect 198 68 202 72
rect 206 68 210 72
rect 222 68 226 72
rect 254 68 258 72
rect 278 68 282 72
rect 342 228 346 232
rect 326 178 330 182
rect 334 148 338 152
rect 310 138 314 142
rect 350 158 354 162
rect 374 178 378 182
rect 454 328 458 332
rect 446 318 450 322
rect 478 348 482 352
rect 486 338 490 342
rect 502 318 506 322
rect 502 278 506 282
rect 502 258 506 262
rect 454 248 458 252
rect 494 218 498 222
rect 414 208 418 212
rect 414 188 418 192
rect 462 168 466 172
rect 382 158 386 162
rect 390 158 394 162
rect 446 148 450 152
rect 398 138 402 142
rect 414 138 418 142
rect 430 138 434 142
rect 366 128 370 132
rect 398 128 402 132
rect 414 128 418 132
rect 430 128 434 132
rect 454 128 458 132
rect 326 78 330 82
rect 318 68 322 72
rect 342 68 346 72
rect 358 68 362 72
rect 374 68 378 72
rect 158 58 162 62
rect 206 58 210 62
rect 294 58 298 62
rect 174 38 178 42
rect 278 18 282 22
rect 158 8 162 12
rect 422 68 426 72
rect 390 58 394 62
rect 350 48 354 52
rect 414 48 418 52
rect 422 48 426 52
rect 478 148 482 152
rect 558 438 562 442
rect 1038 878 1042 882
rect 990 738 994 742
rect 1022 738 1026 742
rect 974 708 978 712
rect 950 688 954 692
rect 894 678 898 682
rect 934 668 938 672
rect 734 628 738 632
rect 758 628 762 632
rect 734 618 738 622
rect 670 578 674 582
rect 710 568 714 572
rect 782 648 786 652
rect 814 638 818 642
rect 798 618 802 622
rect 862 598 866 602
rect 774 588 778 592
rect 926 658 930 662
rect 742 568 746 572
rect 862 568 866 572
rect 886 568 890 572
rect 734 558 738 562
rect 758 558 762 562
rect 574 548 578 552
rect 638 538 642 542
rect 702 538 706 542
rect 646 498 650 502
rect 638 478 642 482
rect 614 468 618 472
rect 582 448 586 452
rect 606 448 610 452
rect 590 438 594 442
rect 574 428 578 432
rect 602 403 606 407
rect 609 403 613 407
rect 758 538 762 542
rect 782 538 786 542
rect 726 528 730 532
rect 758 518 762 522
rect 726 478 730 482
rect 662 468 666 472
rect 718 468 722 472
rect 678 448 682 452
rect 718 448 722 452
rect 670 438 674 442
rect 654 428 658 432
rect 622 388 626 392
rect 590 378 594 382
rect 654 378 658 382
rect 542 368 546 372
rect 534 358 538 362
rect 558 358 562 362
rect 630 358 634 362
rect 566 348 570 352
rect 558 338 562 342
rect 550 328 554 332
rect 534 318 538 322
rect 614 348 618 352
rect 574 338 578 342
rect 582 328 586 332
rect 590 318 594 322
rect 550 268 554 272
rect 598 268 602 272
rect 526 258 530 262
rect 534 258 538 262
rect 678 428 682 432
rect 670 408 674 412
rect 830 558 834 562
rect 966 678 970 682
rect 982 678 986 682
rect 1030 728 1034 732
rect 1006 718 1010 722
rect 1014 688 1018 692
rect 958 668 962 672
rect 990 668 994 672
rect 958 658 962 662
rect 974 658 978 662
rect 998 658 1002 662
rect 998 638 1002 642
rect 1014 628 1018 632
rect 958 568 962 572
rect 950 528 954 532
rect 798 508 802 512
rect 790 498 794 502
rect 990 498 994 502
rect 1006 498 1010 502
rect 790 478 794 482
rect 942 478 946 482
rect 950 478 954 482
rect 750 468 754 472
rect 774 468 778 472
rect 822 468 826 472
rect 894 468 898 472
rect 918 468 922 472
rect 966 468 970 472
rect 702 438 706 442
rect 742 428 746 432
rect 686 378 690 382
rect 646 358 650 362
rect 662 358 666 362
rect 726 378 730 382
rect 702 358 706 362
rect 694 348 698 352
rect 646 338 650 342
rect 766 358 770 362
rect 814 458 818 462
rect 886 458 890 462
rect 830 448 834 452
rect 926 448 930 452
rect 934 448 938 452
rect 798 418 802 422
rect 750 348 754 352
rect 766 348 770 352
rect 734 338 738 342
rect 678 328 682 332
rect 766 338 770 342
rect 782 338 786 342
rect 750 328 754 332
rect 742 318 746 322
rect 678 288 682 292
rect 758 288 762 292
rect 638 278 642 282
rect 694 278 698 282
rect 734 278 738 282
rect 566 258 570 262
rect 582 258 586 262
rect 614 258 618 262
rect 630 258 634 262
rect 534 248 538 252
rect 574 248 578 252
rect 606 248 610 252
rect 542 228 546 232
rect 566 228 570 232
rect 590 218 594 222
rect 622 218 626 222
rect 582 168 586 172
rect 542 158 546 162
rect 518 148 522 152
rect 502 138 506 142
rect 518 138 522 142
rect 526 138 530 142
rect 486 128 490 132
rect 494 118 498 122
rect 574 148 578 152
rect 542 78 546 82
rect 550 78 554 82
rect 582 78 586 82
rect 478 68 482 72
rect 454 48 458 52
rect 478 38 482 42
rect 602 203 606 207
rect 609 203 613 207
rect 654 268 658 272
rect 678 268 682 272
rect 686 258 690 262
rect 670 248 674 252
rect 638 168 642 172
rect 646 168 650 172
rect 622 138 626 142
rect 614 128 618 132
rect 598 118 602 122
rect 694 208 698 212
rect 670 168 674 172
rect 686 168 690 172
rect 734 208 738 212
rect 710 178 714 182
rect 734 168 738 172
rect 710 158 714 162
rect 726 158 730 162
rect 662 148 666 152
rect 694 148 698 152
rect 670 108 674 112
rect 734 148 738 152
rect 750 218 754 222
rect 814 408 818 412
rect 822 358 826 362
rect 822 348 826 352
rect 1046 659 1050 663
rect 1022 568 1026 572
rect 1022 468 1026 472
rect 1030 468 1034 472
rect 1006 458 1010 462
rect 1014 458 1018 462
rect 1046 458 1050 462
rect 846 438 850 442
rect 862 438 866 442
rect 902 438 906 442
rect 958 438 962 442
rect 974 438 978 442
rect 894 408 898 412
rect 950 408 954 412
rect 910 398 914 402
rect 862 378 866 382
rect 886 358 890 362
rect 894 358 898 362
rect 974 378 978 382
rect 982 378 986 382
rect 934 358 938 362
rect 974 358 978 362
rect 998 358 1002 362
rect 1006 358 1010 362
rect 950 348 954 352
rect 830 338 834 342
rect 870 338 874 342
rect 894 338 898 342
rect 910 338 914 342
rect 974 338 978 342
rect 990 338 994 342
rect 838 328 842 332
rect 862 328 866 332
rect 910 318 914 322
rect 918 318 922 322
rect 918 308 922 312
rect 982 308 986 312
rect 814 278 818 282
rect 854 278 858 282
rect 894 278 898 282
rect 782 268 786 272
rect 846 268 850 272
rect 854 268 858 272
rect 798 258 802 262
rect 766 218 770 222
rect 758 148 762 152
rect 782 148 786 152
rect 742 128 746 132
rect 758 128 762 132
rect 790 128 794 132
rect 654 88 658 92
rect 726 118 730 122
rect 774 98 778 102
rect 606 78 610 82
rect 702 78 706 82
rect 710 78 714 82
rect 750 78 754 82
rect 742 68 746 72
rect 558 58 562 62
rect 678 58 682 62
rect 782 58 786 62
rect 806 248 810 252
rect 830 218 834 222
rect 814 168 818 172
rect 838 168 842 172
rect 822 158 826 162
rect 806 148 810 152
rect 814 148 818 152
rect 830 118 834 122
rect 854 218 858 222
rect 870 258 874 262
rect 862 198 866 202
rect 886 268 890 272
rect 878 188 882 192
rect 854 168 858 172
rect 878 168 882 172
rect 854 158 858 162
rect 910 218 914 222
rect 926 298 930 302
rect 1022 438 1026 442
rect 1054 448 1058 452
rect 1062 408 1066 412
rect 1046 398 1050 402
rect 1030 368 1034 372
rect 1022 358 1026 362
rect 1094 928 1098 932
rect 1134 928 1138 932
rect 1118 918 1122 922
rect 1114 903 1118 907
rect 1121 903 1125 907
rect 1134 868 1138 872
rect 1118 858 1122 862
rect 1118 848 1122 852
rect 1094 838 1098 842
rect 1118 768 1122 772
rect 1110 728 1114 732
rect 1114 703 1118 707
rect 1121 703 1125 707
rect 1118 688 1122 692
rect 1102 678 1106 682
rect 1158 928 1162 932
rect 1166 908 1170 912
rect 1182 888 1186 892
rect 1190 888 1194 892
rect 1174 878 1178 882
rect 1254 1058 1258 1062
rect 1238 1018 1242 1022
rect 1270 1118 1274 1122
rect 1318 1118 1322 1122
rect 1278 1078 1282 1082
rect 1302 1078 1306 1082
rect 1646 1538 1650 1542
rect 1614 1528 1618 1532
rect 1606 1518 1610 1522
rect 1598 1508 1602 1512
rect 1574 1488 1578 1492
rect 1614 1478 1618 1482
rect 1550 1468 1554 1472
rect 1526 1458 1530 1462
rect 1510 1438 1514 1442
rect 1558 1438 1562 1442
rect 1582 1448 1586 1452
rect 1574 1428 1578 1432
rect 1526 1398 1530 1402
rect 1550 1398 1554 1402
rect 1510 1388 1514 1392
rect 1590 1408 1594 1412
rect 1534 1378 1538 1382
rect 1574 1378 1578 1382
rect 1662 1468 1666 1472
rect 1662 1458 1666 1462
rect 1614 1438 1618 1442
rect 1670 1438 1674 1442
rect 1614 1418 1618 1422
rect 1694 1478 1698 1482
rect 1678 1428 1682 1432
rect 1502 1368 1506 1372
rect 1574 1368 1578 1372
rect 1630 1368 1634 1372
rect 1510 1358 1514 1362
rect 1590 1358 1594 1362
rect 1678 1358 1682 1362
rect 1462 1328 1466 1332
rect 1470 1308 1474 1312
rect 1454 1298 1458 1302
rect 1422 1278 1426 1282
rect 1446 1278 1450 1282
rect 1398 1228 1402 1232
rect 1374 1218 1378 1222
rect 1446 1228 1450 1232
rect 1510 1338 1514 1342
rect 1494 1298 1498 1302
rect 1486 1278 1490 1282
rect 1558 1340 1562 1344
rect 1646 1348 1650 1352
rect 1662 1348 1666 1352
rect 1582 1338 1586 1342
rect 1598 1338 1602 1342
rect 1622 1338 1626 1342
rect 1654 1338 1658 1342
rect 1670 1338 1674 1342
rect 1566 1318 1570 1322
rect 1542 1298 1546 1302
rect 1550 1288 1554 1292
rect 1358 1158 1362 1162
rect 1390 1158 1394 1162
rect 1358 1148 1362 1152
rect 1406 1148 1410 1152
rect 1366 1068 1370 1072
rect 1270 1058 1274 1062
rect 1302 1058 1306 1062
rect 1326 1058 1330 1062
rect 1302 1048 1306 1052
rect 1262 1018 1266 1022
rect 1246 1008 1250 1012
rect 1262 998 1266 1002
rect 1270 998 1274 1002
rect 1318 1038 1322 1042
rect 1254 898 1258 902
rect 1286 898 1290 902
rect 1198 868 1202 872
rect 1230 868 1234 872
rect 1158 848 1162 852
rect 1166 738 1170 742
rect 1470 1168 1474 1172
rect 1494 1168 1498 1172
rect 1534 1258 1538 1262
rect 1518 1168 1522 1172
rect 1526 1168 1530 1172
rect 1518 1158 1522 1162
rect 1550 1278 1554 1282
rect 1558 1258 1562 1262
rect 1574 1298 1578 1302
rect 1590 1298 1594 1302
rect 1582 1288 1586 1292
rect 1614 1318 1618 1322
rect 1662 1318 1666 1322
rect 1630 1308 1634 1312
rect 1614 1278 1618 1282
rect 1662 1268 1666 1272
rect 1670 1268 1674 1272
rect 1606 1258 1610 1262
rect 1622 1258 1626 1262
rect 1606 1248 1610 1252
rect 1566 1238 1570 1242
rect 1614 1238 1618 1242
rect 1582 1168 1586 1172
rect 1606 1158 1610 1162
rect 1478 1148 1482 1152
rect 1398 1138 1402 1142
rect 1406 1128 1410 1132
rect 1422 1128 1426 1132
rect 1382 1118 1386 1122
rect 1422 1118 1426 1122
rect 1414 1088 1418 1092
rect 1382 1078 1386 1082
rect 1398 1068 1402 1072
rect 1374 1048 1378 1052
rect 1390 1048 1394 1052
rect 1334 1028 1338 1032
rect 1374 1028 1378 1032
rect 1366 1008 1370 1012
rect 1382 1018 1386 1022
rect 1382 988 1386 992
rect 1422 988 1426 992
rect 1350 948 1354 952
rect 1326 938 1330 942
rect 1446 1128 1450 1132
rect 1454 1038 1458 1042
rect 1398 948 1402 952
rect 1398 928 1402 932
rect 1366 888 1370 892
rect 1294 878 1298 882
rect 1262 848 1266 852
rect 1294 858 1298 862
rect 1350 848 1354 852
rect 1278 828 1282 832
rect 1334 828 1338 832
rect 1422 918 1426 922
rect 1422 898 1426 902
rect 1406 888 1410 892
rect 1446 958 1450 962
rect 1438 878 1442 882
rect 1454 908 1458 912
rect 1678 1148 1682 1152
rect 1518 1138 1522 1142
rect 1542 1138 1546 1142
rect 1566 1138 1570 1142
rect 1598 1138 1602 1142
rect 1614 1138 1618 1142
rect 1502 1128 1506 1132
rect 1526 1128 1530 1132
rect 1550 1128 1554 1132
rect 1574 1128 1578 1132
rect 1718 1348 1722 1352
rect 1718 1148 1722 1152
rect 1694 1108 1698 1112
rect 1710 1108 1714 1112
rect 1510 958 1514 962
rect 1590 1038 1594 1042
rect 1510 948 1514 952
rect 1526 948 1530 952
rect 1558 948 1562 952
rect 1478 868 1482 872
rect 1446 848 1450 852
rect 1438 798 1442 802
rect 1366 788 1370 792
rect 1398 788 1402 792
rect 1398 768 1402 772
rect 1366 758 1370 762
rect 1166 718 1170 722
rect 1102 668 1106 672
rect 1150 668 1154 672
rect 1094 638 1098 642
rect 1110 638 1114 642
rect 1430 738 1434 742
rect 1206 678 1210 682
rect 1278 678 1282 682
rect 1334 678 1338 682
rect 1182 668 1186 672
rect 1286 668 1290 672
rect 1302 658 1306 662
rect 1318 658 1322 662
rect 1366 658 1370 662
rect 1222 648 1226 652
rect 1398 728 1402 732
rect 1422 688 1426 692
rect 1422 668 1426 672
rect 1382 658 1386 662
rect 1342 588 1346 592
rect 1078 578 1082 582
rect 1094 578 1098 582
rect 1358 578 1362 582
rect 1422 578 1426 582
rect 1430 578 1434 582
rect 1086 568 1090 572
rect 1182 568 1186 572
rect 1190 568 1194 572
rect 1102 558 1106 562
rect 1150 558 1154 562
rect 1086 538 1090 542
rect 1078 498 1082 502
rect 1086 458 1090 462
rect 1086 448 1090 452
rect 1158 548 1162 552
rect 1118 538 1122 542
rect 1222 548 1226 552
rect 1366 558 1370 562
rect 1406 558 1410 562
rect 1430 558 1434 562
rect 1214 538 1218 542
rect 1230 538 1234 542
rect 1254 538 1258 542
rect 1286 538 1290 542
rect 1350 538 1354 542
rect 1190 528 1194 532
rect 1166 508 1170 512
rect 1114 503 1118 507
rect 1121 503 1125 507
rect 1102 498 1106 502
rect 1182 498 1186 502
rect 1206 498 1210 502
rect 1134 468 1138 472
rect 1126 458 1130 462
rect 1110 428 1114 432
rect 1110 418 1114 422
rect 1102 398 1106 402
rect 1094 378 1098 382
rect 1046 358 1050 362
rect 1086 358 1090 362
rect 1046 348 1050 352
rect 1038 298 1042 302
rect 1054 298 1058 302
rect 958 288 962 292
rect 998 288 1002 292
rect 950 268 954 272
rect 982 268 986 272
rect 1006 268 1010 272
rect 950 248 954 252
rect 1006 248 1010 252
rect 942 218 946 222
rect 958 198 962 202
rect 934 168 938 172
rect 942 158 946 162
rect 910 148 914 152
rect 926 148 930 152
rect 854 118 858 122
rect 878 118 882 122
rect 846 108 850 112
rect 806 88 810 92
rect 854 88 858 92
rect 846 78 850 82
rect 814 68 818 72
rect 838 68 842 72
rect 566 38 570 42
rect 438 28 442 32
rect 510 28 514 32
rect 454 18 458 22
rect 686 18 690 22
rect 790 8 794 12
rect 798 8 802 12
rect 814 8 818 12
rect 602 3 606 7
rect 609 3 613 7
rect 974 168 978 172
rect 894 128 898 132
rect 910 128 914 132
rect 902 108 906 112
rect 1030 208 1034 212
rect 1094 338 1098 342
rect 1174 458 1178 462
rect 1134 448 1138 452
rect 1150 448 1154 452
rect 1142 358 1146 362
rect 1086 328 1090 332
rect 1070 268 1074 272
rect 1114 303 1118 307
rect 1121 303 1125 307
rect 1110 288 1114 292
rect 1102 278 1106 282
rect 1078 248 1082 252
rect 1054 238 1058 242
rect 1006 178 1010 182
rect 1038 178 1042 182
rect 1014 168 1018 172
rect 1022 158 1026 162
rect 1046 158 1050 162
rect 966 108 970 112
rect 990 88 994 92
rect 966 78 970 82
rect 886 68 890 72
rect 926 68 930 72
rect 966 68 970 72
rect 998 78 1002 82
rect 982 58 986 62
rect 1006 58 1010 62
rect 918 28 922 32
rect 950 18 954 22
rect 918 8 922 12
rect 982 8 986 12
rect 1038 148 1042 152
rect 1078 218 1082 222
rect 1086 218 1090 222
rect 1126 268 1130 272
rect 1142 288 1146 292
rect 1278 528 1282 532
rect 1230 508 1234 512
rect 1262 508 1266 512
rect 1286 498 1290 502
rect 1206 478 1210 482
rect 1190 468 1194 472
rect 1214 468 1218 472
rect 1238 458 1242 462
rect 1270 458 1274 462
rect 1302 458 1306 462
rect 1246 448 1250 452
rect 1270 448 1274 452
rect 1206 408 1210 412
rect 1166 398 1170 402
rect 1198 378 1202 382
rect 1166 338 1170 342
rect 1182 358 1186 362
rect 1182 338 1186 342
rect 1190 338 1194 342
rect 1206 338 1210 342
rect 1174 308 1178 312
rect 1246 438 1250 442
rect 1262 438 1266 442
rect 1254 418 1258 422
rect 1246 378 1250 382
rect 1254 338 1258 342
rect 1230 328 1234 332
rect 1174 298 1178 302
rect 1214 298 1218 302
rect 1334 518 1338 522
rect 1326 488 1330 492
rect 1510 918 1514 922
rect 1590 908 1594 912
rect 1526 898 1530 902
rect 1646 1048 1650 1052
rect 1654 1038 1658 1042
rect 1630 918 1634 922
rect 1678 978 1682 982
rect 1630 868 1634 872
rect 1670 868 1674 872
rect 1486 848 1490 852
rect 1454 838 1458 842
rect 1470 808 1474 812
rect 1462 768 1466 772
rect 1558 758 1562 762
rect 1518 748 1522 752
rect 1494 738 1498 742
rect 1526 738 1530 742
rect 1454 728 1458 732
rect 1478 728 1482 732
rect 1470 658 1474 662
rect 1678 858 1682 862
rect 1654 848 1658 852
rect 1550 688 1554 692
rect 1534 678 1538 682
rect 1550 658 1554 662
rect 1590 658 1594 662
rect 1486 648 1490 652
rect 1606 648 1610 652
rect 1662 788 1666 792
rect 1710 938 1714 942
rect 1718 918 1722 922
rect 1710 898 1714 902
rect 1702 858 1706 862
rect 1726 888 1730 892
rect 1726 878 1730 882
rect 1702 848 1706 852
rect 1694 788 1698 792
rect 1702 718 1706 722
rect 1710 718 1714 722
rect 1694 698 1698 702
rect 1734 678 1738 682
rect 1734 628 1738 632
rect 1662 608 1666 612
rect 1486 588 1490 592
rect 1566 588 1570 592
rect 1454 578 1458 582
rect 1462 578 1466 582
rect 1510 578 1514 582
rect 1510 568 1514 572
rect 1494 558 1498 562
rect 1462 548 1466 552
rect 1446 538 1450 542
rect 1438 528 1442 532
rect 1390 478 1394 482
rect 1462 478 1466 482
rect 1374 468 1378 472
rect 1318 438 1322 442
rect 1342 438 1346 442
rect 1302 418 1306 422
rect 1286 408 1290 412
rect 1366 458 1370 462
rect 1374 448 1378 452
rect 1358 388 1362 392
rect 1486 528 1490 532
rect 1422 468 1426 472
rect 1470 468 1474 472
rect 1478 468 1482 472
rect 1382 378 1386 382
rect 1334 368 1338 372
rect 1278 358 1282 362
rect 1374 358 1378 362
rect 1342 348 1346 352
rect 1326 338 1330 342
rect 1278 328 1282 332
rect 1278 298 1282 302
rect 1294 298 1298 302
rect 1246 288 1250 292
rect 1158 278 1162 282
rect 1198 278 1202 282
rect 1150 268 1154 272
rect 1174 268 1178 272
rect 1150 248 1154 252
rect 1158 248 1162 252
rect 1134 228 1138 232
rect 1118 218 1122 222
rect 1166 218 1170 222
rect 1110 208 1114 212
rect 1094 188 1098 192
rect 1062 178 1066 182
rect 1038 118 1042 122
rect 1078 148 1082 152
rect 1222 258 1226 262
rect 1230 258 1234 262
rect 1318 328 1322 332
rect 1342 328 1346 332
rect 1278 278 1282 282
rect 1262 268 1266 272
rect 1230 248 1234 252
rect 1254 248 1258 252
rect 1198 238 1202 242
rect 1238 238 1242 242
rect 1246 208 1250 212
rect 1230 188 1234 192
rect 1134 178 1138 182
rect 1150 178 1154 182
rect 1174 178 1178 182
rect 1238 178 1242 182
rect 1126 168 1130 172
rect 1102 148 1106 152
rect 1222 168 1226 172
rect 1150 158 1154 162
rect 1158 158 1162 162
rect 1166 158 1170 162
rect 1302 268 1306 272
rect 1318 258 1322 262
rect 1366 328 1370 332
rect 1374 328 1378 332
rect 1366 318 1370 322
rect 1358 298 1362 302
rect 1406 458 1410 462
rect 1438 448 1442 452
rect 1470 438 1474 442
rect 1414 418 1418 422
rect 1446 418 1450 422
rect 1398 368 1402 372
rect 1414 368 1418 372
rect 1422 368 1426 372
rect 1550 558 1554 562
rect 1518 528 1522 532
rect 1494 448 1498 452
rect 1510 448 1514 452
rect 1510 438 1514 442
rect 1598 558 1602 562
rect 1574 528 1578 532
rect 1598 528 1602 532
rect 1566 488 1570 492
rect 1542 468 1546 472
rect 1558 468 1562 472
rect 1534 458 1538 462
rect 1486 418 1490 422
rect 1502 418 1506 422
rect 1486 408 1490 412
rect 1478 398 1482 402
rect 1510 398 1514 402
rect 1486 368 1490 372
rect 1390 348 1394 352
rect 1414 348 1418 352
rect 1430 338 1434 342
rect 1438 338 1442 342
rect 1398 298 1402 302
rect 1630 548 1634 552
rect 1646 548 1650 552
rect 1702 538 1706 542
rect 1694 528 1698 532
rect 1662 498 1666 502
rect 1582 468 1586 472
rect 1630 468 1634 472
rect 1574 458 1578 462
rect 1590 428 1594 432
rect 1542 418 1546 422
rect 1566 418 1570 422
rect 1534 388 1538 392
rect 1566 368 1570 372
rect 1526 358 1530 362
rect 1454 348 1458 352
rect 1462 328 1466 332
rect 1446 318 1450 322
rect 1374 278 1378 282
rect 1398 268 1402 272
rect 1422 268 1426 272
rect 1438 258 1442 262
rect 1326 248 1330 252
rect 1350 248 1354 252
rect 1358 248 1362 252
rect 1294 228 1298 232
rect 1286 218 1290 222
rect 1310 188 1314 192
rect 1270 168 1274 172
rect 1246 158 1250 162
rect 1174 148 1178 152
rect 1190 148 1194 152
rect 1086 128 1090 132
rect 1094 128 1098 132
rect 1126 128 1130 132
rect 1150 128 1154 132
rect 1062 118 1066 122
rect 1114 103 1118 107
rect 1121 103 1125 107
rect 1030 88 1034 92
rect 1046 88 1050 92
rect 1102 88 1106 92
rect 1054 78 1058 82
rect 1078 78 1082 82
rect 1134 78 1138 82
rect 1118 68 1122 72
rect 1022 18 1026 22
rect 1038 18 1042 22
rect 1078 18 1082 22
rect 1102 18 1106 22
rect 1062 8 1066 12
rect 1166 68 1170 72
rect 1142 58 1146 62
rect 1206 128 1210 132
rect 1190 118 1194 122
rect 1182 108 1186 112
rect 1246 118 1250 122
rect 1198 108 1202 112
rect 1214 108 1218 112
rect 1238 108 1242 112
rect 1198 88 1202 92
rect 1166 8 1170 12
rect 1174 8 1178 12
rect 1270 158 1274 162
rect 1278 148 1282 152
rect 1294 148 1298 152
rect 1302 128 1306 132
rect 1350 238 1354 242
rect 1390 238 1394 242
rect 1406 238 1410 242
rect 1334 208 1338 212
rect 1438 178 1442 182
rect 1342 158 1346 162
rect 1414 158 1418 162
rect 1350 138 1354 142
rect 1382 138 1386 142
rect 1326 128 1330 132
rect 1286 88 1290 92
rect 1334 118 1338 122
rect 1366 118 1370 122
rect 1366 108 1370 112
rect 1374 98 1378 102
rect 1382 98 1386 102
rect 1406 138 1410 142
rect 1414 108 1418 112
rect 1398 98 1402 102
rect 1334 88 1338 92
rect 1382 88 1386 92
rect 1326 78 1330 82
rect 1230 68 1234 72
rect 1246 68 1250 72
rect 1294 58 1298 62
rect 1278 48 1282 52
rect 1238 38 1242 42
rect 1262 38 1266 42
rect 1214 8 1218 12
rect 1222 8 1226 12
rect 1238 8 1242 12
rect 1438 118 1442 122
rect 1422 98 1426 102
rect 1510 348 1514 352
rect 1542 338 1546 342
rect 1470 318 1474 322
rect 1478 318 1482 322
rect 1494 318 1498 322
rect 1502 318 1506 322
rect 1518 318 1522 322
rect 1486 268 1490 272
rect 1590 348 1594 352
rect 1566 288 1570 292
rect 1534 268 1538 272
rect 1510 258 1514 262
rect 1526 258 1530 262
rect 1478 248 1482 252
rect 1518 248 1522 252
rect 1470 208 1474 212
rect 1502 238 1506 242
rect 1534 238 1538 242
rect 1494 208 1498 212
rect 1518 188 1522 192
rect 1510 168 1514 172
rect 1502 158 1506 162
rect 1494 148 1498 152
rect 1478 138 1482 142
rect 1590 298 1594 302
rect 1702 518 1706 522
rect 1694 478 1698 482
rect 1710 488 1714 492
rect 1662 458 1666 462
rect 1678 458 1682 462
rect 1686 458 1690 462
rect 1606 448 1610 452
rect 1638 448 1642 452
rect 1614 418 1618 422
rect 1614 398 1618 402
rect 1670 448 1674 452
rect 1702 448 1706 452
rect 1654 438 1658 442
rect 1678 438 1682 442
rect 1646 428 1650 432
rect 1638 408 1642 412
rect 1630 388 1634 392
rect 1622 368 1626 372
rect 1654 398 1658 402
rect 1678 378 1682 382
rect 1702 368 1706 372
rect 1622 358 1626 362
rect 1630 358 1634 362
rect 1662 358 1666 362
rect 1702 358 1706 362
rect 1614 348 1618 352
rect 1630 348 1634 352
rect 1614 338 1618 342
rect 1598 278 1602 282
rect 1558 198 1562 202
rect 1590 238 1594 242
rect 1630 258 1634 262
rect 1622 248 1626 252
rect 1582 188 1586 192
rect 1590 168 1594 172
rect 1526 158 1530 162
rect 1542 158 1546 162
rect 1574 158 1578 162
rect 1598 158 1602 162
rect 1542 148 1546 152
rect 1574 148 1578 152
rect 1582 148 1586 152
rect 1454 128 1458 132
rect 1542 108 1546 112
rect 1526 98 1530 102
rect 1566 118 1570 122
rect 1550 98 1554 102
rect 1598 138 1602 142
rect 1590 118 1594 122
rect 1462 88 1466 92
rect 1486 88 1490 92
rect 1518 88 1522 92
rect 1550 88 1554 92
rect 1342 68 1346 72
rect 1350 68 1354 72
rect 1358 58 1362 62
rect 1406 58 1410 62
rect 1526 78 1530 82
rect 1574 78 1578 82
rect 1614 208 1618 212
rect 1662 348 1666 352
rect 1718 348 1722 352
rect 1678 338 1682 342
rect 1694 308 1698 312
rect 1686 288 1690 292
rect 1678 278 1682 282
rect 1710 278 1714 282
rect 1694 268 1698 272
rect 1718 258 1722 262
rect 1646 208 1650 212
rect 1654 198 1658 202
rect 1638 158 1642 162
rect 1710 188 1714 192
rect 1630 148 1634 152
rect 1686 148 1690 152
rect 1662 138 1666 142
rect 1622 108 1626 112
rect 1678 128 1682 132
rect 1694 128 1698 132
rect 1670 98 1674 102
rect 1662 88 1666 92
rect 1662 78 1666 82
rect 1494 68 1498 72
rect 1686 68 1690 72
rect 1430 48 1434 52
rect 1470 38 1474 42
rect 1302 28 1306 32
rect 1374 28 1378 32
rect 1326 8 1330 12
rect 1710 66 1714 70
rect 1694 58 1698 62
rect 1734 58 1738 62
rect 1558 18 1562 22
<< metal3 >>
rect 282 1608 446 1611
rect 626 1608 630 1611
rect 1234 1608 1238 1611
rect 600 1603 602 1607
rect 606 1603 609 1607
rect 614 1603 616 1607
rect 694 1602 697 1608
rect 66 1588 118 1591
rect 122 1588 358 1591
rect 682 1588 710 1591
rect 206 1578 534 1581
rect 538 1578 630 1581
rect 634 1578 646 1581
rect 674 1578 678 1581
rect 206 1572 209 1578
rect 250 1568 686 1571
rect 690 1568 726 1571
rect 1402 1568 1478 1571
rect 1502 1568 1510 1571
rect 1514 1568 1590 1571
rect 206 1561 209 1568
rect 162 1558 209 1561
rect 370 1558 374 1561
rect 426 1558 542 1561
rect 626 1558 702 1561
rect 762 1558 790 1561
rect 902 1561 905 1568
rect 794 1558 905 1561
rect 978 1558 998 1561
rect 1010 1558 1070 1561
rect 1162 1558 1166 1561
rect 1222 1558 1294 1561
rect 1434 1558 1550 1561
rect 402 1548 518 1551
rect 562 1548 582 1551
rect 586 1548 606 1551
rect 610 1548 646 1551
rect 650 1548 718 1551
rect 778 1548 806 1551
rect 810 1548 934 1551
rect 938 1548 1094 1551
rect 1222 1551 1225 1558
rect 1170 1548 1225 1551
rect 1234 1548 1238 1551
rect 1298 1548 1310 1551
rect 1322 1548 1326 1551
rect 1386 1548 1414 1551
rect 1474 1548 1478 1551
rect 1498 1548 1518 1551
rect 1602 1548 1649 1551
rect 190 1542 193 1548
rect 1646 1542 1649 1548
rect 98 1538 126 1541
rect 130 1538 166 1541
rect 170 1538 182 1541
rect 226 1538 254 1541
rect 290 1538 318 1541
rect 354 1538 366 1541
rect 386 1538 422 1541
rect 426 1538 446 1541
rect 482 1538 494 1541
rect 510 1538 702 1541
rect 706 1538 750 1541
rect 754 1538 806 1541
rect 858 1538 942 1541
rect 970 1538 1094 1541
rect 1098 1538 1118 1541
rect 1146 1538 1150 1541
rect 1154 1538 1182 1541
rect 1234 1538 1390 1541
rect 1418 1538 1422 1541
rect 1514 1538 1550 1541
rect 406 1532 409 1538
rect 510 1532 513 1538
rect -26 1531 -22 1532
rect -26 1528 86 1531
rect 90 1528 110 1531
rect 114 1528 286 1531
rect 290 1528 310 1531
rect 338 1528 406 1531
rect 746 1528 766 1531
rect 966 1531 969 1538
rect 914 1528 969 1531
rect 986 1528 998 1531
rect 1002 1528 1094 1531
rect 1226 1528 1254 1531
rect 1306 1528 1310 1531
rect 1322 1528 1326 1531
rect 1342 1528 1438 1531
rect 1442 1528 1470 1531
rect 1474 1528 1526 1531
rect 1554 1528 1614 1531
rect 742 1522 745 1528
rect 870 1522 873 1528
rect 1342 1522 1345 1528
rect 10 1518 182 1521
rect 186 1518 366 1521
rect 466 1518 518 1521
rect 530 1518 550 1521
rect 938 1518 966 1521
rect 986 1518 1006 1521
rect 1042 1518 1046 1521
rect 1226 1518 1238 1521
rect 1378 1518 1446 1521
rect 1538 1518 1606 1521
rect 1062 1512 1065 1518
rect 306 1508 422 1511
rect 426 1508 454 1511
rect 506 1508 574 1511
rect 874 1508 958 1511
rect 994 1508 1014 1511
rect 1274 1508 1374 1511
rect 1490 1508 1542 1511
rect 1546 1508 1598 1511
rect 1112 1503 1114 1507
rect 1118 1503 1121 1507
rect 1126 1503 1128 1507
rect 358 1498 550 1501
rect 554 1498 566 1501
rect 882 1498 910 1501
rect 1178 1498 1190 1501
rect 1202 1498 1462 1501
rect 358 1492 361 1498
rect 66 1488 70 1491
rect 202 1488 358 1491
rect 370 1488 486 1491
rect 490 1488 502 1491
rect 738 1488 766 1491
rect 778 1488 798 1491
rect 802 1488 910 1491
rect 1026 1488 1238 1491
rect 1242 1488 1366 1491
rect 1370 1488 1574 1491
rect -26 1481 -22 1482
rect -26 1478 54 1481
rect 122 1478 190 1481
rect 250 1478 302 1481
rect 450 1478 462 1481
rect 690 1478 702 1481
rect 730 1478 790 1481
rect 794 1478 822 1481
rect 910 1481 913 1488
rect 910 1478 950 1481
rect 954 1478 958 1481
rect 970 1478 1030 1481
rect 1106 1478 1166 1481
rect 1170 1478 1214 1481
rect 1218 1478 1286 1481
rect 1618 1478 1694 1481
rect 58 1468 70 1471
rect 178 1468 182 1471
rect 218 1468 246 1471
rect 322 1468 350 1471
rect 538 1468 582 1471
rect 638 1468 646 1471
rect 650 1468 654 1471
rect 670 1471 673 1478
rect 670 1468 686 1471
rect 746 1468 753 1471
rect 762 1468 790 1471
rect 794 1468 854 1471
rect 862 1471 865 1478
rect 894 1471 897 1478
rect 862 1468 897 1471
rect 906 1468 926 1471
rect 930 1468 998 1471
rect 1098 1468 1126 1471
rect 1130 1468 1142 1471
rect 1162 1468 1206 1471
rect 1258 1468 1318 1471
rect 1426 1468 1446 1471
rect 1466 1468 1550 1471
rect 1658 1468 1662 1471
rect -26 1461 -22 1462
rect -26 1458 6 1461
rect 38 1461 41 1468
rect 34 1458 41 1461
rect 50 1458 62 1461
rect 66 1458 78 1461
rect 138 1458 142 1461
rect 158 1461 161 1468
rect 750 1462 753 1468
rect 146 1458 262 1461
rect 266 1458 278 1461
rect 386 1458 398 1461
rect 506 1458 526 1461
rect 594 1458 678 1461
rect 850 1458 862 1461
rect 930 1458 934 1461
rect 954 1458 974 1461
rect 994 1458 1014 1461
rect 1066 1458 1070 1461
rect 1074 1458 1110 1461
rect 1154 1458 1254 1461
rect 1330 1458 1398 1461
rect 1402 1458 1526 1461
rect 10 1448 118 1451
rect 210 1448 310 1451
rect 462 1451 465 1458
rect 442 1448 465 1451
rect 482 1448 558 1451
rect 562 1448 646 1451
rect 690 1448 758 1451
rect 898 1448 942 1451
rect 1074 1448 1134 1451
rect 1162 1448 1182 1451
rect 1270 1451 1273 1458
rect 1662 1452 1665 1458
rect 1194 1448 1273 1451
rect 1362 1448 1430 1451
rect 1558 1448 1582 1451
rect 1558 1442 1561 1448
rect 66 1438 70 1441
rect 258 1438 622 1441
rect 626 1438 630 1441
rect 650 1438 782 1441
rect 946 1438 1017 1441
rect 1014 1432 1017 1438
rect 1078 1438 1094 1441
rect 1130 1438 1206 1441
rect 1210 1438 1230 1441
rect 1322 1438 1406 1441
rect 1410 1438 1510 1441
rect 1618 1438 1670 1441
rect 1062 1432 1065 1438
rect 1078 1432 1081 1438
rect 58 1428 62 1431
rect 298 1428 334 1431
rect 1214 1428 1422 1431
rect 1426 1428 1574 1431
rect 1650 1428 1678 1431
rect 446 1421 449 1428
rect 446 1418 790 1421
rect 914 1418 1006 1421
rect 1214 1421 1217 1428
rect 1034 1418 1217 1421
rect 1226 1418 1286 1421
rect 1330 1418 1390 1421
rect 1498 1418 1614 1421
rect 34 1408 86 1411
rect 90 1408 198 1411
rect 890 1408 1054 1411
rect 1290 1408 1382 1411
rect 1442 1408 1590 1411
rect 600 1403 602 1407
rect 606 1403 609 1407
rect 614 1403 616 1407
rect 26 1398 38 1401
rect 378 1398 574 1401
rect 1002 1398 1014 1401
rect 1138 1398 1302 1401
rect 1306 1398 1366 1401
rect 1370 1398 1478 1401
rect 1530 1398 1550 1401
rect 234 1388 286 1391
rect 482 1388 510 1391
rect 994 1388 1022 1391
rect 1270 1388 1278 1391
rect 1282 1388 1350 1391
rect 1514 1388 1537 1391
rect 22 1381 25 1388
rect 22 1378 54 1381
rect 138 1378 265 1381
rect 262 1372 265 1378
rect 586 1378 814 1381
rect 926 1378 958 1381
rect 962 1378 998 1381
rect 1390 1381 1393 1388
rect 1298 1378 1393 1381
rect 1534 1382 1537 1388
rect 1578 1378 1662 1381
rect 50 1368 54 1371
rect 114 1368 118 1371
rect 130 1368 214 1371
rect 450 1368 502 1371
rect 566 1371 569 1378
rect 926 1372 929 1378
rect 566 1368 678 1371
rect 818 1368 926 1371
rect 946 1368 966 1371
rect 970 1368 993 1371
rect 1266 1368 1270 1371
rect 1306 1368 1374 1371
rect 1378 1368 1502 1371
rect 1506 1368 1574 1371
rect 1578 1368 1582 1371
rect 154 1358 158 1361
rect 290 1358 302 1361
rect 330 1358 334 1361
rect 406 1361 409 1368
rect 386 1358 409 1361
rect 446 1362 449 1368
rect 550 1362 553 1368
rect 498 1358 534 1361
rect 578 1358 614 1361
rect 654 1358 734 1361
rect 814 1361 817 1368
rect 990 1362 993 1368
rect 754 1358 817 1361
rect 858 1358 942 1361
rect 1314 1358 1414 1361
rect 1418 1358 1510 1361
rect 1514 1358 1518 1361
rect 1630 1361 1633 1368
rect 1594 1358 1678 1361
rect 654 1352 657 1358
rect -26 1351 -22 1352
rect -26 1348 46 1351
rect 58 1348 118 1351
rect 186 1348 294 1351
rect 402 1348 438 1351
rect 442 1348 470 1351
rect 474 1348 502 1351
rect 546 1348 550 1351
rect 562 1348 574 1351
rect 650 1348 654 1351
rect 706 1348 766 1351
rect 842 1348 886 1351
rect 942 1348 958 1351
rect 974 1351 977 1358
rect 1718 1352 1721 1358
rect 974 1348 1094 1351
rect 1146 1348 1150 1351
rect 1162 1348 1166 1351
rect 1210 1348 1246 1351
rect 1338 1348 1438 1351
rect 1442 1348 1646 1351
rect 1650 1348 1662 1351
rect 182 1342 185 1348
rect 942 1342 945 1348
rect 78 1338 94 1341
rect 274 1338 326 1341
rect 530 1338 550 1341
rect 554 1338 566 1341
rect 610 1338 646 1341
rect 650 1338 694 1341
rect 750 1338 774 1341
rect 850 1338 902 1341
rect 906 1338 918 1341
rect 978 1338 1022 1341
rect 1034 1338 1086 1341
rect 1114 1338 1302 1341
rect 1378 1338 1406 1341
rect 1410 1338 1438 1341
rect 1514 1340 1558 1341
rect 1514 1338 1561 1340
rect 1586 1338 1598 1341
rect 1618 1338 1622 1341
rect 1626 1338 1654 1341
rect 78 1332 81 1338
rect 750 1332 753 1338
rect 1334 1332 1337 1338
rect 1670 1332 1673 1338
rect 210 1328 278 1331
rect 282 1328 302 1331
rect 306 1328 358 1331
rect 394 1328 454 1331
rect 570 1328 638 1331
rect 642 1328 702 1331
rect 882 1328 990 1331
rect 1082 1328 1158 1331
rect 1162 1328 1174 1331
rect 1186 1328 1214 1331
rect 1226 1328 1310 1331
rect 1466 1328 1558 1331
rect 26 1318 158 1321
rect 162 1318 214 1321
rect 258 1318 326 1321
rect 330 1318 390 1321
rect 394 1318 406 1321
rect 410 1318 430 1321
rect 814 1321 817 1328
rect 814 1318 982 1321
rect 986 1318 1166 1321
rect 1170 1318 1198 1321
rect 1202 1318 1270 1321
rect 1294 1318 1342 1321
rect 1426 1318 1566 1321
rect 1570 1318 1614 1321
rect 1658 1318 1662 1321
rect 1294 1312 1297 1318
rect 186 1308 190 1311
rect 194 1308 230 1311
rect 410 1308 742 1311
rect 746 1308 766 1311
rect 778 1308 782 1311
rect 786 1308 814 1311
rect 1250 1308 1294 1311
rect 1314 1308 1470 1311
rect 1474 1308 1630 1311
rect 1112 1303 1114 1307
rect 1118 1303 1121 1307
rect 1126 1303 1128 1307
rect 1158 1302 1161 1308
rect 18 1298 86 1301
rect 1042 1298 1046 1301
rect 1242 1298 1278 1301
rect 1282 1298 1430 1301
rect 1434 1298 1454 1301
rect 1458 1298 1494 1301
rect 1498 1298 1542 1301
rect 1546 1298 1574 1301
rect 1578 1298 1590 1301
rect 66 1288 230 1291
rect 234 1288 510 1291
rect 1018 1288 1041 1291
rect 1038 1282 1041 1288
rect 1294 1288 1302 1291
rect 1386 1288 1414 1291
rect 1418 1288 1550 1291
rect 1562 1288 1582 1291
rect 1586 1288 1670 1291
rect -26 1281 -22 1282
rect -26 1278 -15 1281
rect 106 1278 222 1281
rect 274 1278 398 1281
rect 634 1278 646 1281
rect 690 1278 694 1281
rect 706 1278 734 1281
rect 962 1278 982 1281
rect 1182 1281 1185 1288
rect 1294 1282 1297 1288
rect 1130 1278 1278 1281
rect 1322 1278 1358 1281
rect 1362 1278 1366 1281
rect 1426 1278 1446 1281
rect 1450 1278 1486 1281
rect 1554 1278 1614 1281
rect -18 1271 -15 1278
rect -18 1268 78 1271
rect 82 1268 206 1271
rect 282 1268 286 1271
rect 298 1268 326 1271
rect 662 1271 665 1278
rect 662 1268 710 1271
rect 1006 1271 1009 1278
rect 1006 1268 1046 1271
rect 1106 1268 1110 1271
rect 1118 1271 1121 1278
rect 1118 1268 1662 1271
rect 10 1258 14 1261
rect 214 1261 217 1268
rect 178 1258 217 1261
rect 270 1261 273 1268
rect 270 1258 286 1261
rect 462 1261 465 1268
rect 462 1258 478 1261
rect 526 1261 529 1268
rect 526 1258 542 1261
rect 634 1258 662 1261
rect 690 1258 734 1261
rect 914 1259 918 1261
rect 910 1258 918 1259
rect 994 1258 1126 1261
rect 1138 1258 1198 1261
rect 1206 1258 1214 1261
rect 1218 1258 1222 1261
rect 1234 1258 1238 1261
rect 1266 1258 1310 1261
rect 1354 1258 1358 1261
rect 1538 1258 1558 1261
rect 1610 1258 1622 1261
rect 1670 1261 1673 1268
rect 1666 1258 1673 1261
rect -26 1251 -22 1252
rect -26 1248 6 1251
rect 58 1248 110 1251
rect 218 1248 334 1251
rect 386 1248 390 1251
rect 506 1248 566 1251
rect 570 1248 678 1251
rect 682 1248 726 1251
rect 842 1248 862 1251
rect 866 1248 958 1251
rect 986 1248 1022 1251
rect 1042 1248 1214 1251
rect 1218 1248 1238 1251
rect 1610 1248 1614 1251
rect 86 1242 89 1248
rect 710 1242 713 1248
rect 170 1238 198 1241
rect 290 1238 294 1241
rect 358 1238 382 1241
rect 434 1238 470 1241
rect 594 1238 606 1241
rect 986 1238 1150 1241
rect 1210 1238 1566 1241
rect 1570 1238 1614 1241
rect 358 1232 361 1238
rect 10 1228 206 1231
rect 554 1228 622 1231
rect 722 1228 1046 1231
rect 1050 1228 1262 1231
rect 1346 1228 1398 1231
rect 1402 1228 1446 1231
rect 14 1218 22 1221
rect 138 1218 174 1221
rect 178 1218 262 1221
rect 266 1218 302 1221
rect 306 1218 342 1221
rect 426 1218 582 1221
rect 586 1218 590 1221
rect 1146 1218 1222 1221
rect 1250 1218 1286 1221
rect 1290 1218 1374 1221
rect 14 1212 17 1218
rect 322 1208 414 1211
rect 600 1203 602 1207
rect 606 1203 609 1207
rect 614 1203 616 1207
rect 26 1198 110 1201
rect 202 1188 326 1191
rect 338 1188 342 1191
rect 562 1188 710 1191
rect 714 1188 806 1191
rect 922 1188 950 1191
rect 54 1182 57 1188
rect 114 1178 214 1181
rect 526 1181 529 1188
rect 526 1178 574 1181
rect 706 1178 718 1181
rect 694 1172 697 1178
rect 114 1168 118 1171
rect 306 1168 318 1171
rect 338 1168 374 1171
rect 394 1168 454 1171
rect 490 1168 686 1171
rect 810 1168 902 1171
rect 1498 1168 1518 1171
rect 1522 1168 1526 1171
rect 74 1158 126 1161
rect 146 1158 158 1161
rect 318 1158 430 1161
rect 434 1158 446 1161
rect 482 1158 486 1161
rect 634 1158 654 1161
rect 658 1158 670 1161
rect 674 1158 686 1161
rect 690 1158 734 1161
rect 1242 1158 1278 1161
rect 1282 1158 1302 1161
rect 1306 1158 1358 1161
rect 1470 1161 1473 1168
rect 1394 1158 1473 1161
rect 1582 1161 1585 1168
rect 1522 1158 1585 1161
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 10 1148 166 1151
rect 318 1151 321 1158
rect 710 1152 713 1158
rect 170 1148 321 1151
rect 330 1148 382 1151
rect 410 1148 542 1151
rect 546 1148 614 1151
rect 870 1151 873 1158
rect 870 1148 926 1151
rect 1170 1148 1206 1151
rect 1298 1148 1326 1151
rect 1362 1148 1406 1151
rect 1606 1151 1609 1158
rect 1482 1148 1609 1151
rect 1682 1148 1718 1151
rect 782 1142 785 1148
rect 838 1142 841 1148
rect -26 1138 70 1141
rect 74 1138 310 1141
rect 314 1138 326 1141
rect 446 1138 470 1141
rect 498 1138 502 1141
rect 510 1138 566 1141
rect 1402 1138 1449 1141
rect 1522 1138 1542 1141
rect 1546 1138 1566 1141
rect 1570 1138 1598 1141
rect 1610 1138 1614 1141
rect -26 1132 -23 1138
rect 446 1132 449 1138
rect 510 1132 513 1138
rect 1446 1132 1449 1138
rect -26 1128 -22 1132
rect 18 1128 22 1131
rect 26 1128 38 1131
rect 218 1128 286 1131
rect 522 1128 590 1131
rect 1410 1128 1422 1131
rect 1506 1128 1526 1131
rect 1530 1128 1550 1131
rect 1554 1128 1574 1131
rect 114 1118 134 1121
rect 138 1118 174 1121
rect 178 1118 198 1121
rect 202 1118 238 1121
rect 242 1118 310 1121
rect 394 1118 414 1121
rect 418 1118 486 1121
rect 490 1118 518 1121
rect 802 1118 902 1121
rect 1242 1118 1270 1121
rect 1274 1118 1318 1121
rect 1322 1118 1382 1121
rect 1386 1118 1422 1121
rect 1426 1118 1462 1121
rect 550 1112 553 1118
rect 258 1108 262 1111
rect 274 1108 334 1111
rect 338 1108 342 1111
rect 674 1108 966 1111
rect 978 1108 1030 1111
rect 1698 1108 1710 1111
rect 1112 1103 1114 1107
rect 1118 1103 1121 1107
rect 1126 1103 1128 1107
rect -26 1101 -22 1102
rect -26 1098 6 1101
rect 10 1098 62 1101
rect 82 1098 102 1101
rect 474 1098 641 1101
rect 650 1098 758 1101
rect 810 1098 814 1101
rect 18 1088 206 1091
rect 514 1088 558 1091
rect 638 1091 641 1098
rect 638 1088 670 1091
rect 706 1088 910 1091
rect 1022 1088 1046 1091
rect 1122 1088 1174 1091
rect 278 1082 281 1088
rect 1022 1082 1025 1088
rect -26 1081 -22 1082
rect -26 1078 209 1081
rect 206 1072 209 1078
rect 338 1078 550 1081
rect 626 1078 926 1081
rect 1282 1078 1302 1081
rect 1414 1081 1417 1088
rect 1386 1078 1417 1081
rect 162 1068 198 1071
rect 210 1068 214 1071
rect 222 1071 225 1078
rect 222 1068 246 1071
rect 578 1068 622 1071
rect 714 1068 766 1071
rect 818 1068 822 1071
rect 1074 1068 1230 1071
rect 1370 1068 1390 1071
rect 1394 1068 1398 1071
rect -26 1061 -22 1062
rect -26 1058 14 1061
rect 42 1058 54 1061
rect 94 1061 97 1068
rect 110 1061 113 1068
rect 94 1058 113 1061
rect 122 1058 150 1061
rect 226 1058 278 1061
rect 314 1058 358 1061
rect 394 1058 398 1061
rect 438 1061 441 1068
rect 438 1058 494 1061
rect 542 1061 545 1068
rect 542 1058 550 1061
rect 578 1058 630 1061
rect 650 1058 678 1061
rect 762 1058 838 1061
rect 842 1058 870 1061
rect 894 1061 897 1068
rect 894 1058 910 1061
rect 990 1058 1014 1061
rect 1106 1058 1150 1061
rect 1258 1058 1270 1061
rect 1306 1058 1326 1061
rect 1642 1058 1649 1061
rect 18 1048 57 1051
rect 54 1042 57 1048
rect 378 1048 398 1051
rect 530 1048 542 1051
rect 642 1048 678 1051
rect 758 1051 761 1058
rect 990 1052 993 1058
rect 1166 1052 1169 1058
rect 1646 1052 1649 1058
rect 690 1048 761 1051
rect 810 1048 822 1051
rect 826 1048 926 1051
rect 1010 1048 1070 1051
rect 1194 1048 1302 1051
rect 1378 1048 1390 1051
rect 86 1041 89 1048
rect 74 1038 89 1041
rect 98 1038 142 1041
rect 170 1038 262 1041
rect 266 1038 278 1041
rect 358 1041 361 1048
rect 330 1038 361 1041
rect 482 1038 486 1041
rect 578 1038 582 1041
rect 770 1038 774 1041
rect 850 1038 854 1041
rect 906 1038 913 1041
rect 930 1038 990 1041
rect 1322 1038 1454 1041
rect 1594 1038 1654 1041
rect 910 1032 913 1038
rect 26 1028 30 1031
rect 194 1028 238 1031
rect 506 1028 662 1031
rect 674 1028 790 1031
rect 858 1028 878 1031
rect 970 1028 1086 1031
rect 1338 1028 1374 1031
rect 30 1022 33 1028
rect 66 1018 454 1021
rect 458 1018 630 1021
rect 702 1018 710 1021
rect 714 1018 974 1021
rect 1242 1018 1262 1021
rect 1266 1018 1358 1021
rect 1362 1018 1382 1021
rect 402 1008 574 1011
rect 826 1008 1142 1011
rect 1250 1008 1366 1011
rect 600 1003 602 1007
rect 606 1003 609 1007
rect 614 1003 616 1007
rect 82 998 126 1001
rect 130 998 414 1001
rect 482 998 582 1001
rect 794 998 881 1001
rect 890 998 910 1001
rect 1226 998 1262 1001
rect 370 988 830 991
rect 838 988 846 991
rect 850 988 870 991
rect 878 991 881 998
rect 878 988 1094 991
rect 1270 991 1273 998
rect 1226 988 1273 991
rect 1386 988 1422 991
rect 6 982 9 988
rect 282 978 294 981
rect 418 978 678 981
rect 1674 978 1678 981
rect -26 971 -22 972
rect -26 968 6 971
rect 54 968 102 971
rect 178 968 206 971
rect 290 968 302 971
rect 354 968 358 971
rect 426 968 462 971
rect 530 968 574 971
rect 610 968 694 971
rect 742 971 745 978
rect 722 968 745 971
rect 778 968 814 971
rect 854 971 857 978
rect 842 968 857 971
rect 922 968 1062 971
rect 54 962 57 968
rect 230 961 233 968
rect 478 962 481 968
rect 138 958 238 961
rect 242 958 254 961
rect 338 958 406 961
rect 482 958 558 961
rect 666 958 710 961
rect 754 958 766 961
rect 810 958 838 961
rect 882 958 902 961
rect 1450 958 1510 961
rect -26 951 -22 952
rect -26 948 6 951
rect 10 948 46 951
rect 82 948 134 951
rect 138 948 158 951
rect 162 948 174 951
rect 270 951 273 958
rect 250 948 273 951
rect 286 948 294 951
rect 326 951 329 958
rect 314 948 329 951
rect 370 948 374 951
rect 454 951 457 958
rect 998 952 1001 958
rect 454 948 470 951
rect 558 948 566 951
rect 690 948 742 951
rect 802 948 814 951
rect 866 948 974 951
rect 1026 948 1206 951
rect 286 942 289 948
rect 94 938 118 941
rect 158 938 222 941
rect 330 938 334 941
rect 378 938 422 941
rect 438 941 441 948
rect 558 942 561 948
rect 1402 948 1406 951
rect 1530 948 1558 951
rect 438 938 446 941
rect 450 938 518 941
rect 694 938 702 941
rect 706 938 718 941
rect 1050 938 1054 941
rect 1098 938 1102 941
rect 1162 938 1326 941
rect 1350 941 1353 948
rect 1510 941 1513 948
rect 1526 941 1529 948
rect 1350 938 1529 941
rect 1686 938 1710 941
rect 94 932 97 938
rect 158 932 161 938
rect 10 928 70 931
rect 254 931 257 938
rect 254 928 342 931
rect 498 928 526 931
rect 706 928 710 931
rect 754 928 758 931
rect 762 928 838 931
rect 842 928 862 931
rect 866 928 910 931
rect 914 928 926 931
rect 1042 928 1046 931
rect 1098 928 1134 931
rect 1138 928 1158 931
rect 1394 928 1398 931
rect 1422 928 1518 931
rect 1522 928 1630 931
rect 1686 931 1689 938
rect 1634 928 1689 931
rect 30 922 33 928
rect 1422 922 1425 928
rect 1718 922 1721 928
rect 194 918 622 921
rect 714 918 774 921
rect 866 918 878 921
rect 994 918 998 921
rect 1110 918 1118 921
rect 1122 918 1158 921
rect 1514 918 1630 921
rect 1166 912 1169 918
rect 10 908 142 911
rect 146 908 542 911
rect 730 908 806 911
rect 1458 908 1590 911
rect 1594 908 1638 911
rect 1112 903 1114 907
rect 1118 903 1121 907
rect 1126 903 1128 907
rect -26 901 -22 902
rect -26 898 6 901
rect 10 898 190 901
rect 474 898 494 901
rect 690 898 798 901
rect 1162 898 1254 901
rect 1290 898 1422 901
rect 1466 898 1526 901
rect 1554 898 1710 901
rect 122 888 238 891
rect 778 888 942 891
rect 1186 888 1190 891
rect 1370 888 1406 891
rect 1706 888 1726 891
rect -26 878 -22 882
rect 62 881 65 888
rect 26 878 65 881
rect 122 878 150 881
rect 178 878 190 881
rect 234 878 262 881
rect 314 878 326 881
rect 346 878 358 881
rect 362 878 366 881
rect 386 878 438 881
rect 490 878 518 881
rect 522 878 582 881
rect 586 878 662 881
rect 754 878 934 881
rect 970 878 990 881
rect 1018 878 1038 881
rect 1042 878 1174 881
rect 1586 878 1726 881
rect -26 871 -23 878
rect -26 868 54 871
rect 58 868 78 871
rect 86 871 89 878
rect 86 868 110 871
rect 194 868 198 871
rect 266 868 278 871
rect 282 868 374 871
rect 546 868 582 871
rect 730 868 758 871
rect 826 868 998 871
rect 1138 868 1198 871
rect 1202 868 1230 871
rect 1294 871 1297 878
rect 1234 868 1297 871
rect 1438 871 1441 878
rect 1438 868 1478 871
rect 1586 868 1630 871
rect 1634 868 1670 871
rect -26 861 -22 862
rect -26 858 14 861
rect 42 858 134 861
rect 222 858 225 868
rect 250 858 254 861
rect 266 858 278 861
rect 298 858 302 861
rect 322 858 342 861
rect 414 861 417 868
rect 354 858 417 861
rect 534 861 537 868
rect 1006 862 1009 868
rect 442 858 449 861
rect 534 858 550 861
rect 626 858 718 861
rect 746 858 750 861
rect 786 858 790 861
rect 834 858 838 861
rect 962 858 966 861
rect 1122 858 1294 861
rect 1682 858 1702 861
rect 446 852 449 858
rect 766 852 769 858
rect 814 852 817 858
rect 870 852 873 858
rect 1654 852 1657 858
rect 178 848 182 851
rect 242 848 310 851
rect 394 848 414 851
rect 490 848 494 851
rect 514 848 574 851
rect 578 848 734 851
rect 770 848 790 851
rect 914 848 926 851
rect 954 848 974 851
rect 1122 848 1158 851
rect 1266 848 1350 851
rect 1450 848 1486 851
rect 1758 851 1762 852
rect 1706 848 1762 851
rect 30 841 33 848
rect 110 842 113 848
rect 30 838 94 841
rect 162 838 470 841
rect 498 838 558 841
rect 634 838 678 841
rect 730 838 785 841
rect 850 838 886 841
rect 930 838 950 841
rect 1098 838 1454 841
rect 782 832 785 838
rect -2 828 118 831
rect 194 828 366 831
rect 370 828 518 831
rect 522 828 542 831
rect 594 828 638 831
rect 642 828 654 831
rect 670 828 718 831
rect 866 828 894 831
rect 922 828 926 831
rect 1282 828 1334 831
rect -26 821 -22 822
rect -2 821 1 828
rect 670 822 673 828
rect -26 818 1 821
rect 106 818 134 821
rect 162 818 206 821
rect 378 818 398 821
rect 506 818 646 821
rect 682 818 686 821
rect 698 818 814 821
rect 18 808 70 811
rect 394 808 422 811
rect 1002 808 1470 811
rect 600 803 602 807
rect 606 803 609 807
rect 614 803 616 807
rect -26 801 -22 802
rect -26 798 38 801
rect 42 798 54 801
rect 74 798 326 801
rect 402 798 438 801
rect 466 798 590 801
rect 638 798 750 801
rect 938 798 1438 801
rect 590 788 598 791
rect 638 791 641 798
rect 602 788 641 791
rect 650 788 694 791
rect 706 788 734 791
rect 986 788 998 791
rect 1370 788 1398 791
rect 1666 788 1694 791
rect -26 781 -22 782
rect -26 778 110 781
rect 210 778 758 781
rect 762 778 838 781
rect 954 778 1390 781
rect 1398 772 1401 778
rect 42 768 46 771
rect 74 768 254 771
rect 258 768 414 771
rect 450 768 486 771
rect 562 768 638 771
rect 650 768 654 771
rect 682 768 726 771
rect 938 768 942 771
rect 962 768 974 771
rect 978 768 1006 771
rect 1010 768 1030 771
rect 1122 768 1238 771
rect 1242 768 1398 771
rect -26 761 -22 762
rect -26 758 6 761
rect 10 758 46 761
rect 58 758 158 761
rect 330 758 430 761
rect 434 758 454 761
rect 542 758 550 761
rect 554 758 590 761
rect 618 758 742 761
rect 746 758 806 761
rect 834 758 961 761
rect 970 758 1366 761
rect 1462 761 1465 768
rect 1462 758 1558 761
rect 50 748 54 751
rect 58 748 78 751
rect 146 748 166 751
rect 298 748 358 751
rect 478 751 481 758
rect 958 752 961 758
rect 478 748 494 751
rect 546 748 550 751
rect 578 748 662 751
rect 738 748 750 751
rect 794 748 942 751
rect 986 748 1169 751
rect 1394 748 1518 751
rect 1166 742 1169 748
rect -26 741 -22 742
rect -26 738 54 741
rect 102 738 134 741
rect 138 738 174 741
rect 178 738 230 741
rect 270 738 694 741
rect 698 738 838 741
rect 994 738 1022 741
rect 1434 738 1494 741
rect 1530 738 1534 741
rect 102 732 105 738
rect 270 732 273 738
rect 26 728 46 731
rect 114 728 214 731
rect 218 728 270 731
rect 322 728 334 731
rect 346 728 350 731
rect 466 728 486 731
rect 490 728 526 731
rect 530 728 553 731
rect 594 728 630 731
rect 650 728 686 731
rect 746 728 774 731
rect 786 728 798 731
rect 1034 728 1110 731
rect 1430 731 1433 738
rect 1402 728 1454 731
rect 1482 728 1486 731
rect 550 722 553 728
rect 50 718 150 721
rect 210 718 278 721
rect 290 718 366 721
rect 370 718 542 721
rect 762 718 822 721
rect 1010 718 1166 721
rect 1706 718 1710 721
rect 58 708 102 711
rect 258 708 302 711
rect 466 708 678 711
rect 738 708 854 711
rect 970 708 974 711
rect 1112 703 1114 707
rect 1118 703 1121 707
rect 1126 703 1128 707
rect -26 701 -22 702
rect -26 698 62 701
rect 66 698 190 701
rect 1758 701 1762 702
rect 1698 698 1762 701
rect 146 688 358 691
rect 362 688 422 691
rect 426 688 494 691
rect 546 688 622 691
rect 626 688 686 691
rect 954 688 1014 691
rect 1098 688 1118 691
rect 1426 688 1550 691
rect 1554 688 1582 691
rect -26 681 -22 682
rect -26 678 6 681
rect 82 678 110 681
rect 138 678 214 681
rect 234 678 262 681
rect 282 678 553 681
rect 674 678 718 681
rect 722 678 766 681
rect 778 678 806 681
rect 810 678 894 681
rect 898 678 966 681
rect 970 678 982 681
rect 986 678 1102 681
rect 1210 678 1278 681
rect 1282 678 1334 681
rect 1758 681 1762 682
rect 1738 678 1762 681
rect 78 668 86 671
rect 90 668 94 671
rect 106 668 126 671
rect 426 668 446 671
rect 550 671 553 678
rect 506 668 537 671
rect 550 668 710 671
rect 730 668 934 671
rect 962 668 990 671
rect 1106 668 1150 671
rect 1206 671 1209 678
rect 1186 668 1209 671
rect 1318 668 1422 671
rect 1534 671 1537 678
rect 1534 668 1590 671
rect 42 658 126 661
rect 154 658 158 661
rect 198 661 201 668
rect 178 658 201 661
rect 294 661 297 668
rect 446 662 449 668
rect 534 662 537 668
rect 974 662 977 668
rect 294 658 302 661
rect 550 658 582 661
rect 594 658 926 661
rect 1002 659 1046 661
rect 1286 661 1289 668
rect 1318 662 1321 668
rect 1590 662 1593 668
rect 1002 658 1049 659
rect 1286 658 1302 661
rect 1370 658 1382 661
rect 1474 658 1550 661
rect 1642 658 1662 661
rect 1758 661 1762 662
rect 1666 658 1762 661
rect -26 651 -22 652
rect -26 648 6 651
rect 34 648 38 651
rect 42 648 94 651
rect 98 648 262 651
rect 266 648 294 651
rect 342 651 345 658
rect 322 648 345 651
rect 386 648 390 651
rect 470 651 473 658
rect 394 648 473 651
rect 498 648 502 651
rect 550 651 553 658
rect 526 648 553 651
rect 562 648 782 651
rect 958 651 961 658
rect 958 648 1222 651
rect 1490 648 1606 651
rect 526 642 529 648
rect 10 638 406 641
rect 426 638 462 641
rect 554 638 574 641
rect 586 638 670 641
rect 706 638 814 641
rect 994 638 998 641
rect 1098 638 1110 641
rect 10 628 214 631
rect 218 628 238 631
rect 266 628 310 631
rect 322 628 334 631
rect 346 628 734 631
rect 762 628 974 631
rect 1018 628 1102 631
rect 1758 631 1762 632
rect 1738 628 1762 631
rect 34 618 38 621
rect 50 618 310 621
rect 314 618 334 621
rect 594 618 734 621
rect 802 618 1046 621
rect 122 608 134 611
rect 186 608 238 611
rect 1758 611 1762 612
rect 1666 608 1762 611
rect 600 603 602 607
rect 606 603 609 607
rect 614 603 616 607
rect -26 601 -22 602
rect -26 598 46 601
rect 138 598 342 601
rect 410 598 590 601
rect 626 598 862 601
rect 210 588 230 591
rect 234 588 241 591
rect 250 588 278 591
rect 450 588 454 591
rect 466 588 774 591
rect 1034 588 1342 591
rect 1758 591 1762 592
rect 1570 588 1762 591
rect -26 581 -22 582
rect -26 578 6 581
rect 66 578 86 581
rect 90 578 158 581
rect 162 578 174 581
rect 178 578 198 581
rect 218 578 222 581
rect 230 578 358 581
rect 530 578 670 581
rect 674 578 865 581
rect 1082 578 1094 581
rect 1362 578 1422 581
rect 1434 578 1454 581
rect 1486 581 1489 588
rect 1466 578 1489 581
rect 1514 578 1734 581
rect 38 572 41 578
rect 58 568 126 571
rect 154 568 158 571
rect 230 571 233 578
rect 862 572 865 578
rect 170 568 233 571
rect 274 568 278 571
rect 706 568 710 571
rect 746 568 750 571
rect 866 568 886 571
rect 890 568 958 571
rect 962 568 1022 571
rect 1090 568 1094 571
rect 1178 568 1182 571
rect 1194 568 1510 571
rect 1758 571 1762 572
rect 1586 568 1762 571
rect -26 561 -22 562
rect -26 558 6 561
rect 114 558 182 561
rect 186 558 254 561
rect 350 561 353 568
rect 350 558 366 561
rect 382 561 385 568
rect 382 558 406 561
rect 414 561 417 568
rect 414 558 729 561
rect 738 558 758 561
rect 1106 558 1150 561
rect 1370 558 1374 561
rect 1434 558 1494 561
rect 1554 558 1598 561
rect 1602 558 1609 561
rect 34 548 198 551
rect 202 548 230 551
rect 250 548 262 551
rect 294 551 297 558
rect 282 548 297 551
rect 386 548 390 551
rect 418 548 422 551
rect 578 548 582 551
rect 726 551 729 558
rect 830 551 833 558
rect 726 548 833 551
rect 1162 548 1198 551
rect 1202 548 1222 551
rect 1406 551 1409 558
rect 1406 548 1462 551
rect 1650 548 1654 551
rect 1758 551 1762 552
rect 1738 548 1762 551
rect 638 542 641 548
rect 1630 542 1633 548
rect -26 538 -22 542
rect 26 538 54 541
rect 154 538 174 541
rect 186 538 190 541
rect 266 538 390 541
rect 410 538 494 541
rect 706 538 758 541
rect 786 538 790 541
rect 1090 538 1118 541
rect 1218 538 1230 541
rect 1234 538 1254 541
rect 1258 538 1286 541
rect 1290 538 1350 541
rect 1450 538 1518 541
rect 1690 538 1702 541
rect -26 531 -23 538
rect 1518 532 1521 538
rect -26 528 86 531
rect 90 528 142 531
rect 218 528 326 531
rect 362 528 390 531
rect 394 528 414 531
rect 418 528 438 531
rect 722 528 726 531
rect 954 528 1190 531
rect 1282 528 1286 531
rect 1442 528 1486 531
rect 1578 528 1582 531
rect 1602 528 1694 531
rect 1758 531 1762 532
rect 1702 528 1762 531
rect 1702 522 1705 528
rect 10 518 134 521
rect 154 518 318 521
rect 378 518 758 521
rect 762 518 1334 521
rect 1338 518 1702 521
rect -26 511 -22 512
rect -26 508 54 511
rect 58 508 62 511
rect 250 508 334 511
rect 490 508 798 511
rect 802 508 1102 511
rect 1170 508 1230 511
rect 1266 508 1270 511
rect 1758 511 1762 512
rect 1554 508 1762 511
rect 1112 503 1114 507
rect 1118 503 1121 507
rect 1126 503 1128 507
rect 10 498 70 501
rect 98 498 430 501
rect 650 498 790 501
rect 994 498 1006 501
rect 1010 498 1078 501
rect 1082 498 1102 501
rect 1186 498 1206 501
rect 1290 498 1662 501
rect 78 492 81 498
rect -26 491 -22 492
rect -26 488 14 491
rect 162 488 278 491
rect 502 488 1326 491
rect 1330 488 1566 491
rect 1758 491 1762 492
rect 1738 488 1762 491
rect 502 482 505 488
rect 74 478 102 481
rect 202 478 286 481
rect 386 478 414 481
rect 418 478 438 481
rect 474 478 502 481
rect 730 478 790 481
rect 946 478 950 481
rect 962 478 1206 481
rect 1394 478 1462 481
rect 1710 481 1713 488
rect 1698 478 1713 481
rect 110 472 113 478
rect -26 471 -22 472
rect -26 468 6 471
rect 234 468 270 471
rect 274 468 382 471
rect 410 468 454 471
rect 538 468 614 471
rect 638 471 641 478
rect 638 468 662 471
rect 722 468 750 471
rect 778 468 822 471
rect 826 468 894 471
rect 914 468 918 471
rect 970 468 1022 471
rect 1034 468 1134 471
rect 1218 468 1374 471
rect 1406 468 1422 471
rect 1474 468 1478 471
rect 1482 468 1542 471
rect 1586 468 1630 471
rect 1758 471 1762 472
rect 1730 468 1762 471
rect 38 461 41 468
rect 222 462 225 468
rect 26 458 41 461
rect 106 458 150 461
rect 194 458 214 461
rect 290 458 294 461
rect 442 458 814 461
rect 818 458 830 461
rect 850 458 886 461
rect 890 458 958 461
rect 1010 458 1014 461
rect 1050 458 1086 461
rect 1090 458 1126 461
rect 1190 461 1193 468
rect 1406 462 1409 468
rect 1178 458 1193 461
rect 1242 458 1254 461
rect 1274 458 1281 461
rect 1306 458 1366 461
rect 1370 458 1377 461
rect 1538 458 1550 461
rect 1558 461 1561 468
rect 1558 458 1574 461
rect 1666 458 1678 461
rect -26 451 -22 452
rect 6 451 9 458
rect -26 448 110 451
rect 154 448 158 451
rect 186 448 206 451
rect 210 448 326 451
rect 466 448 470 451
rect 558 448 582 451
rect 610 448 678 451
rect 722 448 830 451
rect 930 448 934 451
rect 970 448 1054 451
rect 1058 448 1070 451
rect 1138 448 1150 451
rect 1154 448 1246 451
rect 1278 451 1281 458
rect 1278 448 1321 451
rect 1370 448 1374 451
rect 1442 448 1446 451
rect 1498 448 1502 451
rect 1514 448 1529 451
rect 1610 448 1614 451
rect 1642 448 1657 451
rect 1686 451 1689 458
rect 1674 448 1689 451
rect 1758 451 1762 452
rect 1706 448 1762 451
rect 558 442 561 448
rect 34 438 78 441
rect 122 438 246 441
rect 322 438 334 441
rect 354 438 446 441
rect 594 438 670 441
rect 706 438 846 441
rect 866 438 902 441
rect 962 438 974 441
rect 1086 441 1089 448
rect 1270 442 1273 448
rect 1318 442 1321 448
rect 1026 438 1089 441
rect 1250 438 1262 441
rect 1346 438 1470 441
rect 1474 438 1510 441
rect 1526 441 1529 448
rect 1654 442 1657 448
rect 1526 438 1622 441
rect 1682 438 1726 441
rect 254 432 257 438
rect 518 428 521 438
rect 530 428 574 431
rect 618 428 654 431
rect 682 428 710 431
rect 746 428 750 431
rect 1114 428 1582 431
rect 1594 428 1646 431
rect 182 421 185 428
rect 50 418 185 421
rect 250 418 305 421
rect 434 418 798 421
rect 802 418 1110 421
rect 1178 418 1254 421
rect 1266 418 1302 421
rect 1418 418 1446 421
rect 1490 418 1502 421
rect 1546 418 1566 421
rect 1618 418 1726 421
rect 302 412 305 418
rect 138 408 294 411
rect 674 408 814 411
rect 898 408 950 411
rect 1066 408 1206 411
rect 1290 408 1446 411
rect 1482 408 1486 411
rect 1530 408 1638 411
rect 600 403 602 407
rect 606 403 609 407
rect 614 403 616 407
rect 154 398 366 401
rect 914 398 1046 401
rect 1106 398 1166 401
rect 1426 398 1478 401
rect 1514 398 1614 401
rect 1626 398 1654 401
rect 10 388 70 391
rect 74 388 126 391
rect 130 388 158 391
rect 162 388 238 391
rect 282 388 622 391
rect 626 388 1358 391
rect 1362 388 1534 391
rect 1626 388 1630 391
rect 178 378 230 381
rect 306 378 398 381
rect 498 378 510 381
rect 514 378 590 381
rect 658 378 686 381
rect 718 378 726 381
rect 854 378 862 381
rect 866 378 974 381
rect 986 378 1094 381
rect 1098 378 1198 381
rect 1202 378 1246 381
rect 1254 378 1382 381
rect 1522 378 1678 381
rect 18 368 22 371
rect 74 368 542 371
rect 546 368 1030 371
rect 1254 371 1257 378
rect 1034 368 1257 371
rect 1338 368 1398 371
rect 1418 368 1422 371
rect 1478 368 1486 371
rect 1558 368 1566 371
rect 1570 368 1614 371
rect 1626 368 1702 371
rect 58 358 166 361
rect 170 358 174 361
rect 186 358 198 361
rect 234 358 286 361
rect 402 358 422 361
rect 442 358 534 361
rect 562 358 630 361
rect 634 358 646 361
rect 666 358 702 361
rect 770 358 822 361
rect 890 358 894 361
rect 978 358 998 361
rect 1026 358 1046 361
rect 1082 358 1086 361
rect 1146 358 1182 361
rect 1186 358 1278 361
rect 1378 358 1526 361
rect 1530 358 1622 361
rect 1634 358 1638 361
rect 1666 358 1702 361
rect 1758 361 1762 362
rect 1730 358 1762 361
rect 214 352 217 358
rect 50 348 70 351
rect 130 348 182 351
rect 234 348 238 351
rect 254 348 286 351
rect 318 351 321 358
rect 306 348 321 351
rect 462 348 478 351
rect 570 348 582 351
rect 618 348 694 351
rect 698 348 750 351
rect 762 348 766 351
rect 786 348 822 351
rect 934 351 937 358
rect 934 348 950 351
rect 1006 351 1009 358
rect 990 348 1009 351
rect 1050 348 1342 351
rect 1394 348 1414 351
rect 1458 348 1502 351
rect 1506 348 1510 351
rect 1514 348 1521 351
rect 1594 348 1614 351
rect 1626 348 1630 351
rect 1666 348 1718 351
rect 110 342 113 348
rect 254 342 257 348
rect 462 342 465 348
rect 990 342 993 348
rect 10 338 54 341
rect 266 338 390 341
rect 490 338 558 341
rect 578 338 582 341
rect 650 338 654 341
rect 738 338 766 341
rect 786 338 830 341
rect 874 338 894 341
rect 898 338 910 341
rect 978 338 985 341
rect 1050 338 1094 341
rect 1158 338 1166 341
rect 1170 338 1182 341
rect 1194 338 1206 341
rect 1330 338 1430 341
rect 1442 338 1542 341
rect 1594 338 1614 341
rect 1254 332 1257 338
rect 18 328 30 331
rect 34 328 222 331
rect 250 328 366 331
rect 386 328 454 331
rect 458 328 534 331
rect 554 328 582 331
rect 682 328 750 331
rect 834 328 838 331
rect 866 328 870 331
rect 1090 328 1230 331
rect 1266 328 1278 331
rect 1322 328 1326 331
rect 1346 328 1366 331
rect 1378 328 1462 331
rect 1678 331 1681 338
rect 1758 331 1762 332
rect 1482 328 1762 331
rect 26 318 46 321
rect 218 318 270 321
rect 338 318 446 321
rect 506 318 510 321
rect 538 318 590 321
rect 746 318 910 321
rect 922 318 1313 321
rect 1370 318 1422 321
rect 1450 318 1470 321
rect 1482 318 1494 321
rect 1506 318 1518 321
rect 18 308 22 311
rect 446 311 449 318
rect 446 308 918 311
rect 986 308 1094 311
rect 1170 308 1174 311
rect 1310 311 1313 318
rect 1310 308 1694 311
rect 1112 303 1114 307
rect 1118 303 1121 307
rect 1126 303 1128 307
rect -26 301 -22 302
rect -26 298 6 301
rect 10 298 502 301
rect 510 298 926 301
rect 930 298 1038 301
rect 1058 298 1102 301
rect 1178 298 1214 301
rect 1282 298 1294 301
rect 1298 298 1358 301
rect 1362 298 1398 301
rect 1402 298 1590 301
rect -26 288 70 291
rect 74 288 78 291
rect 306 288 342 291
rect 346 288 390 291
rect 394 288 406 291
rect 510 291 513 298
rect 414 288 513 291
rect 682 288 758 291
rect 962 288 998 291
rect 1002 288 1110 291
rect 1114 288 1142 291
rect 1250 288 1377 291
rect -26 282 -23 288
rect -26 278 -22 282
rect 42 278 62 281
rect 110 281 113 288
rect 66 278 113 281
rect 302 281 305 288
rect 290 278 305 281
rect 414 281 417 288
rect 330 278 401 281
rect 398 272 401 278
rect 406 278 417 281
rect 506 278 638 281
rect 678 281 681 288
rect 1374 282 1377 288
rect 1690 288 1694 291
rect 642 278 694 281
rect 738 278 814 281
rect 858 278 894 281
rect 898 278 1102 281
rect 1162 278 1198 281
rect 1202 278 1278 281
rect 1566 281 1569 288
rect 1378 278 1489 281
rect 1566 278 1598 281
rect 1602 278 1678 281
rect 1682 278 1710 281
rect 406 272 409 278
rect 234 268 262 271
rect 274 268 278 271
rect 554 268 598 271
rect 602 268 654 271
rect 658 268 678 271
rect 682 268 782 271
rect 786 268 846 271
rect 858 268 862 271
rect 954 268 982 271
rect 1010 268 1014 271
rect 1074 268 1086 271
rect 1102 271 1105 278
rect 1486 272 1489 278
rect 1090 268 1105 271
rect 1154 268 1174 271
rect 1178 268 1262 271
rect 1362 268 1398 271
rect 1490 268 1518 271
rect 1522 268 1534 271
rect 1758 271 1762 272
rect 1698 268 1762 271
rect 110 262 113 268
rect 122 258 190 261
rect 194 258 278 261
rect 282 258 294 261
rect 366 261 369 268
rect 354 258 369 261
rect 502 262 505 268
rect 518 258 526 261
rect 530 258 534 261
rect 554 258 566 261
rect 586 258 614 261
rect 634 258 686 261
rect 690 258 798 261
rect 886 261 889 268
rect 1126 261 1129 268
rect 886 258 1121 261
rect 1126 258 1198 261
rect 1214 258 1222 261
rect 1226 258 1230 261
rect 1302 261 1305 268
rect 1302 258 1318 261
rect 1422 261 1425 268
rect 1422 258 1438 261
rect 1514 258 1526 261
rect 1634 258 1718 261
rect -26 251 -22 252
rect -26 248 102 251
rect 138 248 158 251
rect 226 248 262 251
rect 266 248 318 251
rect 322 248 342 251
rect 458 248 534 251
rect 578 248 606 251
rect 650 248 670 251
rect 754 248 806 251
rect 870 251 873 258
rect 870 248 950 251
rect 1010 248 1078 251
rect 1082 248 1094 251
rect 1118 251 1121 258
rect 1254 252 1257 258
rect 1118 248 1150 251
rect 1162 248 1230 251
rect 1330 248 1350 251
rect 1362 248 1478 251
rect 1502 248 1510 251
rect 1522 248 1622 251
rect 1502 242 1505 248
rect 74 238 78 241
rect 106 238 134 241
rect 146 238 150 241
rect 202 238 254 241
rect 266 238 310 241
rect 506 238 1054 241
rect 1058 238 1198 241
rect 1242 238 1350 241
rect 1394 238 1406 241
rect 1538 238 1590 241
rect 98 228 238 231
rect 250 228 342 231
rect 546 228 566 231
rect 722 228 1134 231
rect 1138 228 1294 231
rect 178 218 270 221
rect 498 218 550 221
rect 594 218 622 221
rect 754 218 766 221
rect 834 218 854 221
rect 902 218 910 221
rect 914 218 942 221
rect 1010 218 1078 221
rect 1090 218 1118 221
rect 1162 218 1166 221
rect 1178 218 1286 221
rect 186 208 238 211
rect 258 208 414 211
rect 698 208 734 211
rect 802 208 1030 211
rect 1034 208 1054 211
rect 1114 208 1246 211
rect 1338 208 1470 211
rect 1474 208 1494 211
rect 1498 208 1614 211
rect 1618 208 1646 211
rect 600 203 602 207
rect 606 203 609 207
rect 614 203 616 207
rect 10 198 78 201
rect 82 198 158 201
rect 866 198 958 201
rect 962 198 974 201
rect 978 198 1321 201
rect 1562 198 1654 201
rect 18 188 54 191
rect 186 188 329 191
rect 418 188 854 191
rect 858 188 878 191
rect 1098 188 1230 191
rect 1318 191 1321 198
rect 1318 188 1518 191
rect 1586 188 1710 191
rect 326 182 329 188
rect -26 181 -22 182
rect -26 178 6 181
rect 26 178 142 181
rect 146 178 206 181
rect 378 178 710 181
rect 714 178 942 181
rect 1010 178 1038 181
rect 1066 178 1134 181
rect 1154 178 1174 181
rect 1310 181 1313 188
rect 1242 178 1313 181
rect 18 168 30 171
rect 66 168 86 171
rect 214 171 217 178
rect 202 168 217 171
rect 226 168 230 171
rect 290 168 302 171
rect 322 168 462 171
rect 586 168 638 171
rect 650 168 670 171
rect 690 168 729 171
rect 738 168 814 171
rect 842 168 854 171
rect 938 168 974 171
rect 1010 168 1014 171
rect 1130 168 1222 171
rect 1438 171 1441 178
rect 1274 168 1441 171
rect 1514 168 1590 171
rect 726 162 729 168
rect -26 161 -22 162
rect -26 158 22 161
rect 126 158 166 161
rect 170 158 174 161
rect 210 158 238 161
rect 394 158 542 161
rect 546 158 702 161
rect 714 158 718 161
rect 806 158 822 161
rect 878 161 881 168
rect 858 158 881 161
rect 1026 158 1046 161
rect 1050 158 1150 161
rect 1170 158 1193 161
rect 1250 158 1270 161
rect 1370 158 1414 161
rect 1530 158 1534 161
rect 1546 158 1574 161
rect 1602 158 1638 161
rect 62 151 65 158
rect 58 148 65 151
rect 126 152 129 158
rect 186 148 190 151
rect 282 148 321 151
rect 350 151 353 158
rect 338 148 353 151
rect 382 151 385 158
rect 806 152 809 158
rect 370 148 385 151
rect 390 148 417 151
rect 238 142 241 148
rect 50 138 110 141
rect 162 138 230 141
rect 250 138 270 141
rect 318 141 321 148
rect 390 141 393 148
rect 414 142 417 148
rect 522 148 529 151
rect 578 148 662 151
rect 698 148 734 151
rect 762 148 782 151
rect 818 148 910 151
rect 942 151 945 158
rect 930 148 945 151
rect 1042 148 1078 151
rect 1158 151 1161 158
rect 1190 152 1193 158
rect 1106 148 1161 151
rect 1170 148 1174 151
rect 1202 148 1278 151
rect 1282 148 1286 151
rect 1342 151 1345 158
rect 1298 148 1345 151
rect 1502 151 1505 158
rect 1498 148 1505 151
rect 1514 148 1542 151
rect 1578 148 1582 151
rect 1626 148 1630 151
rect 1758 151 1762 152
rect 1690 148 1762 151
rect 318 138 393 141
rect 402 138 406 141
rect 434 138 438 141
rect 446 141 449 148
rect 478 141 481 148
rect 526 142 529 148
rect 446 138 481 141
rect 506 138 518 141
rect 626 138 1345 141
rect 1354 138 1358 141
rect 1386 138 1406 141
rect 1482 138 1598 141
rect 1666 138 1697 141
rect 106 128 174 131
rect 310 131 313 138
rect 310 128 366 131
rect 370 128 398 131
rect 402 128 414 131
rect 418 128 430 131
rect 434 128 454 131
rect 490 128 614 131
rect 746 128 758 131
rect 770 128 790 131
rect 890 128 894 131
rect 914 128 1086 131
rect 1098 128 1126 131
rect 1154 128 1158 131
rect 1202 128 1206 131
rect 1322 128 1326 131
rect 1342 131 1345 138
rect 1694 132 1697 138
rect 1342 128 1454 131
rect 1458 128 1678 131
rect 498 118 598 121
rect 602 118 702 121
rect 730 118 830 121
rect 850 118 854 121
rect 882 118 1006 121
rect 1042 118 1062 121
rect 1074 118 1190 121
rect 1194 118 1230 121
rect 1302 121 1305 128
rect 1250 118 1334 121
rect 1338 118 1366 121
rect 1370 118 1438 121
rect 1514 118 1566 121
rect 1594 118 1678 121
rect 346 108 670 111
rect 850 108 902 111
rect 906 108 966 111
rect 1186 108 1198 111
rect 1202 108 1214 111
rect 1242 108 1358 111
rect 1370 108 1406 111
rect 1418 108 1534 111
rect 1546 108 1622 111
rect 1112 103 1114 107
rect 1118 103 1121 107
rect 1126 103 1128 107
rect 122 98 142 101
rect 146 98 774 101
rect 778 98 958 101
rect 1138 98 1374 101
rect 1386 98 1398 101
rect 1402 98 1422 101
rect 1426 98 1526 101
rect 1530 98 1550 101
rect 1554 98 1670 101
rect 170 88 654 91
rect 658 88 798 91
rect 994 88 1030 91
rect 1034 88 1046 91
rect 1050 88 1102 91
rect 1106 88 1198 91
rect 1338 88 1382 91
rect 1466 88 1486 91
rect 1490 88 1518 91
rect 1522 88 1550 91
rect 1554 88 1662 91
rect 26 78 46 81
rect 126 81 129 88
rect 90 78 129 81
rect 318 78 326 81
rect 330 78 537 81
rect 546 78 550 81
rect 554 78 582 81
rect 586 78 606 81
rect 610 78 702 81
rect 714 78 750 81
rect 806 81 809 88
rect 854 82 857 88
rect 754 78 846 81
rect 962 78 966 81
rect 1058 78 1062 81
rect 1074 78 1078 81
rect 1082 78 1134 81
rect 1286 81 1289 88
rect 1138 78 1289 81
rect 1330 78 1526 81
rect 1578 78 1606 81
rect 18 68 38 71
rect 42 68 86 71
rect 202 68 206 71
rect 226 68 254 71
rect 258 68 278 71
rect 282 68 318 71
rect 322 68 342 71
rect 346 68 358 71
rect 378 68 422 71
rect 426 68 433 71
rect 442 68 478 71
rect 534 71 537 78
rect 534 68 742 71
rect 746 68 798 71
rect 810 68 814 71
rect 842 68 846 71
rect 890 68 926 71
rect 998 71 1001 78
rect 1662 72 1665 78
rect 970 68 1001 71
rect 1090 68 1118 71
rect 1170 68 1230 71
rect 1234 68 1246 71
rect 1338 68 1342 71
rect 1354 68 1494 71
rect 1674 68 1686 71
rect 1706 70 1713 71
rect 1706 68 1710 70
rect 26 58 158 61
rect 210 58 294 61
rect 394 58 558 61
rect 562 58 662 61
rect 682 58 782 61
rect 986 58 1006 61
rect 1050 58 1142 61
rect 1146 58 1214 61
rect 1298 58 1358 61
rect 1402 58 1406 61
rect 1698 58 1734 61
rect 1758 61 1762 62
rect 1738 58 1762 61
rect 42 48 70 51
rect 346 48 350 51
rect 426 48 438 51
rect 458 48 470 51
rect 782 51 785 58
rect 478 48 569 51
rect 782 48 1278 51
rect 1282 48 1430 51
rect 414 41 417 48
rect 178 38 417 41
rect 478 42 481 48
rect 566 42 569 48
rect 570 38 1238 41
rect 1242 38 1262 41
rect 1266 38 1470 41
rect 442 28 510 31
rect 514 28 614 31
rect 922 28 1302 31
rect 1314 28 1374 31
rect 282 18 454 21
rect 466 18 686 21
rect 690 18 950 21
rect 954 18 958 21
rect 1026 18 1038 21
rect 1066 18 1078 21
rect 1098 18 1102 21
rect 1210 18 1558 21
rect 50 8 54 11
rect 138 8 158 11
rect 162 8 502 11
rect 754 8 790 11
rect 802 8 814 11
rect 914 8 918 11
rect 978 8 982 11
rect 1058 8 1062 11
rect 1082 8 1166 11
rect 1178 8 1214 11
rect 1226 8 1238 11
rect 1242 8 1286 11
rect 1330 8 1350 11
rect 600 3 602 7
rect 606 3 609 7
rect 614 3 616 7
<< m4contact >>
rect 446 1608 450 1612
rect 622 1608 626 1612
rect 1238 1608 1242 1612
rect 602 1603 606 1607
rect 610 1603 613 1607
rect 613 1603 614 1607
rect 694 1598 698 1602
rect 678 1578 682 1582
rect 1550 1558 1554 1562
rect 1230 1548 1234 1552
rect 1318 1548 1322 1552
rect 182 1538 186 1542
rect 190 1538 194 1542
rect 366 1538 370 1542
rect 478 1538 482 1542
rect 1094 1538 1098 1542
rect 1414 1538 1418 1542
rect 982 1528 986 1532
rect 1310 1528 1314 1532
rect 366 1518 370 1522
rect 550 1518 554 1522
rect 742 1518 746 1522
rect 870 1518 874 1522
rect 966 1518 970 1522
rect 1038 1518 1042 1522
rect 1062 1508 1066 1512
rect 1114 1503 1118 1507
rect 1122 1503 1125 1507
rect 1125 1503 1126 1507
rect 1190 1498 1194 1502
rect 70 1488 74 1492
rect 366 1488 370 1492
rect 54 1468 58 1472
rect 1318 1468 1322 1472
rect 1654 1468 1658 1472
rect 478 1448 482 1452
rect 1190 1448 1194 1452
rect 1662 1448 1666 1452
rect 62 1438 66 1442
rect 630 1438 634 1442
rect 1062 1438 1066 1442
rect 1230 1438 1234 1442
rect 62 1428 66 1432
rect 1646 1428 1650 1432
rect 602 1403 606 1407
rect 610 1403 613 1407
rect 613 1403 614 1407
rect 814 1378 818 1382
rect 1662 1378 1666 1382
rect 54 1368 58 1372
rect 1262 1368 1266 1372
rect 1302 1368 1306 1372
rect 1582 1368 1586 1372
rect 446 1358 450 1362
rect 534 1358 538 1362
rect 550 1358 554 1362
rect 574 1358 578 1362
rect 1518 1358 1522 1362
rect 1718 1358 1722 1362
rect 46 1348 50 1352
rect 550 1348 554 1352
rect 646 1348 650 1352
rect 766 1348 770 1352
rect 958 1348 962 1352
rect 1142 1348 1146 1352
rect 1158 1348 1162 1352
rect 182 1338 186 1342
rect 270 1338 274 1342
rect 694 1338 698 1342
rect 1334 1338 1338 1342
rect 1614 1338 1618 1342
rect 1214 1328 1218 1332
rect 1558 1328 1562 1332
rect 1670 1328 1674 1332
rect 1654 1318 1658 1322
rect 190 1308 194 1312
rect 742 1308 746 1312
rect 774 1308 778 1312
rect 1158 1308 1162 1312
rect 1114 1303 1118 1307
rect 1122 1303 1125 1307
rect 1125 1303 1126 1307
rect 1046 1298 1050 1302
rect 62 1288 66 1292
rect 1302 1288 1306 1292
rect 1558 1288 1562 1292
rect 1670 1288 1674 1292
rect 630 1278 634 1282
rect 694 1278 698 1282
rect 982 1278 986 1282
rect 1126 1278 1130 1282
rect 1358 1278 1362 1282
rect 278 1268 282 1272
rect 1110 1268 1114 1272
rect 6 1258 10 1262
rect 918 1258 922 1262
rect 1126 1258 1130 1262
rect 1134 1258 1138 1262
rect 1222 1258 1226 1262
rect 1238 1258 1242 1262
rect 1262 1258 1266 1262
rect 1662 1258 1666 1262
rect 1038 1248 1042 1252
rect 1614 1248 1618 1252
rect 286 1238 290 1242
rect 982 1238 986 1242
rect 22 1218 26 1222
rect 590 1218 594 1222
rect 602 1203 606 1207
rect 610 1203 613 1207
rect 613 1203 614 1207
rect 110 1198 114 1202
rect 326 1188 330 1192
rect 342 1188 346 1192
rect 710 1188 714 1192
rect 54 1178 58 1182
rect 214 1178 218 1182
rect 686 1168 690 1172
rect 694 1168 698 1172
rect 158 1158 162 1162
rect 478 1158 482 1162
rect 654 1158 658 1162
rect 670 1158 674 1162
rect 542 1148 546 1152
rect 782 1148 786 1152
rect 838 1148 842 1152
rect 494 1138 498 1142
rect 1606 1138 1610 1142
rect 286 1128 290 1132
rect 902 1118 906 1122
rect 1462 1118 1466 1122
rect 262 1108 266 1112
rect 334 1108 338 1112
rect 550 1108 554 1112
rect 966 1108 970 1112
rect 1114 1103 1118 1107
rect 1122 1103 1125 1107
rect 1125 1103 1126 1107
rect 758 1098 762 1102
rect 806 1098 810 1102
rect 910 1088 914 1092
rect 278 1078 282 1082
rect 550 1078 554 1082
rect 926 1078 930 1082
rect 198 1068 202 1072
rect 206 1068 210 1072
rect 814 1068 818 1072
rect 1390 1068 1394 1072
rect 398 1058 402 1062
rect 1014 1058 1018 1062
rect 1150 1058 1154 1062
rect 1166 1058 1170 1062
rect 1638 1058 1642 1062
rect 542 1048 546 1052
rect 678 1048 682 1052
rect 326 1038 330 1042
rect 766 1038 770 1042
rect 854 1038 858 1042
rect 902 1038 906 1042
rect 22 1028 26 1032
rect 30 1018 34 1022
rect 1358 1018 1362 1022
rect 574 1008 578 1012
rect 602 1003 606 1007
rect 610 1003 613 1007
rect 613 1003 614 1007
rect 78 998 82 1002
rect 582 998 586 1002
rect 6 988 10 992
rect 830 988 834 992
rect 1222 988 1226 992
rect 278 978 282 982
rect 1670 978 1674 982
rect 6 968 10 972
rect 478 968 482 972
rect 774 968 778 972
rect 238 958 242 962
rect 334 958 338 962
rect 766 958 770 962
rect 46 948 50 952
rect 294 948 298 952
rect 374 948 378 952
rect 686 948 690 952
rect 998 948 1002 952
rect 326 938 330 942
rect 422 938 426 942
rect 1406 948 1410 952
rect 446 938 450 942
rect 1046 938 1050 942
rect 1102 938 1106 942
rect 6 928 10 932
rect 70 928 74 932
rect 494 928 498 932
rect 710 928 714 932
rect 750 928 754 932
rect 1038 928 1042 932
rect 1390 928 1394 932
rect 1518 928 1522 932
rect 1630 928 1634 932
rect 1718 928 1722 932
rect 998 918 1002 922
rect 1158 918 1162 922
rect 1166 918 1170 922
rect 6 908 10 912
rect 542 908 546 912
rect 1638 908 1642 912
rect 1114 903 1118 907
rect 1122 903 1125 907
rect 1125 903 1126 907
rect 686 898 690 902
rect 1158 898 1162 902
rect 1462 898 1466 902
rect 1550 898 1554 902
rect 1702 888 1706 892
rect 326 878 330 882
rect 966 878 970 882
rect 1014 878 1018 882
rect 1582 878 1586 882
rect 78 868 82 872
rect 190 868 194 872
rect 222 868 226 872
rect 278 868 282 872
rect 542 868 546 872
rect 1582 868 1586 872
rect 14 858 18 862
rect 246 858 250 862
rect 262 858 266 862
rect 294 858 298 862
rect 350 858 354 862
rect 438 858 442 862
rect 750 858 754 862
rect 790 858 794 862
rect 814 858 818 862
rect 838 858 842 862
rect 870 858 874 862
rect 966 858 970 862
rect 1006 858 1010 862
rect 1654 858 1658 862
rect 110 848 114 852
rect 238 848 242 852
rect 766 848 770 852
rect 910 848 914 852
rect 926 838 930 842
rect 190 828 194 832
rect 590 828 594 832
rect 918 828 922 832
rect 646 818 650 822
rect 678 818 682 822
rect 814 818 818 822
rect 14 808 18 812
rect 602 803 606 807
rect 610 803 613 807
rect 613 803 614 807
rect 54 798 58 802
rect 590 798 594 802
rect 694 788 698 792
rect 1390 778 1394 782
rect 1398 778 1402 782
rect 38 768 42 772
rect 70 768 74 772
rect 654 768 658 772
rect 942 768 946 772
rect 1030 768 1034 772
rect 1238 768 1242 772
rect 6 758 10 762
rect 54 758 58 762
rect 830 758 834 762
rect 46 748 50 752
rect 550 748 554 752
rect 1390 748 1394 752
rect 54 738 58 742
rect 1534 738 1538 742
rect 342 728 346 732
rect 742 728 746 732
rect 782 728 786 732
rect 1486 728 1490 732
rect 206 718 210 722
rect 286 718 290 722
rect 542 718 546 722
rect 678 708 682 712
rect 966 708 970 712
rect 1114 703 1118 707
rect 1122 703 1125 707
rect 1125 703 1126 707
rect 190 698 194 702
rect 142 688 146 692
rect 542 688 546 692
rect 686 688 690 692
rect 1094 688 1098 692
rect 1582 688 1586 692
rect 6 678 10 682
rect 1590 668 1594 672
rect 150 658 154 662
rect 446 658 450 662
rect 590 658 594 662
rect 1638 658 1642 662
rect 1662 658 1666 662
rect 30 648 34 652
rect 390 648 394 652
rect 6 638 10 642
rect 670 638 674 642
rect 990 638 994 642
rect 238 628 242 632
rect 262 628 266 632
rect 342 628 346 632
rect 974 628 978 632
rect 1102 628 1106 632
rect 46 618 50 622
rect 334 618 338 622
rect 1046 618 1050 622
rect 182 608 186 612
rect 602 603 606 607
rect 610 603 613 607
rect 613 603 614 607
rect 46 598 50 602
rect 342 598 346 602
rect 622 598 626 602
rect 446 588 450 592
rect 1030 588 1034 592
rect 6 578 10 582
rect 38 578 42 582
rect 222 578 226 582
rect 1734 578 1738 582
rect 126 568 130 572
rect 158 568 162 572
rect 278 568 282 572
rect 702 568 706 572
rect 750 568 754 572
rect 1094 568 1098 572
rect 1174 568 1178 572
rect 1582 568 1586 572
rect 6 558 10 562
rect 110 558 114 562
rect 366 558 370 562
rect 406 558 410 562
rect 1374 558 1378 562
rect 262 548 266 552
rect 390 548 394 552
rect 422 548 426 552
rect 582 548 586 552
rect 638 548 642 552
rect 1198 548 1202 552
rect 1654 548 1658 552
rect 1734 548 1738 552
rect 190 538 194 542
rect 406 538 410 542
rect 790 538 794 542
rect 1518 538 1522 542
rect 1630 538 1634 542
rect 1686 538 1690 542
rect 142 528 146 532
rect 718 528 722 532
rect 1286 528 1290 532
rect 1582 528 1586 532
rect 6 518 10 522
rect 62 508 66 512
rect 246 508 250 512
rect 1102 508 1106 512
rect 1270 508 1274 512
rect 1550 508 1554 512
rect 1114 503 1118 507
rect 1122 503 1125 507
rect 1125 503 1126 507
rect 6 498 10 502
rect 78 498 82 502
rect 14 488 18 492
rect 278 488 282 492
rect 1734 488 1738 492
rect 958 478 962 482
rect 6 468 10 472
rect 110 468 114 472
rect 222 468 226 472
rect 910 468 914 472
rect 1726 468 1730 472
rect 294 458 298 462
rect 830 458 834 462
rect 846 458 850 462
rect 958 458 962 462
rect 1254 458 1258 462
rect 1550 458 1554 462
rect 110 448 114 452
rect 966 448 970 452
rect 1070 448 1074 452
rect 1366 448 1370 452
rect 1446 448 1450 452
rect 1502 448 1506 452
rect 1614 448 1618 452
rect 246 438 250 442
rect 254 438 258 442
rect 518 438 522 442
rect 1270 438 1274 442
rect 1622 438 1626 442
rect 1726 438 1730 442
rect 614 428 618 432
rect 710 428 714 432
rect 750 428 754 432
rect 1582 428 1586 432
rect 1174 418 1178 422
rect 1262 418 1266 422
rect 1726 418 1730 422
rect 1446 408 1450 412
rect 1478 408 1482 412
rect 1526 408 1530 412
rect 602 403 606 407
rect 610 403 613 407
rect 613 403 614 407
rect 1422 398 1426 402
rect 1622 398 1626 402
rect 6 388 10 392
rect 1622 388 1626 392
rect 726 378 730 382
rect 1518 378 1522 382
rect 14 368 18 372
rect 70 368 74 372
rect 1614 368 1618 372
rect 174 358 178 362
rect 214 358 218 362
rect 1078 358 1082 362
rect 1638 358 1642 362
rect 1726 358 1730 362
rect 230 348 234 352
rect 302 348 306 352
rect 582 348 586 352
rect 750 348 754 352
rect 758 348 762 352
rect 782 348 786 352
rect 1502 348 1506 352
rect 1622 348 1626 352
rect 110 338 114 342
rect 262 338 266 342
rect 582 338 586 342
rect 654 338 658 342
rect 974 338 978 342
rect 1046 338 1050 342
rect 1590 338 1594 342
rect 534 328 538 332
rect 830 328 834 332
rect 870 328 874 332
rect 1254 328 1258 332
rect 1262 328 1266 332
rect 1326 328 1330 332
rect 1478 328 1482 332
rect 510 318 514 322
rect 1422 318 1426 322
rect 14 308 18 312
rect 1094 308 1098 312
rect 1166 308 1170 312
rect 1114 303 1118 307
rect 1122 303 1125 307
rect 1125 303 1126 307
rect 502 298 506 302
rect 1102 298 1106 302
rect 78 288 82 292
rect 1694 288 1698 292
rect 110 268 114 272
rect 262 268 266 272
rect 270 268 274 272
rect 502 268 506 272
rect 862 268 866 272
rect 1014 268 1018 272
rect 1086 268 1090 272
rect 1358 268 1362 272
rect 1518 268 1522 272
rect 550 258 554 262
rect 1198 258 1202 262
rect 1254 258 1258 262
rect 646 248 650 252
rect 750 248 754 252
rect 1094 248 1098 252
rect 1510 248 1514 252
rect 150 238 154 242
rect 254 238 258 242
rect 262 238 266 242
rect 502 238 506 242
rect 246 228 250 232
rect 718 228 722 232
rect 550 218 554 222
rect 1006 218 1010 222
rect 1158 218 1162 222
rect 1174 218 1178 222
rect 798 208 802 212
rect 1054 208 1058 212
rect 602 203 606 207
rect 610 203 613 207
rect 613 203 614 207
rect 6 198 10 202
rect 158 198 162 202
rect 974 198 978 202
rect 182 188 186 192
rect 854 188 858 192
rect 6 178 10 182
rect 942 178 946 182
rect 230 168 234 172
rect 318 168 322 172
rect 1006 168 1010 172
rect 166 158 170 162
rect 702 158 706 162
rect 718 158 722 162
rect 1366 158 1370 162
rect 1534 158 1538 162
rect 182 148 186 152
rect 238 148 242 152
rect 366 148 370 152
rect 1166 148 1170 152
rect 1198 148 1202 152
rect 1286 148 1290 152
rect 1510 148 1514 152
rect 1622 148 1626 152
rect 406 138 410 142
rect 438 138 442 142
rect 1358 138 1362 142
rect 766 128 770 132
rect 886 128 890 132
rect 1158 128 1162 132
rect 1198 128 1202 132
rect 1318 128 1322 132
rect 702 118 706 122
rect 846 118 850 122
rect 1006 118 1010 122
rect 1070 118 1074 122
rect 1230 118 1234 122
rect 1510 118 1514 122
rect 1678 118 1682 122
rect 342 108 346 112
rect 1358 108 1362 112
rect 1406 108 1410 112
rect 1534 108 1538 112
rect 1114 103 1118 107
rect 1122 103 1125 107
rect 1125 103 1126 107
rect 958 98 962 102
rect 1134 98 1138 102
rect 798 88 802 92
rect 854 78 858 82
rect 958 78 962 82
rect 1062 78 1066 82
rect 1070 78 1074 82
rect 1606 78 1610 82
rect 438 68 442 72
rect 798 68 802 72
rect 806 68 810 72
rect 846 68 850 72
rect 1086 68 1090 72
rect 1334 68 1338 72
rect 1662 68 1666 72
rect 1670 68 1674 72
rect 1702 68 1706 72
rect 662 58 666 62
rect 1046 58 1050 62
rect 1214 58 1218 62
rect 1398 58 1402 62
rect 342 48 346 52
rect 438 48 442 52
rect 470 48 474 52
rect 614 28 618 32
rect 1310 28 1314 32
rect 462 18 466 22
rect 958 18 962 22
rect 1062 18 1066 22
rect 1094 18 1098 22
rect 1206 18 1210 22
rect 54 8 58 12
rect 502 8 506 12
rect 750 8 754 12
rect 910 8 914 12
rect 974 8 978 12
rect 1054 8 1058 12
rect 1078 8 1082 12
rect 1286 8 1290 12
rect 1350 8 1354 12
rect 602 3 606 7
rect 610 3 613 7
rect 613 3 614 7
<< metal4 >>
rect 626 1608 633 1611
rect 370 1538 374 1541
rect 54 1372 57 1468
rect 70 1441 73 1488
rect 66 1438 73 1441
rect 46 1342 49 1348
rect 62 1292 65 1428
rect 182 1342 185 1538
rect 190 1312 193 1538
rect 366 1492 369 1518
rect 446 1362 449 1608
rect 600 1603 602 1607
rect 606 1603 609 1607
rect 614 1603 616 1607
rect 474 1538 478 1541
rect 266 1338 270 1341
rect 282 1268 289 1271
rect 6 992 9 1258
rect 286 1242 289 1268
rect 22 1032 25 1218
rect 6 932 9 968
rect 6 762 9 908
rect 14 812 17 858
rect 6 642 9 678
rect 30 652 33 1018
rect 38 582 41 768
rect 46 752 49 948
rect 54 802 57 1178
rect 54 742 57 758
rect 46 602 49 618
rect 10 578 14 581
rect 6 522 9 558
rect 62 512 65 1108
rect 70 772 73 928
rect 78 872 81 998
rect 110 852 113 1198
rect 334 1188 342 1191
rect 78 502 81 578
rect 110 562 113 848
rect 130 568 134 571
rect 6 472 9 498
rect 6 392 9 468
rect 14 462 17 488
rect 110 472 113 558
rect 142 532 145 688
rect 158 661 161 1158
rect 198 1062 201 1068
rect 194 868 198 871
rect 190 702 193 828
rect 206 722 209 1068
rect 154 658 161 661
rect 158 552 161 568
rect 182 541 185 608
rect 214 581 217 1178
rect 258 1108 262 1111
rect 278 982 281 1078
rect 222 862 225 868
rect 238 852 241 958
rect 278 872 281 978
rect 258 858 262 861
rect 246 852 249 858
rect 286 722 289 1128
rect 326 1042 329 1188
rect 334 1112 337 1188
rect 478 1162 481 1448
rect 550 1362 553 1518
rect 630 1442 633 1608
rect 670 1578 678 1581
rect 600 1403 602 1407
rect 606 1403 609 1407
rect 614 1403 616 1407
rect 538 1358 542 1361
rect 570 1358 574 1361
rect 542 1348 550 1351
rect 334 962 337 1108
rect 394 1058 398 1061
rect 478 972 481 1158
rect 542 1152 545 1348
rect 630 1282 633 1438
rect 650 1348 657 1351
rect 654 1342 657 1348
rect 494 1112 497 1138
rect 298 948 302 951
rect 370 948 374 951
rect 330 938 337 941
rect 426 938 430 941
rect 302 861 305 868
rect 298 858 305 861
rect 326 862 329 878
rect 334 732 337 938
rect 346 858 350 861
rect 438 852 441 858
rect 238 632 241 648
rect 214 578 222 581
rect 262 552 265 628
rect 334 622 337 728
rect 342 632 345 728
rect 446 662 449 938
rect 494 932 497 1108
rect 550 1082 553 1108
rect 542 912 545 1048
rect 542 872 545 908
rect 550 752 553 1078
rect 574 952 577 1008
rect 582 1002 585 1038
rect 590 832 593 1218
rect 600 1203 602 1207
rect 606 1203 609 1207
rect 614 1203 616 1207
rect 670 1162 673 1578
rect 694 1342 697 1598
rect 970 1518 974 1521
rect 742 1312 745 1518
rect 694 1172 697 1278
rect 600 1003 602 1007
rect 606 1003 609 1007
rect 614 1003 616 1007
rect 646 822 649 848
rect 600 803 602 807
rect 606 803 609 807
rect 614 803 616 807
rect 542 692 545 718
rect 386 648 390 651
rect 342 602 345 628
rect 450 588 454 591
rect 550 582 553 748
rect 590 662 593 798
rect 654 772 657 1158
rect 678 1052 681 1068
rect 686 952 689 1168
rect 710 932 713 1188
rect 758 931 761 1098
rect 766 1042 769 1348
rect 774 972 777 1308
rect 754 928 761 931
rect 670 642 673 868
rect 678 712 681 818
rect 686 692 689 898
rect 754 858 758 861
rect 766 852 769 958
rect 694 772 697 788
rect 782 732 785 1148
rect 814 1101 817 1378
rect 810 1098 817 1101
rect 810 1068 814 1071
rect 790 852 793 858
rect 814 822 817 858
rect 830 762 833 988
rect 838 862 841 1148
rect 850 1038 854 1041
rect 870 862 873 1518
rect 962 1348 966 1351
rect 982 1282 985 1528
rect 1042 1518 1046 1521
rect 1062 1442 1065 1508
rect 1038 1298 1046 1301
rect 902 1042 905 1118
rect 910 852 913 1088
rect 918 832 921 1258
rect 982 1242 985 1278
rect 1038 1252 1041 1298
rect 926 842 929 1078
rect 966 882 969 1108
rect 994 948 998 951
rect 990 918 998 921
rect 962 858 966 861
rect 938 768 942 771
rect 738 728 742 731
rect 970 708 977 711
rect 974 632 977 708
rect 990 642 993 918
rect 1014 882 1017 1058
rect 1050 938 1054 941
rect 1042 928 1049 931
rect 1006 862 1009 868
rect 600 603 602 607
rect 606 603 609 607
rect 614 603 616 607
rect 622 592 625 598
rect 1030 592 1033 768
rect 1046 622 1049 928
rect 1094 692 1097 1538
rect 1112 1503 1114 1507
rect 1118 1503 1121 1507
rect 1126 1503 1128 1507
rect 1190 1452 1193 1498
rect 1230 1442 1233 1548
rect 1146 1348 1150 1351
rect 1158 1312 1161 1348
rect 1214 1332 1217 1338
rect 1112 1303 1114 1307
rect 1118 1303 1121 1307
rect 1126 1303 1128 1307
rect 1106 1268 1110 1271
rect 1126 1262 1129 1278
rect 1134 1262 1137 1268
rect 1238 1262 1241 1608
rect 1310 1532 1313 1538
rect 1318 1472 1321 1548
rect 1418 1538 1422 1541
rect 1262 1262 1265 1368
rect 1302 1292 1305 1368
rect 1330 1338 1334 1341
rect 1112 1103 1114 1107
rect 1118 1103 1121 1107
rect 1126 1103 1128 1107
rect 1154 1058 1158 1061
rect 1102 632 1105 938
rect 1166 922 1169 1058
rect 1222 992 1225 1258
rect 1112 903 1114 907
rect 1118 903 1121 907
rect 1126 903 1128 907
rect 1158 902 1161 918
rect 1238 772 1241 1258
rect 1358 1022 1361 1278
rect 1390 932 1393 1068
rect 1398 948 1406 951
rect 1398 782 1401 948
rect 1462 902 1465 1118
rect 1518 932 1521 1358
rect 1550 902 1553 1558
rect 1558 1292 1561 1328
rect 1582 882 1585 1368
rect 1614 1252 1617 1338
rect 1390 752 1393 778
rect 1526 738 1534 741
rect 1478 728 1486 731
rect 1112 703 1114 707
rect 1118 703 1121 707
rect 1126 703 1128 707
rect 706 568 713 571
rect 182 538 190 541
rect 110 452 113 468
rect 222 462 225 468
rect 246 442 249 508
rect 278 492 281 568
rect 370 558 374 561
rect 386 548 390 551
rect 406 542 409 558
rect 422 552 425 568
rect 638 552 641 558
rect 286 461 289 468
rect 286 458 294 461
rect 14 312 17 368
rect 70 291 73 368
rect 166 358 174 361
rect 218 358 222 361
rect 70 288 78 291
rect 110 272 113 338
rect 146 238 150 241
rect 6 182 9 198
rect 158 162 161 198
rect 166 162 169 358
rect 234 348 238 351
rect 254 242 257 438
rect 518 432 521 438
rect 262 342 265 358
rect 582 352 585 548
rect 710 432 713 568
rect 722 528 729 531
rect 610 428 614 431
rect 600 403 602 407
rect 606 403 609 407
rect 614 403 616 407
rect 726 382 729 528
rect 750 432 753 568
rect 782 538 790 541
rect 782 352 785 538
rect 906 468 910 471
rect 958 462 961 478
rect 842 458 846 461
rect 830 452 833 458
rect 962 448 966 451
rect 1074 448 1078 451
rect 298 348 302 351
rect 578 338 582 341
rect 646 338 654 341
rect 538 328 542 331
rect 506 318 510 321
rect 502 302 505 318
rect 274 268 278 271
rect 262 242 265 268
rect 502 242 505 268
rect 246 232 249 238
rect 182 152 185 188
rect 226 168 230 171
rect 314 168 318 171
rect 242 148 246 151
rect 362 148 366 151
rect 406 122 409 138
rect 438 132 441 138
rect 342 52 345 108
rect 438 52 441 68
rect 470 52 473 68
rect 462 12 465 18
rect 502 12 505 238
rect 550 222 553 258
rect 646 252 649 338
rect 750 252 753 348
rect 758 342 761 348
rect 978 338 982 341
rect 1042 338 1046 341
rect 866 328 870 331
rect 830 322 833 328
rect 858 268 862 271
rect 1006 268 1014 271
rect 600 203 602 207
rect 606 203 609 207
rect 614 203 616 207
rect 718 162 721 228
rect 714 158 718 161
rect 702 152 705 158
rect 702 112 705 118
rect 666 58 670 61
rect 614 22 617 28
rect 750 12 753 248
rect 1006 222 1009 268
rect 1054 212 1057 238
rect 762 128 766 131
rect 798 92 801 208
rect 798 72 801 78
rect 846 72 849 118
rect 854 82 857 188
rect 942 142 945 178
rect 890 128 897 131
rect 894 122 897 128
rect 958 92 961 98
rect 958 82 961 88
rect 810 68 814 71
rect 954 18 958 21
rect 50 8 54 11
rect 918 11 921 18
rect 914 8 921 11
rect 974 12 977 198
rect 1006 122 1009 168
rect 1042 58 1046 61
rect 1054 12 1057 208
rect 1070 112 1073 118
rect 1062 72 1065 78
rect 1070 72 1073 78
rect 1062 62 1065 68
rect 1062 22 1065 58
rect 1078 12 1081 358
rect 1094 312 1097 568
rect 1102 512 1105 528
rect 1112 503 1114 507
rect 1118 503 1121 507
rect 1126 503 1128 507
rect 1174 422 1177 568
rect 1366 558 1374 561
rect 1170 308 1177 311
rect 1112 303 1114 307
rect 1118 303 1121 307
rect 1126 303 1128 307
rect 1102 292 1105 298
rect 1174 292 1177 308
rect 1086 72 1089 268
rect 1198 262 1201 548
rect 1282 528 1286 531
rect 1254 441 1257 458
rect 1270 442 1273 508
rect 1366 452 1369 558
rect 1254 438 1265 441
rect 1262 422 1265 438
rect 1446 412 1449 448
rect 1478 412 1481 728
rect 1254 262 1257 328
rect 1262 322 1265 328
rect 1094 22 1097 248
rect 1158 132 1161 218
rect 1174 152 1177 218
rect 1198 152 1201 258
rect 1326 242 1329 328
rect 1422 322 1425 398
rect 1502 352 1505 448
rect 1518 382 1521 538
rect 1526 412 1529 738
rect 1582 692 1585 868
rect 1582 532 1585 568
rect 1550 462 1553 508
rect 1582 432 1585 528
rect 1474 328 1478 331
rect 1518 272 1521 378
rect 1590 342 1593 668
rect 1170 148 1174 151
rect 1202 128 1209 131
rect 1206 122 1209 128
rect 1234 118 1238 121
rect 1112 103 1114 107
rect 1118 103 1121 107
rect 1126 103 1128 107
rect 1134 92 1137 98
rect 1206 22 1209 118
rect 1214 52 1217 58
rect 1286 12 1289 148
rect 1358 142 1361 268
rect 1354 138 1358 141
rect 1322 128 1326 131
rect 1338 68 1345 71
rect 1342 62 1345 68
rect 1310 22 1313 28
rect 1350 12 1353 138
rect 1366 131 1369 158
rect 1510 152 1513 248
rect 1358 128 1369 131
rect 1358 112 1361 128
rect 1406 112 1409 148
rect 1506 118 1510 121
rect 1534 112 1537 158
rect 1606 82 1609 1138
rect 1634 1058 1638 1061
rect 1630 542 1633 928
rect 1638 662 1641 908
rect 1646 551 1649 1428
rect 1654 1322 1657 1468
rect 1662 1452 1665 1458
rect 1654 862 1657 1308
rect 1662 1262 1665 1378
rect 1670 1292 1673 1328
rect 1670 982 1673 1288
rect 1674 978 1681 981
rect 1646 548 1654 551
rect 1618 448 1622 451
rect 1622 402 1625 438
rect 1614 362 1617 368
rect 1622 352 1625 388
rect 1630 372 1633 538
rect 1634 358 1638 361
rect 1626 148 1630 151
rect 1662 72 1665 658
rect 1670 72 1673 368
rect 1678 122 1681 978
rect 1718 932 1721 1358
rect 1686 291 1689 538
rect 1686 288 1694 291
rect 1702 72 1705 888
rect 1734 552 1737 578
rect 1726 442 1729 468
rect 1734 452 1737 488
rect 1726 362 1729 418
rect 1402 58 1409 61
rect 1406 52 1409 58
rect 600 3 602 7
rect 606 3 609 7
rect 614 3 616 7
<< m5contact >>
rect 374 1538 378 1542
rect 46 1338 50 1342
rect 602 1603 606 1607
rect 609 1603 610 1607
rect 610 1603 613 1607
rect 470 1538 474 1542
rect 262 1338 266 1342
rect 62 1108 66 1112
rect 14 578 18 582
rect 78 578 82 582
rect 134 568 138 572
rect 198 1058 202 1062
rect 198 868 202 872
rect 158 548 162 552
rect 254 1108 258 1112
rect 222 858 226 862
rect 254 858 258 862
rect 246 848 250 852
rect 602 1403 606 1407
rect 609 1403 610 1407
rect 610 1403 613 1407
rect 542 1358 546 1362
rect 566 1358 570 1362
rect 390 1058 394 1062
rect 654 1338 658 1342
rect 494 1108 498 1112
rect 302 948 306 952
rect 366 948 370 952
rect 430 938 434 942
rect 302 868 306 872
rect 326 858 330 862
rect 342 858 346 862
rect 438 848 442 852
rect 334 728 338 732
rect 238 648 242 652
rect 582 1038 586 1042
rect 574 948 578 952
rect 602 1203 606 1207
rect 609 1203 610 1207
rect 610 1203 613 1207
rect 974 1518 978 1522
rect 602 1003 606 1007
rect 609 1003 610 1007
rect 610 1003 613 1007
rect 646 848 650 852
rect 602 803 606 807
rect 609 803 610 807
rect 610 803 613 807
rect 382 648 386 652
rect 454 588 458 592
rect 678 1068 682 1072
rect 670 868 674 872
rect 758 858 762 862
rect 694 768 698 772
rect 806 1068 810 1072
rect 790 848 794 852
rect 846 1038 850 1042
rect 966 1348 970 1352
rect 1046 1518 1050 1522
rect 990 948 994 952
rect 958 858 962 862
rect 934 768 938 772
rect 734 728 738 732
rect 1054 938 1058 942
rect 1006 868 1010 872
rect 602 603 606 607
rect 609 603 610 607
rect 610 603 613 607
rect 1114 1503 1118 1507
rect 1121 1503 1122 1507
rect 1122 1503 1125 1507
rect 1150 1348 1154 1352
rect 1214 1338 1218 1342
rect 1114 1303 1118 1307
rect 1121 1303 1122 1307
rect 1122 1303 1125 1307
rect 1102 1268 1106 1272
rect 1134 1268 1138 1272
rect 1310 1538 1314 1542
rect 1422 1538 1426 1542
rect 1326 1338 1330 1342
rect 1114 1103 1118 1107
rect 1121 1103 1122 1107
rect 1122 1103 1125 1107
rect 1158 1058 1162 1062
rect 1114 903 1118 907
rect 1121 903 1122 907
rect 1122 903 1125 907
rect 1114 703 1118 707
rect 1121 703 1122 707
rect 1122 703 1125 707
rect 622 588 626 592
rect 550 578 554 582
rect 422 568 426 572
rect 14 458 18 462
rect 222 458 226 462
rect 374 558 378 562
rect 382 548 386 552
rect 638 558 642 562
rect 286 468 290 472
rect 222 358 226 362
rect 142 238 146 242
rect 238 348 242 352
rect 518 428 522 432
rect 262 358 266 362
rect 606 428 610 432
rect 602 403 606 407
rect 609 403 610 407
rect 610 403 613 407
rect 902 468 906 472
rect 838 458 842 462
rect 830 448 834 452
rect 958 448 962 452
rect 1078 448 1082 452
rect 294 348 298 352
rect 574 338 578 342
rect 542 328 546 332
rect 502 318 506 322
rect 278 268 282 272
rect 246 238 250 242
rect 158 158 162 162
rect 222 168 226 172
rect 310 168 314 172
rect 246 148 250 152
rect 358 148 362 152
rect 438 128 442 132
rect 406 118 410 122
rect 470 68 474 72
rect 758 338 762 342
rect 982 338 986 342
rect 1038 338 1042 342
rect 862 328 866 332
rect 830 318 834 322
rect 854 268 858 272
rect 602 203 606 207
rect 609 203 610 207
rect 610 203 613 207
rect 710 158 714 162
rect 702 148 706 152
rect 702 108 706 112
rect 670 58 674 62
rect 614 18 618 22
rect 1054 238 1058 242
rect 758 128 762 132
rect 798 78 802 82
rect 942 138 946 142
rect 894 118 898 122
rect 958 88 962 92
rect 814 68 818 72
rect 918 18 922 22
rect 950 18 954 22
rect 46 8 50 12
rect 462 8 466 12
rect 1038 58 1042 62
rect 1070 108 1074 112
rect 1062 68 1066 72
rect 1070 68 1074 72
rect 1062 58 1066 62
rect 1102 528 1106 532
rect 1114 503 1118 507
rect 1121 503 1122 507
rect 1122 503 1125 507
rect 1114 303 1118 307
rect 1121 303 1122 307
rect 1122 303 1125 307
rect 1102 288 1106 292
rect 1174 288 1178 292
rect 1278 528 1282 532
rect 1262 318 1266 322
rect 1470 328 1474 332
rect 1326 238 1330 242
rect 1174 148 1178 152
rect 1206 118 1210 122
rect 1238 118 1242 122
rect 1114 103 1118 107
rect 1121 103 1122 107
rect 1122 103 1125 107
rect 1134 88 1138 92
rect 1214 48 1218 52
rect 1350 138 1354 142
rect 1326 128 1330 132
rect 1342 58 1346 62
rect 1310 18 1314 22
rect 1406 148 1410 152
rect 1502 118 1506 122
rect 1630 1058 1634 1062
rect 1662 1458 1666 1462
rect 1654 1308 1658 1312
rect 1622 448 1626 452
rect 1614 358 1618 362
rect 1630 368 1634 372
rect 1630 358 1634 362
rect 1630 148 1634 152
rect 1670 368 1674 372
rect 1734 448 1738 452
rect 1406 48 1410 52
rect 602 3 606 7
rect 609 3 610 7
rect 610 3 613 7
<< metal5 >>
rect 606 1603 609 1607
rect 606 1602 610 1603
rect 378 1538 470 1541
rect 1314 1538 1422 1541
rect 978 1518 1046 1521
rect 1118 1503 1121 1507
rect 1118 1502 1122 1503
rect 1662 1453 1665 1458
rect 606 1403 609 1407
rect 606 1402 610 1403
rect 546 1358 566 1361
rect 970 1348 1150 1351
rect 50 1338 262 1341
rect 266 1338 654 1341
rect 1218 1338 1326 1341
rect 1658 1308 1661 1311
rect 1118 1303 1121 1307
rect 1118 1302 1122 1303
rect 1106 1268 1134 1271
rect 606 1203 609 1207
rect 606 1202 610 1203
rect 66 1108 254 1111
rect 258 1108 494 1111
rect 1118 1103 1121 1107
rect 1118 1102 1122 1103
rect 682 1068 806 1071
rect 202 1058 390 1061
rect 1162 1058 1630 1061
rect 586 1038 846 1041
rect 606 1003 609 1007
rect 606 1002 610 1003
rect 306 948 366 951
rect 578 948 990 951
rect 434 938 1054 941
rect 1118 903 1121 907
rect 1118 902 1122 903
rect 202 868 302 871
rect 674 868 1006 871
rect 226 858 254 861
rect 330 858 342 861
rect 762 858 958 861
rect 250 848 438 851
rect 650 848 790 851
rect 606 803 609 807
rect 606 802 610 803
rect 698 768 934 771
rect 338 728 734 731
rect 1118 703 1121 707
rect 1118 702 1122 703
rect 242 648 382 651
rect 606 603 609 607
rect 606 602 610 603
rect 458 588 622 591
rect 18 578 78 581
rect 82 578 550 581
rect 138 568 422 571
rect 378 558 638 561
rect 162 548 382 551
rect 1106 528 1278 531
rect 1118 503 1121 507
rect 1118 502 1122 503
rect 290 468 902 471
rect 18 458 222 461
rect 226 458 838 461
rect 834 448 958 451
rect 1082 448 1622 451
rect 1626 448 1734 451
rect 522 428 606 431
rect 606 403 609 407
rect 606 402 610 403
rect 1634 368 1670 371
rect 226 358 262 361
rect 1618 358 1630 361
rect 242 348 294 351
rect 578 338 758 341
rect 986 338 1038 341
rect 546 328 862 331
rect 866 328 1470 331
rect 506 318 830 321
rect 834 318 1262 321
rect 1118 303 1121 307
rect 1118 302 1122 303
rect 1106 288 1174 291
rect 282 268 854 271
rect 146 238 246 241
rect 1058 238 1326 241
rect 606 203 609 207
rect 606 202 610 203
rect 226 168 310 171
rect 162 158 710 161
rect 250 148 358 151
rect 706 148 1174 151
rect 1410 148 1630 151
rect 946 138 1350 141
rect 442 128 758 131
rect 762 128 1326 131
rect 410 118 894 121
rect 898 118 1206 121
rect 1242 118 1502 121
rect 706 108 1070 111
rect 1118 103 1121 107
rect 1118 102 1122 103
rect 962 88 1134 91
rect 802 78 1073 81
rect 1070 72 1073 78
rect 474 68 814 71
rect 818 68 1062 71
rect 674 58 1038 61
rect 1066 58 1342 61
rect 1218 48 1406 51
rect 618 18 918 21
rect 954 18 1310 21
rect 50 8 462 11
rect 606 3 609 7
rect 606 2 610 3
<< m6contact >>
rect 600 1607 606 1608
rect 610 1607 616 1608
rect 600 1603 602 1607
rect 602 1603 606 1607
rect 610 1603 613 1607
rect 613 1603 616 1607
rect 600 1602 606 1603
rect 610 1602 616 1603
rect 1112 1507 1118 1508
rect 1122 1507 1128 1508
rect 1112 1503 1114 1507
rect 1114 1503 1118 1507
rect 1122 1503 1125 1507
rect 1125 1503 1128 1507
rect 1112 1502 1118 1503
rect 1122 1502 1128 1503
rect 1661 1447 1667 1453
rect 600 1407 606 1408
rect 610 1407 616 1408
rect 600 1403 602 1407
rect 602 1403 606 1407
rect 610 1403 613 1407
rect 613 1403 616 1407
rect 600 1402 606 1403
rect 610 1402 616 1403
rect 1112 1307 1118 1308
rect 1122 1307 1128 1308
rect 1661 1307 1667 1313
rect 1112 1303 1114 1307
rect 1114 1303 1118 1307
rect 1122 1303 1125 1307
rect 1125 1303 1128 1307
rect 1112 1302 1118 1303
rect 1122 1302 1128 1303
rect 600 1207 606 1208
rect 610 1207 616 1208
rect 600 1203 602 1207
rect 602 1203 606 1207
rect 610 1203 613 1207
rect 613 1203 616 1207
rect 600 1202 606 1203
rect 610 1202 616 1203
rect 1112 1107 1118 1108
rect 1122 1107 1128 1108
rect 1112 1103 1114 1107
rect 1114 1103 1118 1107
rect 1122 1103 1125 1107
rect 1125 1103 1128 1107
rect 1112 1102 1118 1103
rect 1122 1102 1128 1103
rect 600 1007 606 1008
rect 610 1007 616 1008
rect 600 1003 602 1007
rect 602 1003 606 1007
rect 610 1003 613 1007
rect 613 1003 616 1007
rect 600 1002 606 1003
rect 610 1002 616 1003
rect 1112 907 1118 908
rect 1122 907 1128 908
rect 1112 903 1114 907
rect 1114 903 1118 907
rect 1122 903 1125 907
rect 1125 903 1128 907
rect 1112 902 1118 903
rect 1122 902 1128 903
rect 600 807 606 808
rect 610 807 616 808
rect 600 803 602 807
rect 602 803 606 807
rect 610 803 613 807
rect 613 803 616 807
rect 600 802 606 803
rect 610 802 616 803
rect 1112 707 1118 708
rect 1122 707 1128 708
rect 1112 703 1114 707
rect 1114 703 1118 707
rect 1122 703 1125 707
rect 1125 703 1128 707
rect 1112 702 1118 703
rect 1122 702 1128 703
rect 600 607 606 608
rect 610 607 616 608
rect 600 603 602 607
rect 602 603 606 607
rect 610 603 613 607
rect 613 603 616 607
rect 600 602 606 603
rect 610 602 616 603
rect 1112 507 1118 508
rect 1122 507 1128 508
rect 1112 503 1114 507
rect 1114 503 1118 507
rect 1122 503 1125 507
rect 1125 503 1128 507
rect 1112 502 1118 503
rect 1122 502 1128 503
rect 600 407 606 408
rect 610 407 616 408
rect 600 403 602 407
rect 602 403 606 407
rect 610 403 613 407
rect 613 403 616 407
rect 600 402 606 403
rect 610 402 616 403
rect 1112 307 1118 308
rect 1122 307 1128 308
rect 1112 303 1114 307
rect 1114 303 1118 307
rect 1122 303 1125 307
rect 1125 303 1128 307
rect 1112 302 1118 303
rect 1122 302 1128 303
rect 600 207 606 208
rect 610 207 616 208
rect 600 203 602 207
rect 602 203 606 207
rect 610 203 613 207
rect 613 203 616 207
rect 600 202 606 203
rect 610 202 616 203
rect 1112 107 1118 108
rect 1122 107 1128 108
rect 1112 103 1114 107
rect 1114 103 1118 107
rect 1122 103 1125 107
rect 1125 103 1128 107
rect 1112 102 1118 103
rect 1122 102 1128 103
rect 600 7 606 8
rect 610 7 616 8
rect 600 3 602 7
rect 602 3 606 7
rect 610 3 613 7
rect 613 3 616 7
rect 600 2 606 3
rect 610 2 616 3
<< metal6 >>
rect 600 1608 616 1640
rect 606 1602 610 1608
rect 600 1408 616 1602
rect 606 1402 610 1408
rect 600 1208 616 1402
rect 606 1202 610 1208
rect 600 1008 616 1202
rect 606 1002 610 1008
rect 600 808 616 1002
rect 606 802 610 808
rect 600 608 616 802
rect 606 602 610 608
rect 600 408 616 602
rect 606 402 610 408
rect 600 208 616 402
rect 606 202 610 208
rect 600 8 616 202
rect 606 2 610 8
rect 600 -30 616 2
rect 1112 1508 1128 1640
rect 1118 1502 1122 1508
rect 1112 1308 1128 1502
rect 1118 1302 1122 1308
rect 1661 1313 1666 1447
rect 1112 1108 1128 1302
rect 1118 1102 1122 1108
rect 1112 908 1128 1102
rect 1118 902 1122 908
rect 1112 708 1128 902
rect 1118 702 1122 708
rect 1112 508 1128 702
rect 1118 502 1122 508
rect 1112 308 1128 502
rect 1118 302 1122 308
rect 1112 108 1128 302
rect 1118 102 1122 108
rect 1112 -30 1128 102
use INVX1  _966_
timestamp 1563080643
transform 1 0 4 0 1 1505
box -2 -3 18 103
use NAND2X1  _967_
timestamp 1563080643
transform -1 0 44 0 1 1505
box -2 -3 26 103
use NAND2X1  _970_
timestamp 1563080643
transform 1 0 44 0 1 1505
box -2 -3 26 103
use INVX1  _1301_
timestamp 1563080643
transform -1 0 84 0 1 1505
box -2 -3 18 103
use OAI21X1  _1303_
timestamp 1563080643
transform 1 0 84 0 1 1505
box -2 -3 34 103
use NAND2X1  _1302_
timestamp 1563080643
transform -1 0 140 0 1 1505
box -2 -3 26 103
use NAND2X1  _1050_
timestamp 1563080643
transform 1 0 140 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_insert37
timestamp 1563080643
transform -1 0 188 0 1 1505
box -2 -3 26 103
use NAND2X1  _1382_
timestamp 1563080643
transform 1 0 188 0 1 1505
box -2 -3 26 103
use NAND2X1  _1047_
timestamp 1563080643
transform 1 0 212 0 1 1505
box -2 -3 26 103
use INVX1  _1046_
timestamp 1563080643
transform -1 0 252 0 1 1505
box -2 -3 18 103
use NAND2X1  _1089_
timestamp 1563080643
transform 1 0 252 0 1 1505
box -2 -3 26 103
use INVX1  _803_
timestamp 1563080643
transform 1 0 276 0 1 1505
box -2 -3 18 103
use INVX1  _1088_
timestamp 1563080643
transform -1 0 308 0 1 1505
box -2 -3 18 103
use INVX1  _1135_
timestamp 1563080643
transform 1 0 308 0 1 1505
box -2 -3 18 103
use OAI21X1  _805_
timestamp 1563080643
transform 1 0 324 0 1 1505
box -2 -3 34 103
use NAND2X1  _804_
timestamp 1563080643
transform -1 0 380 0 1 1505
box -2 -3 26 103
use NAND2X1  _1136_
timestamp 1563080643
transform -1 0 404 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_insert33
timestamp 1563080643
transform -1 0 428 0 1 1505
box -2 -3 26 103
use NAND2X1  _923_
timestamp 1563080643
transform 1 0 428 0 1 1505
box -2 -3 26 103
use NAND2X1  _801_
timestamp 1563080643
transform 1 0 452 0 1 1505
box -2 -3 26 103
use INVX1  _800_
timestamp 1563080643
transform -1 0 492 0 1 1505
box -2 -3 18 103
use NAND2X1  _806_
timestamp 1563080643
transform -1 0 516 0 1 1505
box -2 -3 26 103
use NAND2X1  _1216_
timestamp 1563080643
transform 1 0 516 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_insert32
timestamp 1563080643
transform 1 0 540 0 1 1505
box -2 -3 26 103
use INVX1  _883_
timestamp 1563080643
transform 1 0 564 0 1 1505
box -2 -3 18 103
use OAI21X1  _885_
timestamp 1563080643
transform 1 0 580 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_0_0
timestamp 1563080643
transform -1 0 620 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1563080643
transform -1 0 628 0 1 1505
box -2 -3 10 103
use NAND2X1  _884_
timestamp 1563080643
transform -1 0 652 0 1 1505
box -2 -3 26 103
use NAND2X1  _881_
timestamp 1563080643
transform 1 0 652 0 1 1505
box -2 -3 26 103
use INVX1  _880_
timestamp 1563080643
transform -1 0 692 0 1 1505
box -2 -3 18 103
use NAND2X1  _886_
timestamp 1563080643
transform -1 0 716 0 1 1505
box -2 -3 26 103
use NAND2X1  _920_
timestamp 1563080643
transform 1 0 716 0 1 1505
box -2 -3 26 103
use INVX1  _919_
timestamp 1563080643
transform -1 0 756 0 1 1505
box -2 -3 18 103
use NOR2X1  _1515_
timestamp 1563080643
transform -1 0 780 0 1 1505
box -2 -3 26 103
use NAND2X1  _1514_
timestamp 1563080643
transform -1 0 804 0 1 1505
box -2 -3 26 103
use DFFPOSX1  _1612_
timestamp 1563080643
transform -1 0 900 0 1 1505
box -2 -3 98 103
use INVX2  _1509_
timestamp 1563080643
transform -1 0 916 0 1 1505
box -2 -3 18 103
use OAI22X1  _1511_
timestamp 1563080643
transform 1 0 916 0 1 1505
box -2 -3 42 103
use OAI22X1  _1504_
timestamp 1563080643
transform 1 0 956 0 1 1505
box -2 -3 42 103
use NOR2X1  _1505_
timestamp 1563080643
transform -1 0 1020 0 1 1505
box -2 -3 26 103
use NAND2X1  _1513_
timestamp 1563080643
transform 1 0 1020 0 1 1505
box -2 -3 26 103
use AOI21X1  _1512_
timestamp 1563080643
transform -1 0 1076 0 1 1505
box -2 -3 34 103
use NAND2X1  _1506_
timestamp 1563080643
transform -1 0 1100 0 1 1505
box -2 -3 26 103
use NOR2X1  _1495_
timestamp 1563080643
transform -1 0 1124 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_1_0
timestamp 1563080643
transform 1 0 1124 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1563080643
transform 1 0 1132 0 1 1505
box -2 -3 10 103
use INVX1  _1577_
timestamp 1563080643
transform 1 0 1140 0 1 1505
box -2 -3 18 103
use NAND2X1  _1588_
timestamp 1563080643
transform 1 0 1156 0 1 1505
box -2 -3 26 103
use AOI22X1  _1578_
timestamp 1563080643
transform 1 0 1180 0 1 1505
box -2 -3 42 103
use NOR3X1  _1576_
timestamp 1563080643
transform 1 0 1220 0 1 1505
box -2 -3 66 103
use INVX1  _1499_
timestamp 1563080643
transform 1 0 1284 0 1 1505
box -2 -3 18 103
use OAI21X1  _1589_
timestamp 1563080643
transform -1 0 1332 0 1 1505
box -2 -3 34 103
use AOI21X1  _1548_
timestamp 1563080643
transform -1 0 1364 0 1 1505
box -2 -3 34 103
use OAI21X1  _1547_
timestamp 1563080643
transform -1 0 1396 0 1 1505
box -2 -3 34 103
use NOR2X1  _1598_
timestamp 1563080643
transform -1 0 1420 0 1 1505
box -2 -3 26 103
use AOI21X1  _1590_
timestamp 1563080643
transform -1 0 1452 0 1 1505
box -2 -3 34 103
use NAND2X1  _1572_
timestamp 1563080643
transform -1 0 1476 0 1 1505
box -2 -3 26 103
use NAND3X1  _1599_
timestamp 1563080643
transform 1 0 1476 0 1 1505
box -2 -3 34 103
use NAND3X1  _1587_
timestamp 1563080643
transform -1 0 1540 0 1 1505
box -2 -3 34 103
use NAND2X1  _1591_
timestamp 1563080643
transform 1 0 1540 0 1 1505
box -2 -3 26 103
use OAI21X1  _1600_
timestamp 1563080643
transform 1 0 1564 0 1 1505
box -2 -3 34 103
use NAND2X1  _1592_
timestamp 1563080643
transform 1 0 1596 0 1 1505
box -2 -3 26 103
use DFFPOSX1  _1603_
timestamp 1563080643
transform 1 0 1620 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_1
timestamp 1563080643
transform 1 0 1716 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1563080643
transform 1 0 1724 0 1 1505
box -2 -3 10 103
use NAND3X1  _968_
timestamp 1563080643
transform -1 0 36 0 -1 1505
box -2 -3 34 103
use OR2X2  _965_
timestamp 1563080643
transform -1 0 68 0 -1 1505
box -2 -3 34 103
use OAI21X1  _971_
timestamp 1563080643
transform -1 0 100 0 -1 1505
box -2 -3 34 103
use INVX1  _969_
timestamp 1563080643
transform -1 0 116 0 -1 1505
box -2 -3 18 103
use BUFX2  BUFX2_insert28
timestamp 1563080643
transform 1 0 116 0 -1 1505
box -2 -3 26 103
use OAI21X1  _1051_
timestamp 1563080643
transform -1 0 172 0 -1 1505
box -2 -3 34 103
use INVX1  _1298_
timestamp 1563080643
transform -1 0 188 0 -1 1505
box -2 -3 18 103
use INVX1  _1049_
timestamp 1563080643
transform -1 0 204 0 -1 1505
box -2 -3 18 103
use NAND3X1  _1048_
timestamp 1563080643
transform 1 0 204 0 -1 1505
box -2 -3 34 103
use OR2X2  _1045_
timestamp 1563080643
transform -1 0 268 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1090_
timestamp 1563080643
transform -1 0 300 0 -1 1505
box -2 -3 34 103
use INVX1  _1378_
timestamp 1563080643
transform -1 0 316 0 -1 1505
box -2 -3 18 103
use OAI21X1  _1383_
timestamp 1563080643
transform -1 0 348 0 -1 1505
box -2 -3 34 103
use INVX1  _1381_
timestamp 1563080643
transform -1 0 364 0 -1 1505
box -2 -3 18 103
use OAI21X1  _1137_
timestamp 1563080643
transform 1 0 364 0 -1 1505
box -2 -3 34 103
use BUFX2  BUFX2_insert16
timestamp 1563080643
transform -1 0 420 0 -1 1505
box -2 -3 26 103
use INVX1  _922_
timestamp 1563080643
transform 1 0 420 0 -1 1505
box -2 -3 18 103
use OAI21X1  _924_
timestamp 1563080643
transform 1 0 436 0 -1 1505
box -2 -3 34 103
use OR2X2  _799_
timestamp 1563080643
transform 1 0 468 0 -1 1505
box -2 -3 34 103
use INVX1  _1132_
timestamp 1563080643
transform 1 0 500 0 -1 1505
box -2 -3 18 103
use NAND3X1  _802_
timestamp 1563080643
transform -1 0 548 0 -1 1505
box -2 -3 34 103
use INVX1  _1215_
timestamp 1563080643
transform 1 0 548 0 -1 1505
box -2 -3 18 103
use NAND3X1  _807_
timestamp 1563080643
transform -1 0 596 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_0_0
timestamp 1563080643
transform 1 0 596 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1563080643
transform 1 0 604 0 -1 1505
box -2 -3 10 103
use OR2X2  _879_
timestamp 1563080643
transform 1 0 612 0 -1 1505
box -2 -3 34 103
use NAND3X1  _882_
timestamp 1563080643
transform 1 0 644 0 -1 1505
box -2 -3 34 103
use NAND3X1  _887_
timestamp 1563080643
transform 1 0 676 0 -1 1505
box -2 -3 34 103
use INVX1  _1212_
timestamp 1563080643
transform 1 0 708 0 -1 1505
box -2 -3 18 103
use AOI21X1  _1517_
timestamp 1563080643
transform 1 0 724 0 -1 1505
box -2 -3 34 103
use NOR2X1  _1516_
timestamp 1563080643
transform 1 0 756 0 -1 1505
box -2 -3 26 103
use NAND2X1  _1519_
timestamp 1563080643
transform 1 0 780 0 -1 1505
box -2 -3 26 103
use NAND3X1  _1522_
timestamp 1563080643
transform 1 0 804 0 -1 1505
box -2 -3 34 103
use INVX1  _1502_
timestamp 1563080643
transform 1 0 836 0 -1 1505
box -2 -3 18 103
use INVX2  _1500_
timestamp 1563080643
transform 1 0 852 0 -1 1505
box -2 -3 18 103
use AOI22X1  _1526_
timestamp 1563080643
transform 1 0 868 0 -1 1505
box -2 -3 42 103
use INVX2  _1510_
timestamp 1563080643
transform -1 0 924 0 -1 1505
box -2 -3 18 103
use NAND3X1  _1543_
timestamp 1563080643
transform -1 0 956 0 -1 1505
box -2 -3 34 103
use NAND2X1  _1542_
timestamp 1563080643
transform 1 0 956 0 -1 1505
box -2 -3 26 103
use NOR2X1  _1501_
timestamp 1563080643
transform -1 0 1004 0 -1 1505
box -2 -3 26 103
use NAND3X1  _1544_
timestamp 1563080643
transform -1 0 1036 0 -1 1505
box -2 -3 34 103
use INVX4  _1466_
timestamp 1563080643
transform 1 0 1036 0 -1 1505
box -2 -3 26 103
use OAI21X1  _1497_
timestamp 1563080643
transform -1 0 1092 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1498_
timestamp 1563080643
transform -1 0 1124 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_1_0
timestamp 1563080643
transform -1 0 1132 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1563080643
transform -1 0 1140 0 -1 1505
box -2 -3 10 103
use NAND3X1  _1575_
timestamp 1563080643
transform -1 0 1172 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1583_
timestamp 1563080643
transform 1 0 1172 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1574_
timestamp 1563080643
transform -1 0 1236 0 -1 1505
box -2 -3 34 103
use NAND3X1  _1573_
timestamp 1563080643
transform 1 0 1236 0 -1 1505
box -2 -3 34 103
use AOI21X1  _1582_
timestamp 1563080643
transform -1 0 1300 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1580_
timestamp 1563080643
transform -1 0 1332 0 -1 1505
box -2 -3 34 103
use NOR3X1  _1579_
timestamp 1563080643
transform -1 0 1396 0 -1 1505
box -2 -3 66 103
use OAI21X1  _1554_
timestamp 1563080643
transform 1 0 1396 0 -1 1505
box -2 -3 34 103
use AOI22X1  _1571_
timestamp 1563080643
transform -1 0 1468 0 -1 1505
box -2 -3 42 103
use AOI22X1  _1585_
timestamp 1563080643
transform -1 0 1508 0 -1 1505
box -2 -3 42 103
use NOR2X1  _1595_
timestamp 1563080643
transform 1 0 1508 0 -1 1505
box -2 -3 26 103
use NAND3X1  _1596_
timestamp 1563080643
transform 1 0 1532 0 -1 1505
box -2 -3 34 103
use OAI21X1  _1597_
timestamp 1563080643
transform 1 0 1564 0 -1 1505
box -2 -3 34 103
use NOR2X1  _1586_
timestamp 1563080643
transform 1 0 1596 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  _784_
timestamp 1563080643
transform 1 0 1620 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1563080643
transform -1 0 1724 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1563080643
transform -1 0 1732 0 -1 1505
box -2 -3 10 103
use BUFX2  BUFX2_insert29
timestamp 1563080643
transform 1 0 4 0 1 1305
box -2 -3 26 103
use NAND2X1  _972_
timestamp 1563080643
transform 1 0 28 0 1 1305
box -2 -3 26 103
use OR2X2  _1084_
timestamp 1563080643
transform 1 0 52 0 1 1305
box -2 -3 34 103
use NAND3X1  _1087_
timestamp 1563080643
transform 1 0 84 0 1 1305
box -2 -3 34 103
use NAND2X1  _1086_
timestamp 1563080643
transform 1 0 116 0 1 1305
box -2 -3 26 103
use NAND2X1  _1052_
timestamp 1563080643
transform -1 0 164 0 1 1305
box -2 -3 26 103
use NAND2X1  _1299_
timestamp 1563080643
transform -1 0 188 0 1 1305
box -2 -3 26 103
use NAND2X1  _1304_
timestamp 1563080643
transform -1 0 212 0 1 1305
box -2 -3 26 103
use NAND2X1  _1091_
timestamp 1563080643
transform 1 0 212 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_insert36
timestamp 1563080643
transform 1 0 236 0 1 1305
box -2 -3 26 103
use INVX1  _1085_
timestamp 1563080643
transform -1 0 276 0 1 1305
box -2 -3 18 103
use NAND2X1  _1379_
timestamp 1563080643
transform -1 0 300 0 1 1305
box -2 -3 26 103
use NAND2X1  _1384_
timestamp 1563080643
transform 1 0 300 0 1 1305
box -2 -3 26 103
use OR2X2  _1416_
timestamp 1563080643
transform 1 0 324 0 1 1305
box -2 -3 34 103
use NAND2X1  _1423_
timestamp 1563080643
transform 1 0 356 0 1 1305
box -2 -3 26 103
use INVX1  _1420_
timestamp 1563080643
transform 1 0 380 0 1 1305
box -2 -3 18 103
use OAI21X1  _1422_
timestamp 1563080643
transform 1 0 396 0 1 1305
box -2 -3 34 103
use NAND2X1  _1421_
timestamp 1563080643
transform 1 0 428 0 1 1305
box -2 -3 26 103
use INVX1  _1254_
timestamp 1563080643
transform 1 0 452 0 1 1305
box -2 -3 18 103
use OAI21X1  _1256_
timestamp 1563080643
transform 1 0 468 0 1 1305
box -2 -3 34 103
use NAND2X1  _1255_
timestamp 1563080643
transform -1 0 524 0 1 1305
box -2 -3 26 103
use NAND2X1  _1133_
timestamp 1563080643
transform -1 0 548 0 1 1305
box -2 -3 26 103
use OAI21X1  _1217_
timestamp 1563080643
transform -1 0 580 0 1 1305
box -2 -3 34 103
use NAND2X1  _1138_
timestamp 1563080643
transform -1 0 604 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_0_0
timestamp 1563080643
transform -1 0 612 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1563080643
transform -1 0 620 0 1 1305
box -2 -3 10 103
use NAND2X1  _1257_
timestamp 1563080643
transform -1 0 644 0 1 1305
box -2 -3 26 103
use OR2X2  _1250_
timestamp 1563080643
transform 1 0 644 0 1 1305
box -2 -3 34 103
use NAND2X1  _1218_
timestamp 1563080643
transform -1 0 700 0 1 1305
box -2 -3 26 103
use NAND2X1  _1213_
timestamp 1563080643
transform 1 0 700 0 1 1305
box -2 -3 26 103
use OR2X2  _918_
timestamp 1563080643
transform 1 0 724 0 1 1305
box -2 -3 34 103
use NAND3X1  _921_
timestamp 1563080643
transform -1 0 788 0 1 1305
box -2 -3 34 103
use NAND2X1  _925_
timestamp 1563080643
transform -1 0 812 0 1 1305
box -2 -3 26 103
use OAI21X1  _1528_
timestamp 1563080643
transform -1 0 844 0 1 1305
box -2 -3 34 103
use NOR2X1  _1523_
timestamp 1563080643
transform 1 0 844 0 1 1305
box -2 -3 26 103
use OAI21X1  _1527_
timestamp 1563080643
transform 1 0 868 0 1 1305
box -2 -3 34 103
use INVX2  _1503_
timestamp 1563080643
transform 1 0 900 0 1 1305
box -2 -3 18 103
use NAND3X1  _1555_
timestamp 1563080643
transform 1 0 916 0 1 1305
box -2 -3 34 103
use NAND3X1  _1518_
timestamp 1563080643
transform 1 0 948 0 1 1305
box -2 -3 34 103
use NAND3X1  _1550_
timestamp 1563080643
transform -1 0 1012 0 1 1305
box -2 -3 34 103
use NAND3X1  _1551_
timestamp 1563080643
transform -1 0 1044 0 1 1305
box -2 -3 34 103
use INVX1  _1507_
timestamp 1563080643
transform 1 0 1044 0 1 1305
box -2 -3 18 103
use NOR2X1  _1508_
timestamp 1563080643
transform -1 0 1084 0 1 1305
box -2 -3 26 103
use AOI21X1  _1530_
timestamp 1563080643
transform 1 0 1084 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1563080643
transform -1 0 1124 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1563080643
transform -1 0 1132 0 1 1305
box -2 -3 10 103
use AOI21X1  _1557_
timestamp 1563080643
transform -1 0 1164 0 1 1305
box -2 -3 34 103
use NOR2X1  _1562_
timestamp 1563080643
transform 1 0 1164 0 1 1305
box -2 -3 26 103
use INVX1  _1561_
timestamp 1563080643
transform -1 0 1204 0 1 1305
box -2 -3 18 103
use INVX1  _1531_
timestamp 1563080643
transform -1 0 1220 0 1 1305
box -2 -3 18 103
use NAND2X1  _1539_
timestamp 1563080643
transform 1 0 1220 0 1 1305
box -2 -3 26 103
use NAND3X1  _1541_
timestamp 1563080643
transform 1 0 1244 0 1 1305
box -2 -3 34 103
use OAI21X1  _1546_
timestamp 1563080643
transform 1 0 1276 0 1 1305
box -2 -3 34 103
use NOR2X1  _1545_
timestamp 1563080643
transform 1 0 1308 0 1 1305
box -2 -3 26 103
use OAI22X1  _1566_
timestamp 1563080643
transform 1 0 1332 0 1 1305
box -2 -3 42 103
use OAI21X1  _1581_
timestamp 1563080643
transform -1 0 1404 0 1 1305
box -2 -3 34 103
use OAI21X1  _1565_
timestamp 1563080643
transform -1 0 1436 0 1 1305
box -2 -3 34 103
use NOR2X1  _1564_
timestamp 1563080643
transform -1 0 1460 0 1 1305
box -2 -3 26 103
use NAND3X1  _1560_
timestamp 1563080643
transform -1 0 1492 0 1 1305
box -2 -3 34 103
use NAND2X1  _1558_
timestamp 1563080643
transform -1 0 1516 0 1 1305
box -2 -3 26 103
use OAI21X1  _1553_
timestamp 1563080643
transform -1 0 1548 0 1 1305
box -2 -3 34 103
use AND2X2  _1552_
timestamp 1563080643
transform -1 0 1580 0 1 1305
box -2 -3 34 103
use NAND3X1  _1570_
timestamp 1563080643
transform 1 0 1580 0 1 1305
box -2 -3 34 103
use INVX1  _1491_
timestamp 1563080643
transform 1 0 1612 0 1 1305
box -2 -3 18 103
use AOI21X1  _1569_
timestamp 1563080643
transform -1 0 1660 0 1 1305
box -2 -3 34 103
use OAI21X1  _1584_
timestamp 1563080643
transform 1 0 1660 0 1 1305
box -2 -3 34 103
use OAI21X1  _1594_
timestamp 1563080643
transform 1 0 1692 0 1 1305
box -2 -3 34 103
use FILL  FILL_14_1
timestamp 1563080643
transform 1 0 1724 0 1 1305
box -2 -3 10 103
use INVX4  _955_
timestamp 1563080643
transform -1 0 28 0 -1 1305
box -2 -3 26 103
use NAND3X1  _973_
timestamp 1563080643
transform -1 0 60 0 -1 1305
box -2 -3 34 103
use INVX4  _1287_
timestamp 1563080643
transform -1 0 84 0 -1 1305
box -2 -3 26 103
use NAND3X1  _1092_
timestamp 1563080643
transform 1 0 84 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1053_
timestamp 1563080643
transform 1 0 116 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1300_
timestamp 1563080643
transform -1 0 180 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1305_
timestamp 1563080643
transform -1 0 212 0 -1 1305
box -2 -3 34 103
use OR2X2  _1297_
timestamp 1563080643
transform -1 0 244 0 -1 1305
box -2 -3 34 103
use OR2X2  _1377_
timestamp 1563080643
transform 1 0 244 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1380_
timestamp 1563080643
transform -1 0 308 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1385_
timestamp 1563080643
transform -1 0 340 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1419_
timestamp 1563080643
transform 1 0 340 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1418_
timestamp 1563080643
transform -1 0 396 0 -1 1305
box -2 -3 26 103
use INVX1  _1417_
timestamp 1563080643
transform -1 0 412 0 -1 1305
box -2 -3 18 103
use NAND2X1  _1204_
timestamp 1563080643
transform -1 0 436 0 -1 1305
box -2 -3 26 103
use OR2X2  _1202_
timestamp 1563080643
transform 1 0 436 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1205_
timestamp 1563080643
transform -1 0 500 0 -1 1305
box -2 -3 34 103
use OR2X2  _1131_
timestamp 1563080643
transform 1 0 500 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1134_
timestamp 1563080643
transform -1 0 564 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_insert15
timestamp 1563080643
transform -1 0 588 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_0_0
timestamp 1563080643
transform -1 0 596 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1563080643
transform -1 0 604 0 -1 1305
box -2 -3 10 103
use NAND3X1  _1139_
timestamp 1563080643
transform -1 0 636 0 -1 1305
box -2 -3 34 103
use OR2X2  _1211_
timestamp 1563080643
transform 1 0 636 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1253_
timestamp 1563080643
transform 1 0 668 0 -1 1305
box -2 -3 34 103
use NAND3X1  _1214_
timestamp 1563080643
transform 1 0 700 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1252_
timestamp 1563080643
transform 1 0 732 0 -1 1305
box -2 -3 26 103
use INVX1  _1251_
timestamp 1563080643
transform -1 0 772 0 -1 1305
box -2 -3 18 103
use NAND3X1  _926_
timestamp 1563080643
transform 1 0 772 0 -1 1305
box -2 -3 34 103
use INVX4  _789_
timestamp 1563080643
transform 1 0 804 0 -1 1305
box -2 -3 26 103
use NAND2X1  _1521_
timestamp 1563080643
transform -1 0 852 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  _1611_
timestamp 1563080643
transform -1 0 948 0 -1 1305
box -2 -3 98 103
use INVX1  _1520_
timestamp 1563080643
transform 1 0 948 0 -1 1305
box -2 -3 18 103
use NAND2X1  _1549_
timestamp 1563080643
transform 1 0 964 0 -1 1305
box -2 -3 26 103
use NAND2X1  _1525_
timestamp 1563080643
transform -1 0 1012 0 -1 1305
box -2 -3 26 103
use NAND2X1  _1529_
timestamp 1563080643
transform 1 0 1012 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  _1607_
timestamp 1563080643
transform -1 0 1132 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_1_0
timestamp 1563080643
transform 1 0 1132 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1563080643
transform 1 0 1140 0 -1 1305
box -2 -3 10 103
use NAND2X1  _1556_
timestamp 1563080643
transform 1 0 1148 0 -1 1305
box -2 -3 26 103
use INVX1  _1524_
timestamp 1563080643
transform 1 0 1172 0 -1 1305
box -2 -3 18 103
use AND2X2  _1464_
timestamp 1563080643
transform -1 0 1220 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_insert43
timestamp 1563080643
transform -1 0 1244 0 -1 1305
box -2 -3 26 103
use OAI21X1  _1563_
timestamp 1563080643
transform -1 0 1276 0 -1 1305
box -2 -3 34 103
use AOI21X1  _1567_
timestamp 1563080643
transform 1 0 1276 0 -1 1305
box -2 -3 34 103
use AOI21X1  _1540_
timestamp 1563080643
transform -1 0 1340 0 -1 1305
box -2 -3 34 103
use NOR2X1  _1485_
timestamp 1563080643
transform -1 0 1364 0 -1 1305
box -2 -3 26 103
use INVX1  _1484_
timestamp 1563080643
transform -1 0 1380 0 -1 1305
box -2 -3 18 103
use NAND2X1  _1537_
timestamp 1563080643
transform 1 0 1380 0 -1 1305
box -2 -3 26 103
use AOI22X1  _1494_
timestamp 1563080643
transform 1 0 1404 0 -1 1305
box -2 -3 42 103
use NAND2X1  _1480_
timestamp 1563080643
transform -1 0 1468 0 -1 1305
box -2 -3 26 103
use AOI21X1  _1559_
timestamp 1563080643
transform -1 0 1500 0 -1 1305
box -2 -3 34 103
use NAND2X1  _1489_
timestamp 1563080643
transform 1 0 1500 0 -1 1305
box -2 -3 26 103
use AOI22X1  _1493_
timestamp 1563080643
transform 1 0 1524 0 -1 1305
box -2 -3 42 103
use NAND2X1  _1490_
timestamp 1563080643
transform -1 0 1588 0 -1 1305
box -2 -3 26 103
use NAND2X1  _1568_
timestamp 1563080643
transform -1 0 1612 0 -1 1305
box -2 -3 26 103
use NAND2X1  _1492_
timestamp 1563080643
transform -1 0 1636 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  _1602_
timestamp 1563080643
transform 1 0 1636 0 -1 1305
box -2 -3 98 103
use OR2X2  _1036_
timestamp 1563080643
transform 1 0 4 0 1 1105
box -2 -3 34 103
use NAND2X1  _1038_
timestamp 1563080643
transform 1 0 36 0 1 1105
box -2 -3 26 103
use INVX1  _1037_
timestamp 1563080643
transform -1 0 76 0 1 1105
box -2 -3 18 103
use INVX1  _1369_
timestamp 1563080643
transform 1 0 76 0 1 1105
box -2 -3 18 103
use NAND2X1  _1370_
timestamp 1563080643
transform -1 0 116 0 1 1105
box -2 -3 26 103
use NAND3X1  _1371_
timestamp 1563080643
transform -1 0 148 0 1 1105
box -2 -3 34 103
use OR2X2  _1368_
timestamp 1563080643
transform -1 0 180 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert38
timestamp 1563080643
transform 1 0 180 0 1 1105
box -2 -3 26 103
use INVX1  _1408_
timestamp 1563080643
transform 1 0 204 0 1 1105
box -2 -3 18 103
use NAND2X1  _1409_
timestamp 1563080643
transform -1 0 244 0 1 1105
box -2 -3 26 103
use OR2X2  _1294_
timestamp 1563080643
transform 1 0 244 0 1 1105
box -2 -3 34 103
use NAND3X1  _1295_
timestamp 1563080643
transform 1 0 276 0 1 1105
box -2 -3 34 103
use INVX1  _1203_
timestamp 1563080643
transform 1 0 308 0 1 1105
box -2 -3 18 103
use INVX1  _871_
timestamp 1563080643
transform 1 0 324 0 1 1105
box -2 -3 18 103
use NAND3X1  _1424_
timestamp 1563080643
transform 1 0 340 0 1 1105
box -2 -3 34 103
use NAND2X1  _872_
timestamp 1563080643
transform -1 0 396 0 1 1105
box -2 -3 26 103
use BUFX2  BUFX2_insert31
timestamp 1563080643
transform 1 0 396 0 1 1105
box -2 -3 26 103
use OR2X2  _870_
timestamp 1563080643
transform 1 0 420 0 1 1105
box -2 -3 34 103
use NAND3X1  _873_
timestamp 1563080643
transform -1 0 484 0 1 1105
box -2 -3 34 103
use OR2X2  _796_
timestamp 1563080643
transform 1 0 484 0 1 1105
box -2 -3 34 103
use NAND2X1  _795_
timestamp 1563080643
transform 1 0 516 0 1 1105
box -2 -3 26 103
use INVX1  _794_
timestamp 1563080643
transform -1 0 556 0 1 1105
box -2 -3 18 103
use NAND3X1  _797_
timestamp 1563080643
transform 1 0 556 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert30
timestamp 1563080643
transform -1 0 612 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_0_0
timestamp 1563080643
transform 1 0 612 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1563080643
transform 1 0 620 0 1 1105
box -2 -3 10 103
use BUFX2  BUFX2_insert34
timestamp 1563080643
transform 1 0 628 0 1 1105
box -2 -3 26 103
use NAND3X1  _1258_
timestamp 1563080643
transform -1 0 684 0 1 1105
box -2 -3 34 103
use NAND3X1  _1219_
timestamp 1563080643
transform -1 0 716 0 1 1105
box -2 -3 34 103
use DFFPOSX1  _1609_
timestamp 1563080643
transform -1 0 812 0 1 1105
box -2 -3 98 103
use DFFPOSX1  _1610_
timestamp 1563080643
transform 1 0 812 0 1 1105
box -2 -3 98 103
use DFFPOSX1  _1606_
timestamp 1563080643
transform -1 0 1004 0 1 1105
box -2 -3 98 103
use DFFPOSX1  _1604_
timestamp 1563080643
transform -1 0 1100 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_1_0
timestamp 1563080643
transform 1 0 1100 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1563080643
transform 1 0 1108 0 1 1105
box -2 -3 10 103
use DFFPOSX1  _1617_
timestamp 1563080643
transform 1 0 1116 0 1 1105
box -2 -3 98 103
use OAI21X1  _1496_
timestamp 1563080643
transform -1 0 1244 0 1 1105
box -2 -3 34 103
use NOR2X1  _1472_
timestamp 1563080643
transform -1 0 1268 0 1 1105
box -2 -3 26 103
use AND2X2  _1483_
timestamp 1563080643
transform 1 0 1268 0 1 1105
box -2 -3 34 103
use NOR2X1  _1482_
timestamp 1563080643
transform -1 0 1324 0 1 1105
box -2 -3 26 103
use OAI21X1  _1486_
timestamp 1563080643
transform 1 0 1324 0 1 1105
box -2 -3 34 103
use NAND2X1  _1470_
timestamp 1563080643
transform -1 0 1380 0 1 1105
box -2 -3 26 103
use OAI21X1  _1536_
timestamp 1563080643
transform 1 0 1380 0 1 1105
box -2 -3 34 103
use AND2X2  _1487_
timestamp 1563080643
transform 1 0 1412 0 1 1105
box -2 -3 34 103
use OAI21X1  _1538_
timestamp 1563080643
transform 1 0 1444 0 1 1105
box -2 -3 34 103
use OAI21X1  _1479_
timestamp 1563080643
transform -1 0 1508 0 1 1105
box -2 -3 34 103
use NAND2X1  _1534_
timestamp 1563080643
transform -1 0 1532 0 1 1105
box -2 -3 26 103
use INVX2  _1475_
timestamp 1563080643
transform -1 0 1548 0 1 1105
box -2 -3 18 103
use NAND2X1  _1488_
timestamp 1563080643
transform 1 0 1548 0 1 1105
box -2 -3 26 103
use INVX2  _1476_
timestamp 1563080643
transform 1 0 1572 0 1 1105
box -2 -3 18 103
use OAI22X1  _1478_
timestamp 1563080643
transform 1 0 1588 0 1 1105
box -2 -3 42 103
use DFFPOSX1  _1601_
timestamp 1563080643
transform 1 0 1628 0 1 1105
box -2 -3 98 103
use FILL  FILL_12_1
timestamp 1563080643
transform 1 0 1724 0 1 1105
box -2 -3 10 103
use INVX1  _1372_
timestamp 1563080643
transform 1 0 4 0 -1 1105
box -2 -3 18 103
use NAND3X1  _1039_
timestamp 1563080643
transform 1 0 20 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1373_
timestamp 1563080643
transform -1 0 76 0 -1 1105
box -2 -3 26 103
use NAND3X1  _1375_
timestamp 1563080643
transform -1 0 108 0 -1 1105
box -2 -3 34 103
use OR2X2  _1374_
timestamp 1563080643
transform -1 0 140 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1376_
timestamp 1563080643
transform -1 0 172 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_insert35
timestamp 1563080643
transform -1 0 196 0 -1 1105
box -2 -3 26 103
use OR2X2  _1407_
timestamp 1563080643
transform 1 0 196 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1410_
timestamp 1563080643
transform -1 0 260 0 -1 1105
box -2 -3 34 103
use INVX2  _1286_
timestamp 1563080643
transform -1 0 276 0 -1 1105
box -2 -3 18 103
use NAND3X1  _1296_
timestamp 1563080643
transform 1 0 276 0 -1 1105
box -2 -3 34 103
use NAND2X1  _1293_
timestamp 1563080643
transform 1 0 308 0 -1 1105
box -2 -3 26 103
use INVX1  _1292_
timestamp 1563080643
transform -1 0 348 0 -1 1105
box -2 -3 18 103
use NAND3X1  _1306_
timestamp 1563080643
transform -1 0 380 0 -1 1105
box -2 -3 34 103
use NAND3X1  _1386_
timestamp 1563080643
transform -1 0 412 0 -1 1105
box -2 -3 34 103
use OR2X2  _876_
timestamp 1563080643
transform 1 0 412 0 -1 1105
box -2 -3 34 103
use INVX1  _874_
timestamp 1563080643
transform -1 0 460 0 -1 1105
box -2 -3 18 103
use NAND2X1  _875_
timestamp 1563080643
transform -1 0 484 0 -1 1105
box -2 -3 26 103
use NAND3X1  _877_
timestamp 1563080643
transform -1 0 516 0 -1 1105
box -2 -3 34 103
use OR2X2  _790_
timestamp 1563080643
transform 1 0 516 0 -1 1105
box -2 -3 34 103
use NAND3X1  _793_
timestamp 1563080643
transform 1 0 548 0 -1 1105
box -2 -3 34 103
use NAND2X1  _792_
timestamp 1563080643
transform 1 0 580 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_0_0
timestamp 1563080643
transform -1 0 612 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1563080643
transform -1 0 620 0 -1 1105
box -2 -3 10 103
use NAND3X1  _798_
timestamp 1563080643
transform -1 0 652 0 -1 1105
box -2 -3 34 103
use NAND3X1  _878_
timestamp 1563080643
transform -1 0 684 0 -1 1105
box -2 -3 34 103
use NAND3X1  _848_
timestamp 1563080643
transform -1 0 716 0 -1 1105
box -2 -3 34 103
use INVX4  _1121_
timestamp 1563080643
transform 1 0 716 0 -1 1105
box -2 -3 26 103
use INVX2  _1120_
timestamp 1563080643
transform 1 0 740 0 -1 1105
box -2 -3 18 103
use INVX2  _788_
timestamp 1563080643
transform -1 0 772 0 -1 1105
box -2 -3 18 103
use NAND3X1  _888_
timestamp 1563080643
transform -1 0 804 0 -1 1105
box -2 -3 34 103
use NAND3X1  _808_
timestamp 1563080643
transform -1 0 836 0 -1 1105
box -2 -3 34 103
use NAND3X1  _839_
timestamp 1563080643
transform 1 0 836 0 -1 1105
box -2 -3 34 103
use NAND3X1  _917_
timestamp 1563080643
transform 1 0 868 0 -1 1105
box -2 -3 34 103
use NAND3X1  _927_
timestamp 1563080643
transform -1 0 932 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  _949_
timestamp 1563080643
transform 1 0 932 0 -1 1105
box -2 -3 98 103
use AND2X2  _1463_
timestamp 1563080643
transform -1 0 1060 0 -1 1105
box -2 -3 34 103
use AND2X2  _777_
timestamp 1563080643
transform 1 0 1060 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1563080643
transform -1 0 1100 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1563080643
transform -1 0 1108 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  _1605_
timestamp 1563080643
transform -1 0 1204 0 -1 1105
box -2 -3 98 103
use AND2X2  _1450_
timestamp 1563080643
transform -1 0 1236 0 -1 1105
box -2 -3 34 103
use AND2X2  _1532_
timestamp 1563080643
transform 1 0 1236 0 -1 1105
box -2 -3 34 103
use OAI22X1  _1533_
timestamp 1563080643
transform -1 0 1308 0 -1 1105
box -2 -3 42 103
use INVX1  _1473_
timestamp 1563080643
transform 1 0 1308 0 -1 1105
box -2 -3 18 103
use AOI22X1  _1474_
timestamp 1563080643
transform -1 0 1364 0 -1 1105
box -2 -3 42 103
use NAND2X1  _1469_
timestamp 1563080643
transform -1 0 1388 0 -1 1105
box -2 -3 26 103
use NAND2X1  _1481_
timestamp 1563080643
transform 1 0 1388 0 -1 1105
box -2 -3 26 103
use INVX1  _1467_
timestamp 1563080643
transform -1 0 1428 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  _1618_
timestamp 1563080643
transform 1 0 1428 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  _1614_
timestamp 1563080643
transform -1 0 1620 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  _785_
timestamp 1563080643
transform 1 0 1620 0 -1 1105
box -2 -3 98 103
use FILL  FILL_11_1
timestamp 1563080643
transform -1 0 1724 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1563080643
transform -1 0 1732 0 -1 1105
box -2 -3 10 103
use BUFX2  BUFX2_insert27
timestamp 1563080643
transform 1 0 4 0 1 905
box -2 -3 26 103
use INVX1  _1330_
timestamp 1563080643
transform 1 0 28 0 1 905
box -2 -3 18 103
use NAND2X1  _1331_
timestamp 1563080643
transform -1 0 68 0 1 905
box -2 -3 26 103
use OR2X2  _1329_
timestamp 1563080643
transform 1 0 68 0 1 905
box -2 -3 34 103
use NAND3X1  _1332_
timestamp 1563080643
transform -1 0 132 0 1 905
box -2 -3 34 103
use OR2X2  _1288_
timestamp 1563080643
transform 1 0 132 0 1 905
box -2 -3 34 103
use NAND2X1  _1290_
timestamp 1563080643
transform 1 0 164 0 1 905
box -2 -3 26 103
use INVX1  _1289_
timestamp 1563080643
transform 1 0 188 0 1 905
box -2 -3 18 103
use NAND3X1  _1291_
timestamp 1563080643
transform -1 0 236 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_insert39
timestamp 1563080643
transform 1 0 236 0 1 905
box -2 -3 26 103
use NAND3X1  _1415_
timestamp 1563080643
transform 1 0 260 0 1 905
box -2 -3 34 103
use NAND3X1  _1414_
timestamp 1563080643
transform 1 0 292 0 1 905
box -2 -3 34 103
use OR2X2  _1413_
timestamp 1563080643
transform -1 0 356 0 1 905
box -2 -3 34 103
use NAND3X1  _1425_
timestamp 1563080643
transform -1 0 388 0 1 905
box -2 -3 34 103
use INVX1  _832_
timestamp 1563080643
transform 1 0 388 0 1 905
box -2 -3 18 103
use NAND2X1  _833_
timestamp 1563080643
transform -1 0 428 0 1 905
box -2 -3 26 103
use OR2X2  _831_
timestamp 1563080643
transform 1 0 428 0 1 905
box -2 -3 34 103
use NAND3X1  _834_
timestamp 1563080643
transform -1 0 492 0 1 905
box -2 -3 34 103
use INVX1  _841_
timestamp 1563080643
transform 1 0 492 0 1 905
box -2 -3 18 103
use NAND2X1  _842_
timestamp 1563080643
transform -1 0 532 0 1 905
box -2 -3 26 103
use OR2X2  _840_
timestamp 1563080643
transform 1 0 532 0 1 905
box -2 -3 34 103
use NAND3X1  _843_
timestamp 1563080643
transform 1 0 564 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1563080643
transform -1 0 604 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1563080643
transform -1 0 612 0 1 905
box -2 -3 10 103
use INVX1  _791_
timestamp 1563080643
transform -1 0 628 0 1 905
box -2 -3 18 103
use INVX1  _1206_
timestamp 1563080643
transform 1 0 628 0 1 905
box -2 -3 18 103
use NAND2X1  _1207_
timestamp 1563080643
transform -1 0 668 0 1 905
box -2 -3 26 103
use OR2X2  _1208_
timestamp 1563080643
transform 1 0 668 0 1 905
box -2 -3 34 103
use NAND3X1  _1209_
timestamp 1563080643
transform -1 0 732 0 1 905
box -2 -3 34 103
use NAND3X1  _1210_
timestamp 1563080643
transform -1 0 764 0 1 905
box -2 -3 34 103
use OR2X2  _909_
timestamp 1563080643
transform 1 0 764 0 1 905
box -2 -3 34 103
use INVX1  _910_
timestamp 1563080643
transform 1 0 796 0 1 905
box -2 -3 18 103
use NAND3X1  _912_
timestamp 1563080643
transform 1 0 812 0 1 905
box -2 -3 34 103
use NAND2X1  _911_
timestamp 1563080643
transform -1 0 868 0 1 905
box -2 -3 26 103
use NAND3X1  _838_
timestamp 1563080643
transform 1 0 868 0 1 905
box -2 -3 34 103
use NAND3X1  _916_
timestamp 1563080643
transform 1 0 900 0 1 905
box -2 -3 34 103
use OR2X2  _915_
timestamp 1563080643
transform 1 0 932 0 1 905
box -2 -3 34 103
use NAND3X1  _849_
timestamp 1563080643
transform -1 0 996 0 1 905
box -2 -3 34 103
use AOI21X1  _1406_
timestamp 1563080643
transform 1 0 996 0 1 905
box -2 -3 34 103
use AOI21X1  _1445_
timestamp 1563080643
transform -1 0 1060 0 1 905
box -2 -3 34 103
use AOI21X1  _947_
timestamp 1563080643
transform 1 0 1060 0 1 905
box -2 -3 34 103
use AOI21X1  _908_
timestamp 1563080643
transform 1 0 1092 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1563080643
transform 1 0 1124 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1563080643
transform 1 0 1132 0 1 905
box -2 -3 10 103
use AOI21X1  _830_
timestamp 1563080643
transform 1 0 1140 0 1 905
box -2 -3 34 103
use DFFPOSX1  _1446_
timestamp 1563080643
transform 1 0 1172 0 1 905
box -2 -3 98 103
use DFFPOSX1  _950_
timestamp 1563080643
transform -1 0 1364 0 1 905
box -2 -3 98 103
use NAND2X1  _1471_
timestamp 1563080643
transform -1 0 1388 0 1 905
box -2 -3 26 103
use INVX1  _1468_
timestamp 1563080643
transform -1 0 1404 0 1 905
box -2 -3 18 103
use BUFX2  BUFX2_insert42
timestamp 1563080643
transform 1 0 1404 0 1 905
box -2 -3 26 103
use DFFPOSX1  _1615_
timestamp 1563080643
transform -1 0 1524 0 1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_insert45
timestamp 1563080643
transform -1 0 1596 0 1 905
box -2 -3 74 103
use DFFPOSX1  _1613_
timestamp 1563080643
transform 1 0 1596 0 1 905
box -2 -3 98 103
use AND2X2  _774_
timestamp 1563080643
transform -1 0 1724 0 1 905
box -2 -3 34 103
use FILL  FILL_10_1
timestamp 1563080643
transform 1 0 1724 0 1 905
box -2 -3 10 103
use INVX1  _957_
timestamp 1563080643
transform 1 0 4 0 -1 905
box -2 -3 18 103
use NAND2X1  _1041_
timestamp 1563080643
transform 1 0 20 0 -1 905
box -2 -3 26 103
use INVX1  _1040_
timestamp 1563080643
transform -1 0 60 0 -1 905
box -2 -3 18 103
use OR2X2  _1042_
timestamp 1563080643
transform 1 0 60 0 -1 905
box -2 -3 34 103
use NAND3X1  _1043_
timestamp 1563080643
transform -1 0 124 0 -1 905
box -2 -3 34 103
use NAND3X1  _1044_
timestamp 1563080643
transform -1 0 156 0 -1 905
box -2 -3 34 103
use INVX1  _1339_
timestamp 1563080643
transform 1 0 156 0 -1 905
box -2 -3 18 103
use NAND2X1  _1340_
timestamp 1563080643
transform 1 0 172 0 -1 905
box -2 -3 26 103
use OR2X2  _1335_
timestamp 1563080643
transform 1 0 196 0 -1 905
box -2 -3 34 103
use NAND3X1  _1337_
timestamp 1563080643
transform 1 0 228 0 -1 905
box -2 -3 34 103
use NAND3X1  _1336_
timestamp 1563080643
transform 1 0 260 0 -1 905
box -2 -3 34 103
use NAND3X1  _1341_
timestamp 1563080643
transform -1 0 324 0 -1 905
box -2 -3 34 103
use NAND2X1  _1412_
timestamp 1563080643
transform -1 0 348 0 -1 905
box -2 -3 26 103
use OR2X2  _1338_
timestamp 1563080643
transform -1 0 380 0 -1 905
box -2 -3 34 103
use NAND2X1  _1345_
timestamp 1563080643
transform 1 0 380 0 -1 905
box -2 -3 26 103
use NAND3X1  _1346_
timestamp 1563080643
transform 1 0 404 0 -1 905
box -2 -3 34 103
use NAND3X1  _1347_
timestamp 1563080643
transform 1 0 436 0 -1 905
box -2 -3 34 103
use INVX1  _1173_
timestamp 1563080643
transform 1 0 468 0 -1 905
box -2 -3 18 103
use NAND2X1  _1174_
timestamp 1563080643
transform 1 0 484 0 -1 905
box -2 -3 26 103
use OR2X2  _1172_
timestamp 1563080643
transform 1 0 508 0 -1 905
box -2 -3 34 103
use NAND3X1  _1175_
timestamp 1563080643
transform -1 0 572 0 -1 905
box -2 -3 34 103
use OR2X2  _1122_
timestamp 1563080643
transform 1 0 572 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1563080643
transform 1 0 604 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1563080643
transform 1 0 612 0 -1 905
box -2 -3 10 103
use INVX1  _1123_
timestamp 1563080643
transform 1 0 620 0 -1 905
box -2 -3 18 103
use BUFX2  BUFX2_insert18
timestamp 1563080643
transform 1 0 636 0 -1 905
box -2 -3 26 103
use NAND2X1  _1124_
timestamp 1563080643
transform 1 0 660 0 -1 905
box -2 -3 26 103
use NAND2X1  _847_
timestamp 1563080643
transform -1 0 708 0 -1 905
box -2 -3 26 103
use NAND3X1  _1125_
timestamp 1563080643
transform -1 0 740 0 -1 905
box -2 -3 34 103
use NAND3X1  _1130_
timestamp 1563080643
transform -1 0 772 0 -1 905
box -2 -3 34 103
use NAND3X1  _1171_
timestamp 1563080643
transform -1 0 804 0 -1 905
box -2 -3 34 103
use NAND3X1  _1249_
timestamp 1563080643
transform 1 0 804 0 -1 905
box -2 -3 34 103
use OR2X2  _837_
timestamp 1563080643
transform 1 0 836 0 -1 905
box -2 -3 34 103
use NAND2X1  _836_
timestamp 1563080643
transform 1 0 868 0 -1 905
box -2 -3 26 103
use NAND2X1  _914_
timestamp 1563080643
transform -1 0 916 0 -1 905
box -2 -3 26 103
use NAND3X1  _1220_
timestamp 1563080643
transform -1 0 948 0 -1 905
box -2 -3 34 103
use NAND3X1  _1140_
timestamp 1563080643
transform -1 0 980 0 -1 905
box -2 -3 34 103
use NAND3X1  _1259_
timestamp 1563080643
transform -1 0 1012 0 -1 905
box -2 -3 34 103
use DFFPOSX1  _1447_
timestamp 1563080643
transform 1 0 1012 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_1_0
timestamp 1563080643
transform -1 0 1116 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1563080643
transform -1 0 1124 0 -1 905
box -2 -3 10 103
use INVX2  _786_
timestamp 1563080643
transform -1 0 1140 0 -1 905
box -2 -3 18 103
use BUFX2  BUFX2_insert40
timestamp 1563080643
transform -1 0 1164 0 -1 905
box -2 -3 26 103
use AND2X2  _1462_
timestamp 1563080643
transform -1 0 1196 0 -1 905
box -2 -3 34 103
use DFFPOSX1  _948_
timestamp 1563080643
transform -1 0 1292 0 -1 905
box -2 -3 98 103
use AND2X2  _1451_
timestamp 1563080643
transform 1 0 1292 0 -1 905
box -2 -3 34 103
use DFFPOSX1  _1619_
timestamp 1563080643
transform 1 0 1324 0 -1 905
box -2 -3 98 103
use AOI21X1  _1535_
timestamp 1563080643
transform -1 0 1452 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_insert46
timestamp 1563080643
transform 1 0 1452 0 -1 905
box -2 -3 74 103
use DFFPOSX1  _1616_
timestamp 1563080643
transform -1 0 1620 0 -1 905
box -2 -3 98 103
use AND2X2  _1454_
timestamp 1563080643
transform 1 0 1620 0 -1 905
box -2 -3 34 103
use AND2X2  _1455_
timestamp 1563080643
transform -1 0 1684 0 -1 905
box -2 -3 34 103
use BUFX2  _780_
timestamp 1563080643
transform 1 0 1684 0 -1 905
box -2 -3 26 103
use NAND2X1  _1593_
timestamp 1563080643
transform -1 0 1732 0 -1 905
box -2 -3 26 103
use NAND2X1  _958_
timestamp 1563080643
transform -1 0 28 0 1 705
box -2 -3 26 103
use OR2X2  _956_
timestamp 1563080643
transform -1 0 60 0 1 705
box -2 -3 34 103
use BUFX2  BUFX2_insert26
timestamp 1563080643
transform 1 0 60 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_insert25
timestamp 1563080643
transform 1 0 84 0 1 705
box -2 -3 26 103
use INVX1  _1007_
timestamp 1563080643
transform -1 0 124 0 1 705
box -2 -3 18 103
use NAND2X1  _1008_
timestamp 1563080643
transform -1 0 148 0 1 705
box -2 -3 26 103
use OR2X2  _1003_
timestamp 1563080643
transform 1 0 148 0 1 705
box -2 -3 34 103
use NAND2X1  _1002_
timestamp 1563080643
transform 1 0 180 0 1 705
box -2 -3 26 103
use INVX1  _1001_
timestamp 1563080643
transform -1 0 220 0 1 705
box -2 -3 18 103
use NAND2X1  _999_
timestamp 1563080643
transform 1 0 220 0 1 705
box -2 -3 26 103
use INVX1  _998_
timestamp 1563080643
transform -1 0 260 0 1 705
box -2 -3 18 103
use INVX1  _1333_
timestamp 1563080643
transform 1 0 260 0 1 705
box -2 -3 18 103
use NAND2X1  _1334_
timestamp 1563080643
transform -1 0 300 0 1 705
box -2 -3 26 103
use OR2X2  _997_
timestamp 1563080643
transform -1 0 332 0 1 705
box -2 -3 34 103
use INVX1  _1411_
timestamp 1563080643
transform -1 0 348 0 1 705
box -2 -3 18 103
use INVX1  _1342_
timestamp 1563080643
transform -1 0 364 0 1 705
box -2 -3 18 103
use OAI21X1  _1344_
timestamp 1563080643
transform 1 0 364 0 1 705
box -2 -3 34 103
use INVX2  _1285_
timestamp 1563080643
transform -1 0 412 0 1 705
box -2 -3 18 103
use INVX1  _1164_
timestamp 1563080643
transform 1 0 412 0 1 705
box -2 -3 18 103
use NAND2X1  _1165_
timestamp 1563080643
transform -1 0 452 0 1 705
box -2 -3 26 103
use OR2X2  _1163_
timestamp 1563080643
transform 1 0 452 0 1 705
box -2 -3 34 103
use NAND3X1  _1166_
timestamp 1563080643
transform -1 0 516 0 1 705
box -2 -3 34 103
use OR2X2  _1128_
timestamp 1563080643
transform 1 0 516 0 1 705
box -2 -3 34 103
use BUFX2  BUFX2_insert17
timestamp 1563080643
transform -1 0 572 0 1 705
box -2 -3 26 103
use NAND3X1  _1129_
timestamp 1563080643
transform -1 0 604 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1563080643
transform -1 0 612 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1563080643
transform -1 0 620 0 1 705
box -2 -3 10 103
use NAND3X1  _1180_
timestamp 1563080643
transform -1 0 652 0 1 705
box -2 -3 34 103
use BUFX2  BUFX2_insert19
timestamp 1563080643
transform 1 0 652 0 1 705
box -2 -3 26 103
use NAND3X1  _1244_
timestamp 1563080643
transform -1 0 708 0 1 705
box -2 -3 34 103
use NAND3X1  _1170_
timestamp 1563080643
transform -1 0 740 0 1 705
box -2 -3 34 103
use OR2X2  _1169_
timestamp 1563080643
transform -1 0 772 0 1 705
box -2 -3 34 103
use OR2X2  _1247_
timestamp 1563080643
transform 1 0 772 0 1 705
box -2 -3 34 103
use NAND3X1  _1248_
timestamp 1563080643
transform 1 0 804 0 1 705
box -2 -3 34 103
use INVX1  _835_
timestamp 1563080643
transform 1 0 836 0 1 705
box -2 -3 18 103
use INVX1  _913_
timestamp 1563080643
transform 1 0 852 0 1 705
box -2 -3 18 103
use AND2X2  _1461_
timestamp 1563080643
transform -1 0 900 0 1 705
box -2 -3 34 103
use AND2X2  _1460_
timestamp 1563080643
transform 1 0 900 0 1 705
box -2 -3 34 103
use NAND3X1  _1181_
timestamp 1563080643
transform -1 0 964 0 1 705
box -2 -3 34 103
use AOI21X1  _1328_
timestamp 1563080643
transform 1 0 964 0 1 705
box -2 -3 34 103
use AOI21X1  _869_
timestamp 1563080643
transform 1 0 996 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_insert47
timestamp 1563080643
transform -1 0 1100 0 1 705
box -2 -3 74 103
use BUFX2  BUFX2_insert41
timestamp 1563080643
transform -1 0 1124 0 1 705
box -2 -3 26 103
use FILL  FILL_7_1_0
timestamp 1563080643
transform 1 0 1124 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1563080643
transform 1 0 1132 0 1 705
box -2 -3 10 103
use DFFPOSX1  _1448_
timestamp 1563080643
transform 1 0 1140 0 1 705
box -2 -3 98 103
use AND2X2  _1452_
timestamp 1563080643
transform 1 0 1236 0 1 705
box -2 -3 34 103
use DFFPOSX1  _1620_
timestamp 1563080643
transform 1 0 1268 0 1 705
box -2 -3 98 103
use AOI21X1  _1162_
timestamp 1563080643
transform 1 0 1364 0 1 705
box -2 -3 34 103
use BUFX2  BUFX2_insert44
timestamp 1563080643
transform 1 0 1396 0 1 705
box -2 -3 26 103
use INVX2  _1118_
timestamp 1563080643
transform 1 0 1420 0 1 705
box -2 -3 18 103
use AOI21X1  _1240_
timestamp 1563080643
transform 1 0 1436 0 1 705
box -2 -3 34 103
use AOI21X1  _1279_
timestamp 1563080643
transform 1 0 1468 0 1 705
box -2 -3 34 103
use AOI21X1  _1201_
timestamp 1563080643
transform -1 0 1532 0 1 705
box -2 -3 34 103
use DFFPOSX1  _1280_
timestamp 1563080643
transform 1 0 1532 0 1 705
box -2 -3 98 103
use DFFPOSX1  _782_
timestamp 1563080643
transform 1 0 1628 0 1 705
box -2 -3 98 103
use FILL  FILL_8_1
timestamp 1563080643
transform 1 0 1724 0 1 705
box -2 -3 10 103
use NAND3X1  _959_
timestamp 1563080643
transform -1 0 36 0 -1 705
box -2 -3 34 103
use INVX2  _954_
timestamp 1563080643
transform 1 0 36 0 -1 705
box -2 -3 18 103
use OR2X2  _1006_
timestamp 1563080643
transform 1 0 52 0 -1 705
box -2 -3 34 103
use NAND3X1  _1009_
timestamp 1563080643
transform 1 0 84 0 -1 705
box -2 -3 34 103
use NAND3X1  _1014_
timestamp 1563080643
transform 1 0 116 0 -1 705
box -2 -3 34 103
use NAND3X1  _1054_
timestamp 1563080643
transform -1 0 180 0 -1 705
box -2 -3 34 103
use NAND3X1  _1004_
timestamp 1563080643
transform 1 0 180 0 -1 705
box -2 -3 34 103
use NAND2X1  _1011_
timestamp 1563080643
transform -1 0 236 0 -1 705
box -2 -3 26 103
use NAND3X1  _1000_
timestamp 1563080643
transform -1 0 268 0 -1 705
box -2 -3 34 103
use OR2X2  _1075_
timestamp 1563080643
transform 1 0 268 0 -1 705
box -2 -3 34 103
use NAND3X1  _1078_
timestamp 1563080643
transform 1 0 300 0 -1 705
box -2 -3 34 103
use NAND2X1  _1077_
timestamp 1563080643
transform 1 0 332 0 -1 705
box -2 -3 26 103
use INVX1  _1076_
timestamp 1563080643
transform -1 0 372 0 -1 705
box -2 -3 18 103
use NAND2X1  _1343_
timestamp 1563080643
transform 1 0 372 0 -1 705
box -2 -3 26 103
use NAND2X1  _845_
timestamp 1563080643
transform -1 0 420 0 -1 705
box -2 -3 26 103
use INVX1  _844_
timestamp 1563080643
transform 1 0 420 0 -1 705
box -2 -3 18 103
use OAI21X1  _846_
timestamp 1563080643
transform 1 0 436 0 -1 705
box -2 -3 34 103
use NAND2X1  _1177_
timestamp 1563080643
transform -1 0 492 0 -1 705
box -2 -3 26 103
use INVX1  _1176_
timestamp 1563080643
transform 1 0 492 0 -1 705
box -2 -3 18 103
use OAI21X1  _1178_
timestamp 1563080643
transform -1 0 540 0 -1 705
box -2 -3 34 103
use INVX1  _1126_
timestamp 1563080643
transform 1 0 540 0 -1 705
box -2 -3 18 103
use NAND2X1  _1127_
timestamp 1563080643
transform 1 0 556 0 -1 705
box -2 -3 26 103
use NAND2X1  _1179_
timestamp 1563080643
transform -1 0 604 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_0_0
timestamp 1563080643
transform 1 0 604 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1563080643
transform 1 0 612 0 -1 705
box -2 -3 10 103
use INVX1  _1242_
timestamp 1563080643
transform 1 0 620 0 -1 705
box -2 -3 18 103
use NAND2X1  _1243_
timestamp 1563080643
transform -1 0 660 0 -1 705
box -2 -3 26 103
use NAND2X1  _1168_
timestamp 1563080643
transform 1 0 660 0 -1 705
box -2 -3 26 103
use INVX1  _1167_
timestamp 1563080643
transform -1 0 700 0 -1 705
box -2 -3 18 103
use OR2X2  _1241_
timestamp 1563080643
transform -1 0 732 0 -1 705
box -2 -3 34 103
use INVX1  _1245_
timestamp 1563080643
transform 1 0 732 0 -1 705
box -2 -3 18 103
use NAND2X1  _1246_
timestamp 1563080643
transform -1 0 772 0 -1 705
box -2 -3 26 103
use AND2X2  _1458_
timestamp 1563080643
transform 1 0 772 0 -1 705
box -2 -3 34 103
use AND2X2  _1459_
timestamp 1563080643
transform 1 0 804 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1116_
timestamp 1563080643
transform 1 0 836 0 -1 705
box -2 -3 98 103
use AOI21X1  _1367_
timestamp 1563080643
transform 1 0 932 0 -1 705
box -2 -3 34 103
use INVX2  _1284_
timestamp 1563080643
transform 1 0 964 0 -1 705
box -2 -3 18 103
use AND2X2  _1465_
timestamp 1563080643
transform 1 0 980 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1608_
timestamp 1563080643
transform 1 0 1012 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_1_0
timestamp 1563080643
transform 1 0 1108 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1563080643
transform 1 0 1116 0 -1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_insert50
timestamp 1563080643
transform 1 0 1124 0 -1 705
box -2 -3 74 103
use DFFPOSX1  _1449_
timestamp 1563080643
transform 1 0 1196 0 -1 705
box -2 -3 98 103
use AND2X2  _1453_
timestamp 1563080643
transform -1 0 1324 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1282_
timestamp 1563080643
transform 1 0 1324 0 -1 705
box -2 -3 98 103
use AND2X2  _1456_
timestamp 1563080643
transform 1 0 1420 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1283_
timestamp 1563080643
transform -1 0 1548 0 -1 705
box -2 -3 98 103
use AND2X2  _1457_
timestamp 1563080643
transform 1 0 1548 0 -1 705
box -2 -3 34 103
use DFFPOSX1  _1281_
timestamp 1563080643
transform 1 0 1580 0 -1 705
box -2 -3 98 103
use BUFX2  _781_
timestamp 1563080643
transform 1 0 1676 0 -1 705
box -2 -3 26 103
use BUFX2  _778_
timestamp 1563080643
transform 1 0 1700 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1563080643
transform -1 0 1732 0 -1 705
box -2 -3 10 103
use NAND3X1  _964_
timestamp 1563080643
transform -1 0 36 0 1 505
box -2 -3 34 103
use NAND3X1  _974_
timestamp 1563080643
transform -1 0 68 0 1 505
box -2 -3 34 103
use INVX2  _953_
timestamp 1563080643
transform 1 0 68 0 1 505
box -2 -3 18 103
use INVX1  _1010_
timestamp 1563080643
transform -1 0 100 0 1 505
box -2 -3 18 103
use OAI21X1  _1012_
timestamp 1563080643
transform 1 0 100 0 1 505
box -2 -3 34 103
use NAND3X1  _1015_
timestamp 1563080643
transform -1 0 164 0 1 505
box -2 -3 34 103
use NAND3X1  _1005_
timestamp 1563080643
transform -1 0 196 0 1 505
box -2 -3 34 103
use NAND3X1  _1093_
timestamp 1563080643
transform 1 0 196 0 1 505
box -2 -3 34 103
use NAND3X1  _1083_
timestamp 1563080643
transform 1 0 228 0 1 505
box -2 -3 34 103
use NAND3X1  _1082_
timestamp 1563080643
transform 1 0 260 0 1 505
box -2 -3 34 103
use OR2X2  _1081_
timestamp 1563080643
transform -1 0 324 0 1 505
box -2 -3 34 103
use AOI21X1  _1113_
timestamp 1563080643
transform 1 0 324 0 1 505
box -2 -3 34 103
use AOI21X1  _1074_
timestamp 1563080643
transform 1 0 356 0 1 505
box -2 -3 34 103
use AOI21X1  _1035_
timestamp 1563080643
transform 1 0 388 0 1 505
box -2 -3 34 103
use AOI21X1  _996_
timestamp 1563080643
transform 1 0 420 0 1 505
box -2 -3 34 103
use INVX2  _952_
timestamp 1563080643
transform -1 0 468 0 1 505
box -2 -3 18 103
use DFFPOSX1  _1114_
timestamp 1563080643
transform 1 0 468 0 1 505
box -2 -3 98 103
use NAND3X1  _1405_
timestamp 1563080643
transform -1 0 596 0 1 505
box -2 -3 34 103
use FILL  FILL_5_0_0
timestamp 1563080643
transform 1 0 596 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1563080643
transform 1 0 604 0 1 505
box -2 -3 10 103
use DFFPOSX1  _1115_
timestamp 1563080643
transform 1 0 612 0 1 505
box -2 -3 98 103
use NAND3X1  _1366_
timestamp 1563080643
transform -1 0 740 0 1 505
box -2 -3 34 103
use NAND3X1  _1327_
timestamp 1563080643
transform -1 0 772 0 1 505
box -2 -3 34 103
use NAND3X1  _1444_
timestamp 1563080643
transform 1 0 772 0 1 505
box -2 -3 34 103
use DFFPOSX1  _1117_
timestamp 1563080643
transform 1 0 804 0 1 505
box -2 -3 98 103
use DFFPOSX1  _951_
timestamp 1563080643
transform 1 0 900 0 1 505
box -2 -3 98 103
use INVX2  _787_
timestamp 1563080643
transform -1 0 1012 0 1 505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_insert49
timestamp 1563080643
transform -1 0 1084 0 1 505
box -2 -3 74 103
use NAND3X1  _829_
timestamp 1563080643
transform -1 0 1116 0 1 505
box -2 -3 34 103
use FILL  FILL_5_1_0
timestamp 1563080643
transform -1 0 1124 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1563080643
transform -1 0 1132 0 1 505
box -2 -3 10 103
use BUFX2  BUFX2_insert21
timestamp 1563080643
transform -1 0 1156 0 1 505
box -2 -3 26 103
use NAND3X1  _868_
timestamp 1563080643
transform 1 0 1156 0 1 505
box -2 -3 34 103
use INVX1  _815_
timestamp 1563080643
transform 1 0 1188 0 1 505
box -2 -3 18 103
use NAND2X1  _816_
timestamp 1563080643
transform -1 0 1228 0 1 505
box -2 -3 26 103
use BUFX2  BUFX2_insert23
timestamp 1563080643
transform 1 0 1228 0 1 505
box -2 -3 26 103
use NAND2X1  _855_
timestamp 1563080643
transform 1 0 1252 0 1 505
box -2 -3 26 103
use INVX1  _854_
timestamp 1563080643
transform -1 0 1292 0 1 505
box -2 -3 18 103
use NAND2X1  _852_
timestamp 1563080643
transform 1 0 1292 0 1 505
box -2 -3 26 103
use INVX1  _851_
timestamp 1563080643
transform -1 0 1332 0 1 505
box -2 -3 18 103
use INVX2  _1119_
timestamp 1563080643
transform -1 0 1348 0 1 505
box -2 -3 18 103
use NAND3X1  _1161_
timestamp 1563080643
transform 1 0 1348 0 1 505
box -2 -3 34 103
use OR2X2  _1149_
timestamp 1563080643
transform 1 0 1380 0 1 505
box -2 -3 34 103
use NAND3X1  _1151_
timestamp 1563080643
transform 1 0 1412 0 1 505
box -2 -3 34 103
use NAND3X1  _1150_
timestamp 1563080643
transform 1 0 1444 0 1 505
box -2 -3 34 103
use NAND2X1  _1148_
timestamp 1563080643
transform 1 0 1476 0 1 505
box -2 -3 26 103
use INVX1  _1147_
timestamp 1563080643
transform -1 0 1516 0 1 505
box -2 -3 18 103
use NAND2X1  _1237_
timestamp 1563080643
transform 1 0 1516 0 1 505
box -2 -3 26 103
use NAND2X1  _1184_
timestamp 1563080643
transform 1 0 1540 0 1 505
box -2 -3 26 103
use INVX1  _1183_
timestamp 1563080643
transform 1 0 1564 0 1 505
box -2 -3 18 103
use INVX1  _1234_
timestamp 1563080643
transform 1 0 1580 0 1 505
box -2 -3 18 103
use OAI21X1  _1236_
timestamp 1563080643
transform 1 0 1596 0 1 505
box -2 -3 34 103
use AND2X2  _776_
timestamp 1563080643
transform 1 0 1628 0 1 505
box -2 -3 34 103
use INVX1  _1186_
timestamp 1563080643
transform 1 0 1660 0 1 505
box -2 -3 18 103
use NAND2X1  _1187_
timestamp 1563080643
transform -1 0 1700 0 1 505
box -2 -3 26 103
use BUFX2  _779_
timestamp 1563080643
transform 1 0 1700 0 1 505
box -2 -3 26 103
use FILL  FILL_6_1
timestamp 1563080643
transform 1 0 1724 0 1 505
box -2 -3 10 103
use NAND3X1  _963_
timestamp 1563080643
transform 1 0 4 0 -1 505
box -2 -3 34 103
use OR2X2  _962_
timestamp 1563080643
transform -1 0 68 0 -1 505
box -2 -3 34 103
use INVX1  _960_
timestamp 1563080643
transform -1 0 84 0 -1 505
box -2 -3 18 103
use NAND2X1  _961_
timestamp 1563080643
transform -1 0 108 0 -1 505
box -2 -3 26 103
use NAND2X1  _1013_
timestamp 1563080643
transform 1 0 108 0 -1 505
box -2 -3 26 103
use INVX1  _1079_
timestamp 1563080643
transform 1 0 132 0 -1 505
box -2 -3 18 103
use NAND2X1  _1080_
timestamp 1563080643
transform 1 0 148 0 -1 505
box -2 -3 26 103
use NAND3X1  _984_
timestamp 1563080643
transform 1 0 172 0 -1 505
box -2 -3 34 103
use OR2X2  _983_
timestamp 1563080643
transform -1 0 236 0 -1 505
box -2 -3 34 103
use NAND3X1  _1034_
timestamp 1563080643
transform 1 0 236 0 -1 505
box -2 -3 34 103
use NAND2X1  _982_
timestamp 1563080643
transform 1 0 268 0 -1 505
box -2 -3 26 103
use NAND3X1  _1024_
timestamp 1563080643
transform 1 0 292 0 -1 505
box -2 -3 34 103
use NAND3X1  _1023_
timestamp 1563080643
transform 1 0 324 0 -1 505
box -2 -3 34 103
use OR2X2  _1022_
timestamp 1563080643
transform -1 0 388 0 -1 505
box -2 -3 34 103
use NAND2X1  _1018_
timestamp 1563080643
transform 1 0 388 0 -1 505
box -2 -3 26 103
use NAND2X1  _1069_
timestamp 1563080643
transform 1 0 412 0 -1 505
box -2 -3 26 103
use NAND2X1  _1021_
timestamp 1563080643
transform 1 0 436 0 -1 505
box -2 -3 26 103
use INVX1  _1017_
timestamp 1563080643
transform -1 0 476 0 -1 505
box -2 -3 18 103
use INVX1  _1020_
timestamp 1563080643
transform -1 0 492 0 -1 505
box -2 -3 18 103
use INVX1  _1349_
timestamp 1563080643
transform 1 0 492 0 -1 505
box -2 -3 18 103
use NAND2X1  _1350_
timestamp 1563080643
transform -1 0 532 0 -1 505
box -2 -3 26 103
use OR2X2  _1309_
timestamp 1563080643
transform 1 0 532 0 -1 505
box -2 -3 34 103
use NAND3X1  _1312_
timestamp 1563080643
transform -1 0 596 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1563080643
transform 1 0 596 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1563080643
transform 1 0 604 0 -1 505
box -2 -3 10 103
use OR2X2  _1348_
timestamp 1563080643
transform 1 0 612 0 -1 505
box -2 -3 34 103
use NAND3X1  _1351_
timestamp 1563080643
transform -1 0 676 0 -1 505
box -2 -3 34 103
use NAND3X1  _1317_
timestamp 1563080643
transform 1 0 676 0 -1 505
box -2 -3 34 103
use NAND3X1  _1355_
timestamp 1563080643
transform 1 0 708 0 -1 505
box -2 -3 34 103
use OR2X2  _1354_
timestamp 1563080643
transform -1 0 772 0 -1 505
box -2 -3 34 103
use NAND2X1  _1353_
timestamp 1563080643
transform 1 0 772 0 -1 505
box -2 -3 26 103
use INVX1  _1352_
timestamp 1563080643
transform 1 0 796 0 -1 505
box -2 -3 18 103
use NAND2X1  _1401_
timestamp 1563080643
transform -1 0 836 0 -1 505
box -2 -3 26 103
use NAND3X1  _1316_
timestamp 1563080643
transform 1 0 836 0 -1 505
box -2 -3 34 103
use OR2X2  _1315_
timestamp 1563080643
transform -1 0 900 0 -1 505
box -2 -3 34 103
use NAND2X1  _1314_
timestamp 1563080643
transform 1 0 900 0 -1 505
box -2 -3 26 103
use INVX1  _981_
timestamp 1563080643
transform -1 0 940 0 -1 505
box -2 -3 18 103
use INVX1  _1313_
timestamp 1563080643
transform -1 0 956 0 -1 505
box -2 -3 18 103
use NAND3X1  _906_
timestamp 1563080643
transform -1 0 988 0 -1 505
box -2 -3 34 103
use NAND3X1  _907_
timestamp 1563080643
transform 1 0 988 0 -1 505
box -2 -3 34 103
use NAND2X1  _905_
timestamp 1563080643
transform -1 0 1044 0 -1 505
box -2 -3 26 103
use NAND2X1  _903_
timestamp 1563080643
transform 1 0 1044 0 -1 505
box -2 -3 26 103
use OAI21X1  _904_
timestamp 1563080643
transform -1 0 1100 0 -1 505
box -2 -3 34 103
use INVX1  _902_
timestamp 1563080643
transform -1 0 1116 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_1_0
timestamp 1563080643
transform 1 0 1116 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1563080643
transform 1 0 1124 0 -1 505
box -2 -3 10 103
use INVX4  _810_
timestamp 1563080643
transform 1 0 1132 0 -1 505
box -2 -3 26 103
use NAND3X1  _818_
timestamp 1563080643
transform 1 0 1156 0 -1 505
box -2 -3 34 103
use OR2X2  _817_
timestamp 1563080643
transform -1 0 1220 0 -1 505
box -2 -3 34 103
use NAND3X1  _858_
timestamp 1563080643
transform 1 0 1220 0 -1 505
box -2 -3 34 103
use NAND3X1  _857_
timestamp 1563080643
transform 1 0 1252 0 -1 505
box -2 -3 34 103
use NAND3X1  _853_
timestamp 1563080643
transform 1 0 1284 0 -1 505
box -2 -3 34 103
use OR2X2  _856_
timestamp 1563080643
transform -1 0 1348 0 -1 505
box -2 -3 34 103
use OR2X2  _850_
timestamp 1563080643
transform 1 0 1348 0 -1 505
box -2 -3 34 103
use OR2X2  _1143_
timestamp 1563080643
transform 1 0 1380 0 -1 505
box -2 -3 34 103
use NAND3X1  _1146_
timestamp 1563080643
transform 1 0 1412 0 -1 505
box -2 -3 34 103
use NAND2X1  _1145_
timestamp 1563080643
transform -1 0 1468 0 -1 505
box -2 -3 26 103
use NAND3X1  _1239_
timestamp 1563080643
transform 1 0 1468 0 -1 505
box -2 -3 34 103
use NAND3X1  _1238_
timestamp 1563080643
transform 1 0 1500 0 -1 505
box -2 -3 34 103
use OR2X2  _1182_
timestamp 1563080643
transform 1 0 1532 0 -1 505
box -2 -3 34 103
use NAND3X1  _1185_
timestamp 1563080643
transform -1 0 1596 0 -1 505
box -2 -3 34 103
use NAND2X1  _1235_
timestamp 1563080643
transform 1 0 1596 0 -1 505
box -2 -3 26 103
use NAND3X1  _1190_
timestamp 1563080643
transform 1 0 1620 0 -1 505
box -2 -3 34 103
use NAND3X1  _1189_
timestamp 1563080643
transform -1 0 1684 0 -1 505
box -2 -3 34 103
use OR2X2  _1188_
timestamp 1563080643
transform -1 0 1716 0 -1 505
box -2 -3 34 103
use FILL  FILL_5_1
timestamp 1563080643
transform -1 0 1724 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1563080643
transform -1 0 1732 0 -1 505
box -2 -3 10 103
use NAND3X1  _980_
timestamp 1563080643
transform -1 0 36 0 1 305
box -2 -3 34 103
use NAND3X1  _985_
timestamp 1563080643
transform -1 0 68 0 1 305
box -2 -3 34 103
use NAND3X1  _995_
timestamp 1563080643
transform 1 0 68 0 1 305
box -2 -3 34 103
use NAND3X1  _1112_
timestamp 1563080643
transform -1 0 132 0 1 305
box -2 -3 34 103
use NAND3X1  _1073_
timestamp 1563080643
transform -1 0 164 0 1 305
box -2 -3 34 103
use NAND3X1  _1072_
timestamp 1563080643
transform 1 0 164 0 1 305
box -2 -3 34 103
use NAND2X1  _1071_
timestamp 1563080643
transform 1 0 196 0 1 305
box -2 -3 26 103
use NAND3X1  _1067_
timestamp 1563080643
transform 1 0 220 0 1 305
box -2 -3 34 103
use OR2X2  _1016_
timestamp 1563080643
transform -1 0 284 0 1 305
box -2 -3 34 103
use NAND3X1  _1019_
timestamp 1563080643
transform 1 0 284 0 1 305
box -2 -3 34 103
use OR2X2  _1064_
timestamp 1563080643
transform -1 0 348 0 1 305
box -2 -3 34 103
use NAND2X1  _1066_
timestamp 1563080643
transform 1 0 348 0 1 305
box -2 -3 26 103
use INVX1  _1065_
timestamp 1563080643
transform -1 0 388 0 1 305
box -2 -3 18 103
use OAI21X1  _1070_
timestamp 1563080643
transform -1 0 420 0 1 305
box -2 -3 34 103
use INVX1  _1068_
timestamp 1563080643
transform -1 0 436 0 1 305
box -2 -3 18 103
use OR2X2  _1396_
timestamp 1563080643
transform 1 0 436 0 1 305
box -2 -3 34 103
use NAND3X1  _1399_
timestamp 1563080643
transform -1 0 500 0 1 305
box -2 -3 34 103
use INVX1  _1310_
timestamp 1563080643
transform 1 0 500 0 1 305
box -2 -3 18 103
use NAND2X1  _1311_
timestamp 1563080643
transform -1 0 540 0 1 305
box -2 -3 26 103
use NAND3X1  _1404_
timestamp 1563080643
transform -1 0 572 0 1 305
box -2 -3 34 103
use NAND2X1  _1403_
timestamp 1563080643
transform -1 0 596 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1563080643
transform 1 0 596 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1563080643
transform 1 0 604 0 1 305
box -2 -3 10 103
use INVX2  _1307_
timestamp 1563080643
transform 1 0 612 0 1 305
box -2 -3 18 103
use NAND3X1  _1443_
timestamp 1563080643
transform -1 0 660 0 1 305
box -2 -3 34 103
use NAND3X1  _1365_
timestamp 1563080643
transform -1 0 692 0 1 305
box -2 -3 34 103
use NAND3X1  _1356_
timestamp 1563080643
transform 1 0 692 0 1 305
box -2 -3 34 103
use NAND3X1  _1326_
timestamp 1563080643
transform -1 0 756 0 1 305
box -2 -3 34 103
use OAI21X1  _1402_
timestamp 1563080643
transform -1 0 788 0 1 305
box -2 -3 34 103
use INVX1  _1400_
timestamp 1563080643
transform -1 0 804 0 1 305
box -2 -3 18 103
use INVX4  _1308_
timestamp 1563080643
transform -1 0 828 0 1 305
box -2 -3 26 103
use INVX1  _812_
timestamp 1563080643
transform 1 0 828 0 1 305
box -2 -3 18 103
use NAND2X1  _813_
timestamp 1563080643
transform -1 0 868 0 1 305
box -2 -3 26 103
use INVX1  _899_
timestamp 1563080643
transform 1 0 868 0 1 305
box -2 -3 18 103
use NAND2X1  _900_
timestamp 1563080643
transform 1 0 884 0 1 305
box -2 -3 26 103
use OR2X2  _898_
timestamp 1563080643
transform 1 0 908 0 1 305
box -2 -3 34 103
use NAND3X1  _901_
timestamp 1563080643
transform -1 0 972 0 1 305
box -2 -3 34 103
use NAND3X1  _814_
timestamp 1563080643
transform -1 0 1004 0 1 305
box -2 -3 34 103
use OR2X2  _811_
timestamp 1563080643
transform -1 0 1036 0 1 305
box -2 -3 34 103
use INVX1  _1153_
timestamp 1563080643
transform 1 0 1036 0 1 305
box -2 -3 18 103
use NAND3X1  _946_
timestamp 1563080643
transform -1 0 1084 0 1 305
box -2 -3 34 103
use NAND3X1  _819_
timestamp 1563080643
transform 1 0 1084 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1563080643
transform 1 0 1116 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1563080643
transform 1 0 1124 0 1 305
box -2 -3 10 103
use OR2X2  _937_
timestamp 1563080643
transform 1 0 1132 0 1 305
box -2 -3 34 103
use NAND3X1  _940_
timestamp 1563080643
transform -1 0 1196 0 1 305
box -2 -3 34 103
use NAND3X1  _945_
timestamp 1563080643
transform 1 0 1196 0 1 305
box -2 -3 34 103
use INVX2  _809_
timestamp 1563080643
transform 1 0 1228 0 1 305
box -2 -3 18 103
use NAND3X1  _867_
timestamp 1563080643
transform 1 0 1244 0 1 305
box -2 -3 34 103
use INVX1  _1144_
timestamp 1563080643
transform 1 0 1276 0 1 305
box -2 -3 18 103
use OR2X2  _1269_
timestamp 1563080643
transform 1 0 1292 0 1 305
box -2 -3 34 103
use INVX1  _1270_
timestamp 1563080643
transform 1 0 1324 0 1 305
box -2 -3 18 103
use NAND2X1  _1154_
timestamp 1563080643
transform -1 0 1364 0 1 305
box -2 -3 26 103
use NAND3X1  _1160_
timestamp 1563080643
transform 1 0 1364 0 1 305
box -2 -3 34 103
use NAND2X1  _1271_
timestamp 1563080643
transform -1 0 1420 0 1 305
box -2 -3 26 103
use NAND3X1  _1272_
timestamp 1563080643
transform -1 0 1452 0 1 305
box -2 -3 34 103
use NAND3X1  _1277_
timestamp 1563080643
transform 1 0 1452 0 1 305
box -2 -3 34 103
use NAND3X1  _1278_
timestamp 1563080643
transform -1 0 1516 0 1 305
box -2 -3 34 103
use INVX2  _1141_
timestamp 1563080643
transform -1 0 1532 0 1 305
box -2 -3 18 103
use NAND3X1  _1199_
timestamp 1563080643
transform 1 0 1532 0 1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert6
timestamp 1563080643
transform -1 0 1588 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert9
timestamp 1563080643
transform -1 0 1612 0 1 305
box -2 -3 26 103
use NAND3X1  _1200_
timestamp 1563080643
transform 1 0 1612 0 1 305
box -2 -3 34 103
use NAND3X1  _1233_
timestamp 1563080643
transform 1 0 1644 0 1 305
box -2 -3 34 103
use INVX1  _1231_
timestamp 1563080643
transform 1 0 1676 0 1 305
box -2 -3 18 103
use NAND2X1  _1232_
timestamp 1563080643
transform -1 0 1716 0 1 305
box -2 -3 26 103
use FILL  FILL_4_1
timestamp 1563080643
transform 1 0 1716 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1563080643
transform 1 0 1724 0 1 305
box -2 -3 10 103
use INVX1  _978_
timestamp 1563080643
transform 1 0 4 0 -1 305
box -2 -3 18 103
use NAND2X1  _979_
timestamp 1563080643
transform -1 0 44 0 -1 305
box -2 -3 26 103
use OR2X2  _977_
timestamp 1563080643
transform -1 0 76 0 -1 305
box -2 -3 34 103
use NAND3X1  _994_
timestamp 1563080643
transform -1 0 108 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert10
timestamp 1563080643
transform -1 0 132 0 -1 305
box -2 -3 26 103
use NAND3X1  _1063_
timestamp 1563080643
transform 1 0 132 0 -1 305
box -2 -3 34 103
use NAND3X1  _1102_
timestamp 1563080643
transform 1 0 164 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert14
timestamp 1563080643
transform 1 0 196 0 -1 305
box -2 -3 26 103
use NAND3X1  _989_
timestamp 1563080643
transform 1 0 220 0 -1 305
box -2 -3 34 103
use OR2X2  _986_
timestamp 1563080643
transform -1 0 284 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert11
timestamp 1563080643
transform 1 0 284 0 -1 305
box -2 -3 26 103
use NAND2X1  _988_
timestamp 1563080643
transform 1 0 308 0 -1 305
box -2 -3 26 103
use NAND3X1  _1058_
timestamp 1563080643
transform 1 0 332 0 -1 305
box -2 -3 34 103
use OR2X2  _1055_
timestamp 1563080643
transform -1 0 396 0 -1 305
box -2 -3 34 103
use INVX1  _987_
timestamp 1563080643
transform -1 0 412 0 -1 305
box -2 -3 18 103
use INVX1  _1391_
timestamp 1563080643
transform 1 0 412 0 -1 305
box -2 -3 18 103
use NAND2X1  _1392_
timestamp 1563080643
transform -1 0 452 0 -1 305
box -2 -3 26 103
use INVX1  _1397_
timestamp 1563080643
transform 1 0 452 0 -1 305
box -2 -3 18 103
use NAND2X1  _1398_
timestamp 1563080643
transform -1 0 492 0 -1 305
box -2 -3 26 103
use OR2X2  _1393_
timestamp 1563080643
transform 1 0 492 0 -1 305
box -2 -3 34 103
use NAND3X1  _1394_
timestamp 1563080643
transform -1 0 556 0 -1 305
box -2 -3 34 103
use NAND3X1  _1395_
timestamp 1563080643
transform -1 0 588 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert4
timestamp 1563080643
transform -1 0 612 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_0_0
timestamp 1563080643
transform -1 0 620 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1563080643
transform -1 0 628 0 -1 305
box -2 -3 10 103
use NAND2X1  _1442_
timestamp 1563080643
transform -1 0 652 0 -1 305
box -2 -3 26 103
use NAND2X1  _1364_
timestamp 1563080643
transform -1 0 676 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert0
timestamp 1563080643
transform -1 0 700 0 -1 305
box -2 -3 26 103
use OR2X2  _1357_
timestamp 1563080643
transform 1 0 700 0 -1 305
box -2 -3 34 103
use NAND3X1  _1360_
timestamp 1563080643
transform 1 0 732 0 -1 305
box -2 -3 34 103
use NAND2X1  _1325_
timestamp 1563080643
transform -1 0 788 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert3
timestamp 1563080643
transform -1 0 812 0 -1 305
box -2 -3 26 103
use NAND3X1  _1434_
timestamp 1563080643
transform 1 0 812 0 -1 305
box -2 -3 34 103
use OR2X2  _820_
timestamp 1563080643
transform 1 0 844 0 -1 305
box -2 -3 34 103
use INVX1  _1225_
timestamp 1563080643
transform 1 0 876 0 -1 305
box -2 -3 18 103
use NAND2X1  _822_
timestamp 1563080643
transform 1 0 892 0 -1 305
box -2 -3 26 103
use INVX1  _821_
timestamp 1563080643
transform -1 0 932 0 -1 305
box -2 -3 18 103
use NAND3X1  _823_
timestamp 1563080643
transform -1 0 964 0 -1 305
box -2 -3 34 103
use NAND3X1  _828_
timestamp 1563080643
transform -1 0 996 0 -1 305
box -2 -3 34 103
use NAND3X1  _897_
timestamp 1563080643
transform 1 0 996 0 -1 305
box -2 -3 34 103
use INVX1  _938_
timestamp 1563080643
transform 1 0 1028 0 -1 305
box -2 -3 18 103
use NAND2X1  _939_
timestamp 1563080643
transform -1 0 1068 0 -1 305
box -2 -3 26 103
use NAND3X1  _936_
timestamp 1563080643
transform 1 0 1068 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_insert20
timestamp 1563080643
transform -1 0 1124 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_1_0
timestamp 1563080643
transform -1 0 1132 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1563080643
transform -1 0 1140 0 -1 305
box -2 -3 10 103
use NAND2X1  _1226_
timestamp 1563080643
transform -1 0 1164 0 -1 305
box -2 -3 26 103
use NAND2X1  _944_
timestamp 1563080643
transform -1 0 1188 0 -1 305
box -2 -3 26 103
use OR2X2  _1227_
timestamp 1563080643
transform 1 0 1188 0 -1 305
box -2 -3 34 103
use NAND3X1  _1228_
timestamp 1563080643
transform -1 0 1252 0 -1 305
box -2 -3 34 103
use NAND2X1  _866_
timestamp 1563080643
transform 1 0 1252 0 -1 305
box -2 -3 26 103
use OR2X2  _1221_
timestamp 1563080643
transform 1 0 1276 0 -1 305
box -2 -3 34 103
use NAND3X1  _1224_
timestamp 1563080643
transform -1 0 1340 0 -1 305
box -2 -3 34 103
use NAND3X1  _1229_
timestamp 1563080643
transform 1 0 1340 0 -1 305
box -2 -3 34 103
use NAND2X1  _1159_
timestamp 1563080643
transform 1 0 1372 0 -1 305
box -2 -3 26 103
use OR2X2  _1191_
timestamp 1563080643
transform 1 0 1396 0 -1 305
box -2 -3 34 103
use NAND3X1  _1194_
timestamp 1563080643
transform -1 0 1460 0 -1 305
box -2 -3 34 103
use INVX4  _1142_
timestamp 1563080643
transform -1 0 1484 0 -1 305
box -2 -3 26 103
use NAND2X1  _1276_
timestamp 1563080643
transform 1 0 1484 0 -1 305
box -2 -3 26 103
use NAND3X1  _1268_
timestamp 1563080643
transform 1 0 1508 0 -1 305
box -2 -3 34 103
use NAND2X1  _1198_
timestamp 1563080643
transform 1 0 1540 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_insert8
timestamp 1563080643
transform -1 0 1588 0 -1 305
box -2 -3 26 103
use DFFPOSX1  _783_
timestamp 1563080643
transform 1 0 1588 0 -1 305
box -2 -3 98 103
use OR2X2  _1230_
timestamp 1563080643
transform 1 0 1684 0 -1 305
box -2 -3 34 103
use FILL  FILL_3_1
timestamp 1563080643
transform -1 0 1724 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1563080643
transform -1 0 1732 0 -1 305
box -2 -3 10 103
use INVX4  _976_
timestamp 1563080643
transform -1 0 28 0 1 105
box -2 -3 26 103
use NAND3X1  _1106_
timestamp 1563080643
transform -1 0 60 0 1 105
box -2 -3 34 103
use OR2X2  _1103_
timestamp 1563080643
transform -1 0 92 0 1 105
box -2 -3 34 103
use NAND3X1  _1111_
timestamp 1563080643
transform -1 0 124 0 1 105
box -2 -3 34 103
use INVX2  _975_
timestamp 1563080643
transform -1 0 140 0 1 105
box -2 -3 18 103
use NAND3X1  _1062_
timestamp 1563080643
transform 1 0 140 0 1 105
box -2 -3 34 103
use NAND3X1  _1033_
timestamp 1563080643
transform 1 0 172 0 1 105
box -2 -3 34 103
use NAND2X1  _1032_
timestamp 1563080643
transform 1 0 204 0 1 105
box -2 -3 26 103
use NAND3X1  _1101_
timestamp 1563080643
transform 1 0 228 0 1 105
box -2 -3 34 103
use NAND3X1  _1097_
timestamp 1563080643
transform 1 0 260 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert13
timestamp 1563080643
transform 1 0 292 0 1 105
box -2 -3 26 103
use NAND3X1  _1028_
timestamp 1563080643
transform 1 0 316 0 1 105
box -2 -3 34 103
use OR2X2  _1025_
timestamp 1563080643
transform -1 0 380 0 1 105
box -2 -3 34 103
use OR2X2  _1100_
timestamp 1563080643
transform -1 0 412 0 1 105
box -2 -3 34 103
use OR2X2  _1094_
timestamp 1563080643
transform -1 0 444 0 1 105
box -2 -3 34 103
use OAI21X1  _1031_
timestamp 1563080643
transform 1 0 444 0 1 105
box -2 -3 34 103
use INVX1  _1029_
timestamp 1563080643
transform -1 0 492 0 1 105
box -2 -3 18 103
use NAND3X1  _1390_
timestamp 1563080643
transform -1 0 524 0 1 105
box -2 -3 34 103
use OR2X2  _1387_
timestamp 1563080643
transform -1 0 556 0 1 105
box -2 -3 34 103
use OAI21X1  _1441_
timestamp 1563080643
transform -1 0 588 0 1 105
box -2 -3 34 103
use INVX1  _1439_
timestamp 1563080643
transform -1 0 604 0 1 105
box -2 -3 18 103
use FILL  FILL_1_0_0
timestamp 1563080643
transform 1 0 604 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1563080643
transform 1 0 612 0 1 105
box -2 -3 10 103
use INVX1  _1361_
timestamp 1563080643
transform 1 0 620 0 1 105
box -2 -3 18 103
use OAI21X1  _1363_
timestamp 1563080643
transform 1 0 636 0 1 105
box -2 -3 34 103
use NAND3X1  _1438_
timestamp 1563080643
transform -1 0 700 0 1 105
box -2 -3 34 103
use OR2X2  _1435_
timestamp 1563080643
transform 1 0 700 0 1 105
box -2 -3 34 103
use OAI21X1  _1324_
timestamp 1563080643
transform -1 0 764 0 1 105
box -2 -3 34 103
use INVX1  _1322_
timestamp 1563080643
transform -1 0 780 0 1 105
box -2 -3 18 103
use OR2X2  _1426_
timestamp 1563080643
transform 1 0 780 0 1 105
box -2 -3 34 103
use NAND3X1  _1429_
timestamp 1563080643
transform 1 0 812 0 1 105
box -2 -3 34 103
use NAND3X1  _1433_
timestamp 1563080643
transform 1 0 844 0 1 105
box -2 -3 34 103
use OR2X2  _1432_
timestamp 1563080643
transform -1 0 908 0 1 105
box -2 -3 34 103
use NAND3X1  _1321_
timestamp 1563080643
transform 1 0 908 0 1 105
box -2 -3 34 103
use OR2X2  _1318_
timestamp 1563080643
transform -1 0 972 0 1 105
box -2 -3 34 103
use NAND2X1  _1320_
timestamp 1563080643
transform 1 0 972 0 1 105
box -2 -3 26 103
use INVX1  _1319_
timestamp 1563080643
transform -1 0 1012 0 1 105
box -2 -3 18 103
use NAND3X1  _896_
timestamp 1563080643
transform -1 0 1044 0 1 105
box -2 -3 34 103
use OR2X2  _895_
timestamp 1563080643
transform 1 0 1044 0 1 105
box -2 -3 34 103
use NAND3X1  _892_
timestamp 1563080643
transform -1 0 1108 0 1 105
box -2 -3 34 103
use FILL  FILL_1_1_0
timestamp 1563080643
transform -1 0 1116 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1563080643
transform -1 0 1124 0 1 105
box -2 -3 10 103
use NAND3X1  _935_
timestamp 1563080643
transform -1 0 1156 0 1 105
box -2 -3 34 103
use OR2X2  _889_
timestamp 1563080643
transform -1 0 1188 0 1 105
box -2 -3 34 103
use OR2X2  _934_
timestamp 1563080643
transform -1 0 1220 0 1 105
box -2 -3 34 103
use NAND3X1  _931_
timestamp 1563080643
transform -1 0 1252 0 1 105
box -2 -3 34 103
use NAND3X1  _862_
timestamp 1563080643
transform -1 0 1284 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_insert22
timestamp 1563080643
transform 1 0 1284 0 1 105
box -2 -3 26 103
use OR2X2  _928_
timestamp 1563080643
transform -1 0 1340 0 1 105
box -2 -3 34 103
use OR2X2  _859_
timestamp 1563080643
transform -1 0 1372 0 1 105
box -2 -3 34 103
use INVX1  _1156_
timestamp 1563080643
transform 1 0 1372 0 1 105
box -2 -3 18 103
use OAI21X1  _1158_
timestamp 1563080643
transform -1 0 1420 0 1 105
box -2 -3 34 103
use OAI21X1  _865_
timestamp 1563080643
transform -1 0 1452 0 1 105
box -2 -3 34 103
use INVX1  _863_
timestamp 1563080643
transform -1 0 1468 0 1 105
box -2 -3 18 103
use NAND3X1  _1155_
timestamp 1563080643
transform -1 0 1500 0 1 105
box -2 -3 34 103
use OR2X2  _1152_
timestamp 1563080643
transform -1 0 1532 0 1 105
box -2 -3 34 103
use OAI21X1  _1275_
timestamp 1563080643
transform -1 0 1564 0 1 105
box -2 -3 34 103
use INVX1  _1273_
timestamp 1563080643
transform 1 0 1564 0 1 105
box -2 -3 18 103
use NAND3X1  _1267_
timestamp 1563080643
transform 1 0 1580 0 1 105
box -2 -3 34 103
use NAND3X1  _1263_
timestamp 1563080643
transform 1 0 1612 0 1 105
box -2 -3 34 103
use OAI21X1  _1197_
timestamp 1563080643
transform -1 0 1676 0 1 105
box -2 -3 34 103
use INVX1  _1195_
timestamp 1563080643
transform -1 0 1692 0 1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert7
timestamp 1563080643
transform -1 0 1716 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1563080643
transform 1 0 1716 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1563080643
transform 1 0 1724 0 1 105
box -2 -3 10 103
use NAND2X1  _1105_
timestamp 1563080643
transform 1 0 4 0 -1 105
box -2 -3 26 103
use NAND2X1  _991_
timestamp 1563080643
transform 1 0 28 0 -1 105
box -2 -3 26 103
use NAND2X1  _993_
timestamp 1563080643
transform 1 0 52 0 -1 105
box -2 -3 26 103
use OAI21X1  _992_
timestamp 1563080643
transform -1 0 108 0 -1 105
box -2 -3 34 103
use INVX1  _990_
timestamp 1563080643
transform -1 0 124 0 -1 105
box -2 -3 18 103
use OR2X2  _1061_
timestamp 1563080643
transform 1 0 124 0 -1 105
box -2 -3 34 103
use INVX1  _1104_
timestamp 1563080643
transform -1 0 172 0 -1 105
box -2 -3 18 103
use NAND2X1  _1110_
timestamp 1563080643
transform -1 0 196 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert12
timestamp 1563080643
transform 1 0 196 0 -1 105
box -2 -3 26 103
use NAND2X1  _1060_
timestamp 1563080643
transform 1 0 220 0 -1 105
box -2 -3 26 103
use INVX1  _1059_
timestamp 1563080643
transform -1 0 260 0 -1 105
box -2 -3 18 103
use NAND2X1  _1099_
timestamp 1563080643
transform 1 0 260 0 -1 105
box -2 -3 26 103
use NAND2X1  _1096_
timestamp 1563080643
transform 1 0 284 0 -1 105
box -2 -3 26 103
use INVX1  _1095_
timestamp 1563080643
transform -1 0 324 0 -1 105
box -2 -3 18 103
use NAND2X1  _1027_
timestamp 1563080643
transform 1 0 324 0 -1 105
box -2 -3 26 103
use NAND2X1  _1057_
timestamp 1563080643
transform 1 0 348 0 -1 105
box -2 -3 26 103
use NAND2X1  _1108_
timestamp 1563080643
transform 1 0 372 0 -1 105
box -2 -3 26 103
use OAI21X1  _1109_
timestamp 1563080643
transform -1 0 428 0 -1 105
box -2 -3 34 103
use INVX1  _1056_
timestamp 1563080643
transform -1 0 444 0 -1 105
box -2 -3 18 103
use INVX1  _1098_
timestamp 1563080643
transform -1 0 460 0 -1 105
box -2 -3 18 103
use NAND2X1  _1030_
timestamp 1563080643
transform 1 0 460 0 -1 105
box -2 -3 26 103
use INVX1  _1107_
timestamp 1563080643
transform -1 0 500 0 -1 105
box -2 -3 18 103
use INVX1  _1388_
timestamp 1563080643
transform -1 0 516 0 -1 105
box -2 -3 18 103
use NAND2X1  _1389_
timestamp 1563080643
transform -1 0 540 0 -1 105
box -2 -3 26 103
use NAND2X1  _1440_
timestamp 1563080643
transform 1 0 540 0 -1 105
box -2 -3 26 103
use NAND2X1  _1362_
timestamp 1563080643
transform -1 0 588 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_insert2
timestamp 1563080643
transform 1 0 588 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_0
timestamp 1563080643
transform 1 0 612 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1563080643
transform 1 0 620 0 -1 105
box -2 -3 10 103
use NAND2X1  _1437_
timestamp 1563080643
transform 1 0 628 0 -1 105
box -2 -3 26 103
use INVX1  _1436_
timestamp 1563080643
transform 1 0 652 0 -1 105
box -2 -3 18 103
use INVX1  _1026_
timestamp 1563080643
transform -1 0 684 0 -1 105
box -2 -3 18 103
use NAND2X1  _1323_
timestamp 1563080643
transform -1 0 708 0 -1 105
box -2 -3 26 103
use NAND2X1  _1428_
timestamp 1563080643
transform 1 0 708 0 -1 105
box -2 -3 26 103
use INVX1  _1427_
timestamp 1563080643
transform -1 0 748 0 -1 105
box -2 -3 18 103
use NAND2X1  _1359_
timestamp 1563080643
transform 1 0 748 0 -1 105
box -2 -3 26 103
use INVX1  _1358_
timestamp 1563080643
transform -1 0 788 0 -1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert1
timestamp 1563080643
transform 1 0 788 0 -1 105
box -2 -3 26 103
use INVX1  _1430_
timestamp 1563080643
transform 1 0 812 0 -1 105
box -2 -3 18 103
use NAND2X1  _1431_
timestamp 1563080643
transform -1 0 852 0 -1 105
box -2 -3 26 103
use INVX1  _893_
timestamp 1563080643
transform 1 0 852 0 -1 105
box -2 -3 18 103
use NAND2X1  _894_
timestamp 1563080643
transform -1 0 892 0 -1 105
box -2 -3 26 103
use NAND2X1  _891_
timestamp 1563080643
transform 1 0 892 0 -1 105
box -2 -3 26 103
use INVX1  _890_
timestamp 1563080643
transform -1 0 932 0 -1 105
box -2 -3 18 103
use NAND2X1  _825_
timestamp 1563080643
transform 1 0 932 0 -1 105
box -2 -3 26 103
use INVX1  _824_
timestamp 1563080643
transform 1 0 956 0 -1 105
box -2 -3 18 103
use OAI21X1  _826_
timestamp 1563080643
transform -1 0 1004 0 -1 105
box -2 -3 34 103
use NAND2X1  _827_
timestamp 1563080643
transform -1 0 1028 0 -1 105
box -2 -3 26 103
use NAND2X1  _933_
timestamp 1563080643
transform 1 0 1028 0 -1 105
box -2 -3 26 103
use INVX1  _932_
timestamp 1563080643
transform -1 0 1068 0 -1 105
box -2 -3 18 103
use INVX1  _929_
timestamp 1563080643
transform 1 0 1068 0 -1 105
box -2 -3 18 103
use NAND2X1  _930_
timestamp 1563080643
transform -1 0 1108 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_1_0
timestamp 1563080643
transform 1 0 1108 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1563080643
transform 1 0 1116 0 -1 105
box -2 -3 10 103
use NAND2X1  _942_
timestamp 1563080643
transform 1 0 1124 0 -1 105
box -2 -3 26 103
use OAI21X1  _943_
timestamp 1563080643
transform -1 0 1180 0 -1 105
box -2 -3 34 103
use INVX1  _941_
timestamp 1563080643
transform -1 0 1196 0 -1 105
box -2 -3 18 103
use BUFX2  BUFX2_insert24
timestamp 1563080643
transform -1 0 1220 0 -1 105
box -2 -3 26 103
use NAND2X1  _864_
timestamp 1563080643
transform 1 0 1220 0 -1 105
box -2 -3 26 103
use NAND2X1  _861_
timestamp 1563080643
transform 1 0 1244 0 -1 105
box -2 -3 26 103
use INVX1  _860_
timestamp 1563080643
transform -1 0 1284 0 -1 105
box -2 -3 18 103
use INVX1  _1261_
timestamp 1563080643
transform 1 0 1284 0 -1 105
box -2 -3 18 103
use INVX1  _1222_
timestamp 1563080643
transform 1 0 1300 0 -1 105
box -2 -3 18 103
use NAND2X1  _1223_
timestamp 1563080643
transform -1 0 1340 0 -1 105
box -2 -3 26 103
use INVX1  _1264_
timestamp 1563080643
transform 1 0 1340 0 -1 105
box -2 -3 18 103
use NAND2X1  _1262_
timestamp 1563080643
transform -1 0 1380 0 -1 105
box -2 -3 26 103
use NAND2X1  _1157_
timestamp 1563080643
transform -1 0 1404 0 -1 105
box -2 -3 26 103
use NAND2X1  _1274_
timestamp 1563080643
transform -1 0 1428 0 -1 105
box -2 -3 26 103
use INVX1  _1192_
timestamp 1563080643
transform 1 0 1428 0 -1 105
box -2 -3 18 103
use NAND2X1  _1193_
timestamp 1563080643
transform -1 0 1468 0 -1 105
box -2 -3 26 103
use NAND2X1  _1196_
timestamp 1563080643
transform -1 0 1492 0 -1 105
box -2 -3 26 103
use NAND2X1  _1265_
timestamp 1563080643
transform -1 0 1516 0 -1 105
box -2 -3 26 103
use OR2X2  _1260_
timestamp 1563080643
transform 1 0 1516 0 -1 105
box -2 -3 34 103
use OR2X2  _1266_
timestamp 1563080643
transform 1 0 1548 0 -1 105
box -2 -3 34 103
use INVX2  _1477_
timestamp 1563080643
transform -1 0 1596 0 -1 105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_insert48
timestamp 1563080643
transform -1 0 1668 0 -1 105
box -2 -3 74 103
use BUFX2  BUFX2_insert5
timestamp 1563080643
transform -1 0 1692 0 -1 105
box -2 -3 26 103
use AND2X2  _775_
timestamp 1563080643
transform 1 0 1692 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1563080643
transform -1 0 1732 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 600 -30 616 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 1112 -30 1128 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s 1758 658 1762 662 3 FreeSans 24 0 0 0 CLK
port 2 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 DATA_A[31]
port 3 nsew
flabel metal2 s 62 1638 66 1642 7 FreeSans 24 90 0 0 DATA_A[30]
port 4 nsew
flabel metal2 s 446 1638 450 1642 3 FreeSans 24 90 0 0 DATA_A[29]
port 5 nsew
flabel metal2 s 646 1638 650 1642 3 FreeSans 24 90 0 0 DATA_A[28]
port 6 nsew
flabel metal3 s -26 778 -22 782 7 FreeSans 24 0 0 0 DATA_A[27]
port 7 nsew
flabel metal3 s -26 578 -22 582 7 FreeSans 24 0 0 0 DATA_A[26]
port 8 nsew
flabel metal3 s -26 558 -22 562 7 FreeSans 24 0 0 0 DATA_A[25]
port 9 nsew
flabel metal3 s -26 1098 -22 1102 7 FreeSans 24 0 0 0 DATA_A[24]
port 10 nsew
flabel metal3 s -26 818 -22 822 7 FreeSans 24 0 0 0 DATA_A[23]
port 11 nsew
flabel metal3 s -26 1458 -22 1462 7 FreeSans 24 0 0 0 DATA_A[22]
port 12 nsew
flabel metal2 s 766 1638 770 1642 3 FreeSans 24 90 0 0 DATA_A[21]
port 13 nsew
flabel metal2 s 726 1638 730 1642 3 FreeSans 24 90 0 0 DATA_A[20]
port 14 nsew
flabel metal3 s -26 968 -22 972 7 FreeSans 24 0 0 0 DATA_A[19]
port 15 nsew
flabel metal3 s -26 898 -22 902 7 FreeSans 24 0 0 0 DATA_A[18]
port 16 nsew
flabel metal3 s -26 1058 -22 1062 7 FreeSans 24 0 0 0 DATA_A[17]
port 17 nsew
flabel metal3 s -26 1128 -22 1132 7 FreeSans 24 0 0 0 DATA_A[16]
port 18 nsew
flabel metal3 s -26 538 -22 542 7 FreeSans 24 0 0 0 DATA_A[15]
port 19 nsew
flabel metal3 s -26 1528 -22 1532 7 FreeSans 24 0 0 0 DATA_A[14]
port 20 nsew
flabel metal2 s 294 1638 298 1642 3 FreeSans 24 90 0 0 DATA_A[13]
port 21 nsew
flabel metal2 s 566 1638 570 1642 3 FreeSans 24 90 0 0 DATA_A[12]
port 22 nsew
flabel metal3 s -26 738 -22 742 7 FreeSans 24 0 0 0 DATA_A[11]
port 23 nsew
flabel metal3 s -26 508 -22 512 7 FreeSans 24 0 0 0 DATA_A[10]
port 24 nsew
flabel metal3 s -26 598 -22 602 7 FreeSans 24 0 0 0 DATA_A[9]
port 25 nsew
flabel metal3 s -26 878 -22 882 7 FreeSans 24 0 0 0 DATA_A[8]
port 26 nsew
flabel metal3 s -26 698 -22 702 7 FreeSans 24 0 0 0 DATA_A[7]
port 27 nsew
flabel metal3 s -26 1478 -22 1482 7 FreeSans 24 0 0 0 DATA_A[6]
port 28 nsew
flabel metal3 s -26 1348 -22 1352 7 FreeSans 24 0 0 0 DATA_A[5]
port 29 nsew
flabel metal2 s 630 1638 634 1642 3 FreeSans 24 90 0 0 DATA_A[4]
port 30 nsew
flabel metal3 s -26 858 -22 862 7 FreeSans 24 0 0 0 DATA_A[3]
port 31 nsew
flabel metal3 s -26 758 -22 762 7 FreeSans 24 0 0 0 DATA_A[2]
port 32 nsew
flabel metal3 s -26 1078 -22 1082 7 FreeSans 24 0 0 0 DATA_A[1]
port 33 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 DATA_A[0]
port 34 nsew
flabel metal3 s 1758 608 1762 612 3 FreeSans 24 0 0 0 DATA_B[31]
port 35 nsew
flabel metal2 s 46 -22 50 -18 7 FreeSans 24 270 0 0 DATA_B[30]
port 36 nsew
flabel metal2 s 1078 -22 1082 -18 7 FreeSans 24 270 0 0 DATA_B[29]
port 37 nsew
flabel metal2 s 862 -22 866 -18 7 FreeSans 24 270 0 0 DATA_B[28]
port 38 nsew
flabel metal2 s 1262 -22 1266 -18 7 FreeSans 24 270 0 0 DATA_B[27]
port 39 nsew
flabel metal3 s 1758 548 1762 552 3 FreeSans 24 0 0 0 DATA_B[26]
port 40 nsew
flabel metal2 s 1150 -22 1154 -18 7 FreeSans 24 270 0 0 DATA_B[25]
port 41 nsew
flabel metal3 s 1758 488 1762 492 3 FreeSans 24 0 0 0 DATA_B[24]
port 42 nsew
flabel metal3 s 1758 588 1762 592 3 FreeSans 24 0 0 0 DATA_B[23]
port 43 nsew
flabel metal2 s 1022 -22 1026 -18 7 FreeSans 24 270 0 0 DATA_B[22]
port 44 nsew
flabel metal2 s 1134 -22 1138 -18 7 FreeSans 24 270 0 0 DATA_B[21]
port 45 nsew
flabel metal2 s 918 -22 922 -18 7 FreeSans 24 270 0 0 DATA_B[20]
port 46 nsew
flabel metal2 s 1278 -22 1282 -18 7 FreeSans 24 270 0 0 DATA_B[19]
port 47 nsew
flabel metal3 s -26 298 -22 302 7 FreeSans 24 0 0 0 DATA_B[18]
port 48 nsew
flabel metal2 s 1062 -22 1066 -18 7 FreeSans 24 270 0 0 DATA_B[17]
port 49 nsew
flabel metal3 s 1758 328 1762 332 3 FreeSans 24 0 0 0 DATA_B[16]
port 50 nsew
flabel metal3 s 1758 528 1762 532 3 FreeSans 24 0 0 0 DATA_B[15]
port 51 nsew
flabel metal2 s 134 -22 138 -18 7 FreeSans 24 270 0 0 DATA_B[14]
port 52 nsew
flabel metal2 s 1558 -22 1562 -18 7 FreeSans 24 270 0 0 DATA_B[13]
port 53 nsew
flabel metal2 s 158 -22 162 -18 7 FreeSans 24 270 0 0 DATA_B[12]
port 54 nsew
flabel metal3 s 1758 148 1762 152 3 FreeSans 24 0 0 0 DATA_B[11]
port 55 nsew
flabel metal3 s -26 488 -22 492 7 FreeSans 24 0 0 0 DATA_B[10]
port 56 nsew
flabel metal2 s 1198 -22 1202 -18 7 FreeSans 24 270 0 0 DATA_B[9]
port 57 nsew
flabel metal3 s 1758 568 1762 572 3 FreeSans 24 0 0 0 DATA_B[8]
port 58 nsew
flabel metal3 s 1758 508 1762 512 3 FreeSans 24 0 0 0 DATA_B[7]
port 59 nsew
flabel metal2 s 982 -22 986 -18 7 FreeSans 24 270 0 0 DATA_B[6]
port 60 nsew
flabel metal2 s 1526 -22 1530 -18 7 FreeSans 24 270 0 0 DATA_B[5]
port 61 nsew
flabel metal2 s 1222 -22 1226 -18 7 FreeSans 24 270 0 0 DATA_B[4]
port 62 nsew
flabel metal2 s 1326 -22 1330 -18 7 FreeSans 24 270 0 0 DATA_B[3]
port 63 nsew
flabel metal3 s -26 278 -22 282 7 FreeSans 24 0 0 0 DATA_B[2]
port 64 nsew
flabel metal3 s -26 178 -22 182 7 FreeSans 24 0 0 0 DATA_B[1]
port 65 nsew
flabel metal3 s 1758 268 1762 272 3 FreeSans 24 0 0 0 DATA_B[0]
port 66 nsew
flabel metal3 s 1758 698 1762 702 3 FreeSans 24 0 0 0 DATA_OUT[3]
port 67 nsew
flabel metal3 s 1758 848 1762 852 3 FreeSans 24 0 0 0 DATA_OUT[2]
port 68 nsew
flabel metal3 s 1758 628 1762 632 3 FreeSans 24 0 0 0 DATA_OUT[1]
port 69 nsew
flabel metal3 s 1758 678 1762 682 3 FreeSans 24 0 0 0 DATA_OUT[0]
port 70 nsew
flabel metal2 s 1230 1638 1234 1642 3 FreeSans 24 90 0 0 RESET_L
port 71 nsew
flabel metal2 s 198 1638 202 1642 3 FreeSans 24 90 0 0 SEL_A[11]
port 72 nsew
flabel metal3 s -26 1278 -22 1282 7 FreeSans 24 0 0 0 SEL_A[10]
port 73 nsew
flabel metal3 s -26 1248 -22 1252 7 FreeSans 24 0 0 0 SEL_A[9]
port 74 nsew
flabel metal2 s 414 1638 418 1642 3 FreeSans 24 90 0 0 SEL_A[8]
port 75 nsew
flabel metal2 s 694 1638 698 1642 3 FreeSans 24 90 0 0 SEL_A[7]
port 76 nsew
flabel metal2 s 670 1638 674 1642 3 FreeSans 24 90 0 0 SEL_A[6]
port 77 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 SEL_A[5]
port 78 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 SEL_A[4]
port 79 nsew
flabel metal3 s -26 798 -22 802 7 FreeSans 24 0 0 0 SEL_A[3]
port 80 nsew
flabel metal2 s 550 1638 554 1642 3 FreeSans 24 90 0 0 SEL_A[2]
port 81 nsew
flabel metal2 s 750 1638 754 1642 3 FreeSans 24 90 0 0 SEL_A[1]
port 82 nsew
flabel metal2 s 710 1638 714 1642 3 FreeSans 24 90 0 0 SEL_A[0]
port 83 nsew
flabel metal3 s -26 678 -22 682 7 FreeSans 24 0 0 0 SEL_AB[3]
port 84 nsew
flabel metal3 s 1758 358 1762 362 3 FreeSans 24 0 0 0 SEL_AB[2]
port 85 nsew
flabel metal3 s -26 468 -22 472 7 FreeSans 24 0 0 0 SEL_AB[1]
port 86 nsew
flabel metal2 s 1166 -22 1170 -18 7 FreeSans 24 270 0 0 SEL_AB[0]
port 87 nsew
flabel metal2 s 814 -22 818 -18 7 FreeSans 24 270 0 0 SEL_B[11]
port 88 nsew
flabel metal2 s 838 -22 842 -18 7 FreeSans 24 270 0 0 SEL_B[10]
port 89 nsew
flabel metal2 s 798 -22 802 -18 7 FreeSans 24 270 0 0 SEL_B[9]
port 90 nsew
flabel metal3 s 1758 58 1762 62 3 FreeSans 24 270 0 0 SEL_B[8]
port 91 nsew
flabel metal3 s 1758 468 1762 472 3 FreeSans 24 0 0 0 SEL_B[7]
port 92 nsew
flabel metal3 s 1758 448 1762 452 3 FreeSans 24 0 0 0 SEL_B[6]
port 93 nsew
flabel metal2 s 294 -22 298 -18 7 FreeSans 24 270 0 0 SEL_B[5]
port 94 nsew
flabel metal3 s -26 158 -22 162 7 FreeSans 24 0 0 0 SEL_B[4]
port 95 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 0 0 0 SEL_B[3]
port 96 nsew
flabel metal2 s 1238 -22 1242 -18 7 FreeSans 24 270 0 0 SEL_B[2]
port 97 nsew
flabel metal2 s 1038 -22 1042 -18 7 FreeSans 24 270 0 0 SEL_B[1]
port 98 nsew
flabel metal2 s 1102 -22 1106 -18 7 FreeSans 24 270 0 0 SEL_B[0]
port 99 nsew
<< end >>
