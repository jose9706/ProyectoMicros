/*
 *Universidad de Costa Rica - Escuela de Ingenieria Electrica
 *Proyecto #1 - IE-0411 - Arvhivo de includes 
 *@author Giancarlo Marin H.
 *@date   08/06/2019
 *@brief  Contiene la lsiatd e archivos necesarios para crear el selector de nibble mayor
*/

// Si no se ha creado 
`ifndef _my_incl_vh_
`define _my_incl_vh_

// includes
`include "../Selector/selector4.v"
`include "../nm2/nm2.v"

`endif

